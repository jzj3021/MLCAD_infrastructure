module fpu (clk,
    div_by_zero,
    ine,
    inf,
    overflow,
    qnan,
    snan,
    underflow,
    zero,
    fpu_op,
    opa,
    opb,
    out,
    rmode);
 input clk;
 output div_by_zero;
 output ine;
 output inf;
 output overflow;
 output qnan;
 output snan;
 output underflow;
 output zero;
 input [2:0] fpu_op;
 input [31:0] opa;
 input [31:0] opb;
 output [31:0] out;
 input [1:0] rmode;

 wire UNCONNECTED;
 wire UNCONNECTED0;
 wire UNCONNECTED1;
 wire UNCONNECTED10;
 wire UNCONNECTED100;
 wire UNCONNECTED101;
 wire UNCONNECTED102;
 wire UNCONNECTED103;
 wire UNCONNECTED104;
 wire UNCONNECTED105;
 wire UNCONNECTED106;
 wire UNCONNECTED107;
 wire UNCONNECTED108;
 wire UNCONNECTED109;
 wire UNCONNECTED11;
 wire UNCONNECTED110;
 wire UNCONNECTED111;
 wire UNCONNECTED112;
 wire UNCONNECTED113;
 wire UNCONNECTED114;
 wire UNCONNECTED115;
 wire UNCONNECTED116;
 wire UNCONNECTED117;
 wire UNCONNECTED118;
 wire UNCONNECTED119;
 wire UNCONNECTED12;
 wire UNCONNECTED120;
 wire UNCONNECTED121;
 wire UNCONNECTED122;
 wire UNCONNECTED123;
 wire UNCONNECTED124;
 wire UNCONNECTED125;
 wire UNCONNECTED126;
 wire UNCONNECTED127;
 wire UNCONNECTED128;
 wire UNCONNECTED129;
 wire UNCONNECTED13;
 wire UNCONNECTED130;
 wire UNCONNECTED131;
 wire UNCONNECTED132;
 wire UNCONNECTED133;
 wire UNCONNECTED134;
 wire UNCONNECTED135;
 wire UNCONNECTED136;
 wire UNCONNECTED137;
 wire UNCONNECTED138;
 wire UNCONNECTED139;
 wire UNCONNECTED14;
 wire UNCONNECTED140;
 wire UNCONNECTED141;
 wire UNCONNECTED142;
 wire UNCONNECTED143;
 wire UNCONNECTED144;
 wire UNCONNECTED145;
 wire UNCONNECTED146;
 wire UNCONNECTED147;
 wire UNCONNECTED148;
 wire UNCONNECTED149;
 wire UNCONNECTED15;
 wire UNCONNECTED150;
 wire UNCONNECTED151;
 wire UNCONNECTED152;
 wire UNCONNECTED153;
 wire UNCONNECTED154;
 wire UNCONNECTED155;
 wire UNCONNECTED156;
 wire UNCONNECTED157;
 wire UNCONNECTED158;
 wire UNCONNECTED159;
 wire UNCONNECTED16;
 wire UNCONNECTED160;
 wire UNCONNECTED161;
 wire UNCONNECTED162;
 wire UNCONNECTED163;
 wire UNCONNECTED164;
 wire UNCONNECTED165;
 wire UNCONNECTED166;
 wire UNCONNECTED167;
 wire UNCONNECTED168;
 wire UNCONNECTED169;
 wire UNCONNECTED17;
 wire UNCONNECTED170;
 wire UNCONNECTED171;
 wire UNCONNECTED172;
 wire UNCONNECTED173;
 wire UNCONNECTED174;
 wire UNCONNECTED175;
 wire UNCONNECTED176;
 wire UNCONNECTED177;
 wire UNCONNECTED178;
 wire UNCONNECTED179;
 wire UNCONNECTED18;
 wire UNCONNECTED180;
 wire UNCONNECTED181;
 wire UNCONNECTED182;
 wire UNCONNECTED183;
 wire UNCONNECTED184;
 wire UNCONNECTED185;
 wire UNCONNECTED186;
 wire UNCONNECTED187;
 wire UNCONNECTED188;
 wire UNCONNECTED189;
 wire UNCONNECTED19;
 wire UNCONNECTED190;
 wire UNCONNECTED191;
 wire UNCONNECTED2;
 wire UNCONNECTED20;
 wire UNCONNECTED21;
 wire UNCONNECTED22;
 wire UNCONNECTED23;
 wire UNCONNECTED24;
 wire UNCONNECTED25;
 wire UNCONNECTED26;
 wire UNCONNECTED27;
 wire UNCONNECTED28;
 wire UNCONNECTED29;
 wire UNCONNECTED3;
 wire UNCONNECTED30;
 wire UNCONNECTED31;
 wire UNCONNECTED32;
 wire UNCONNECTED33;
 wire UNCONNECTED34;
 wire UNCONNECTED35;
 wire UNCONNECTED36;
 wire UNCONNECTED37;
 wire UNCONNECTED38;
 wire UNCONNECTED39;
 wire UNCONNECTED4;
 wire UNCONNECTED40;
 wire UNCONNECTED41;
 wire UNCONNECTED42;
 wire UNCONNECTED43;
 wire UNCONNECTED44;
 wire UNCONNECTED45;
 wire UNCONNECTED46;
 wire UNCONNECTED47;
 wire UNCONNECTED48;
 wire UNCONNECTED49;
 wire UNCONNECTED5;
 wire UNCONNECTED50;
 wire UNCONNECTED51;
 wire UNCONNECTED52;
 wire UNCONNECTED53;
 wire UNCONNECTED54;
 wire UNCONNECTED55;
 wire UNCONNECTED56;
 wire UNCONNECTED57;
 wire UNCONNECTED58;
 wire UNCONNECTED59;
 wire UNCONNECTED6;
 wire UNCONNECTED60;
 wire UNCONNECTED61;
 wire UNCONNECTED62;
 wire UNCONNECTED63;
 wire UNCONNECTED64;
 wire UNCONNECTED65;
 wire UNCONNECTED66;
 wire UNCONNECTED67;
 wire UNCONNECTED68;
 wire UNCONNECTED69;
 wire UNCONNECTED7;
 wire UNCONNECTED70;
 wire UNCONNECTED71;
 wire UNCONNECTED72;
 wire UNCONNECTED73;
 wire UNCONNECTED74;
 wire UNCONNECTED75;
 wire UNCONNECTED76;
 wire UNCONNECTED77;
 wire UNCONNECTED78;
 wire UNCONNECTED79;
 wire UNCONNECTED8;
 wire UNCONNECTED80;
 wire UNCONNECTED81;
 wire UNCONNECTED82;
 wire UNCONNECTED83;
 wire UNCONNECTED84;
 wire UNCONNECTED85;
 wire UNCONNECTED86;
 wire UNCONNECTED87;
 wire UNCONNECTED88;
 wire UNCONNECTED89;
 wire UNCONNECTED9;
 wire UNCONNECTED90;
 wire UNCONNECTED91;
 wire UNCONNECTED92;
 wire UNCONNECTED93;
 wire UNCONNECTED94;
 wire UNCONNECTED95;
 wire UNCONNECTED96;
 wire UNCONNECTED97;
 wire UNCONNECTED98;
 wire UNCONNECTED99;
 wire fasu_op;
 wire fasu_op_r1;
 wire fasu_op_r2;
 wire inc_u4_add_230_34_n_185;
 wire inc_u4_add_230_34_n_189;
 wire inc_u4_add_230_34_n_192;
 wire inc_u4_add_230_34_n_196;
 wire inc_u4_add_230_34_n_200;
 wire inc_u4_add_230_34_n_203;
 wire inc_u4_add_230_34_n_204;
 wire inc_u4_add_230_34_n_208;
 wire inc_u4_add_230_34_n_209;
 wire inc_u4_add_230_34_n_213;
 wire inc_u4_add_230_34_n_217;
 wire inc_u4_add_230_34_n_221;
 wire inc_u4_add_230_34_n_226;
 wire inc_u4_add_230_34_n_230;
 wire inc_u4_add_230_34_n_235;
 wire inc_u4_add_230_34_n_239;
 wire inc_u4_add_230_34_n_242;
 wire inc_u4_add_230_34_n_246;
 wire inc_u4_add_230_34_n_250;
 wire inc_u4_add_230_34_n_254;
 wire inc_u4_add_230_34_n_259;
 wire inc_u4_add_230_34_n_263;
 wire inc_u4_add_230_34_n_267;
 wire inc_u4_add_230_34_n_270;
 wire inc_u4_add_230_34_n_272;
 wire inc_u4_add_230_34_n_274;
 wire inc_u4_add_230_34_n_277;
 wire inc_u4_add_230_34_n_278;
 wire inc_u4_add_230_34_n_280;
 wire inc_u4_add_230_34_n_284;
 wire inc_u4_add_230_34_n_286;
 wire inc_u4_add_230_34_n_289;
 wire inc_u4_add_230_34_n_290;
 wire ind_d;
 wire inf_d;
 wire inf_mul;
 wire inf_mul2;
 wire inf_mul_r;
 wire n_1;
 wire n_10;
 wire n_100;
 wire n_1000;
 wire n_1001;
 wire n_1002;
 wire n_1003;
 wire n_1004;
 wire n_1005;
 wire n_1006;
 wire n_1007;
 wire n_1008;
 wire n_1009;
 wire n_101;
 wire n_1010;
 wire n_1011;
 wire n_1014;
 wire n_1015;
 wire n_1016;
 wire n_1017;
 wire n_1018;
 wire n_1019;
 wire n_102;
 wire n_1020;
 wire n_1021;
 wire n_1022;
 wire n_1023;
 wire n_1024;
 wire n_1025;
 wire n_1026;
 wire n_1027;
 wire n_1028;
 wire n_1029;
 wire n_103;
 wire n_1032;
 wire n_1033;
 wire n_1034;
 wire n_1035;
 wire n_1036;
 wire n_1037;
 wire n_1038;
 wire n_1039;
 wire n_104;
 wire n_1040;
 wire n_1042;
 wire n_1044;
 wire n_1045;
 wire n_1046;
 wire n_1047;
 wire n_1048;
 wire n_1049;
 wire n_105;
 wire n_1050;
 wire n_1051;
 wire n_1052;
 wire n_1053;
 wire n_1054;
 wire n_1055;
 wire n_1056;
 wire n_1057;
 wire n_1058;
 wire n_1059;
 wire n_106;
 wire n_1060;
 wire n_1061;
 wire n_1063;
 wire n_1064;
 wire n_1065;
 wire n_1066;
 wire n_1067;
 wire n_1068;
 wire n_1069;
 wire n_107;
 wire n_1070;
 wire n_1071;
 wire n_1072;
 wire n_1073;
 wire n_1074;
 wire n_1075;
 wire n_1076;
 wire n_1077;
 wire n_1078;
 wire n_1079;
 wire n_108;
 wire n_1080;
 wire n_1081;
 wire n_1082;
 wire n_1083;
 wire n_1084;
 wire n_1085;
 wire n_1086;
 wire n_1087;
 wire n_1088;
 wire n_1089;
 wire n_109;
 wire n_1090;
 wire n_1091;
 wire n_1092;
 wire n_1093;
 wire n_1094;
 wire n_1095;
 wire n_1096;
 wire n_1097;
 wire n_1098;
 wire n_1099;
 wire n_11;
 wire n_110;
 wire n_1100;
 wire n_1101;
 wire n_1102;
 wire n_1103;
 wire n_1104;
 wire n_1105;
 wire n_1106;
 wire n_1107;
 wire n_1108;
 wire n_1109;
 wire n_1110;
 wire n_1111;
 wire n_1112;
 wire n_1113;
 wire n_1114;
 wire n_1115;
 wire n_1116;
 wire n_1117;
 wire n_1118;
 wire n_1119;
 wire n_112;
 wire n_1120;
 wire n_1121;
 wire n_1122;
 wire n_1123;
 wire n_1124;
 wire n_1125;
 wire n_1126;
 wire n_1127;
 wire n_1128;
 wire n_1129;
 wire n_113;
 wire n_1130;
 wire n_1131;
 wire n_1132;
 wire n_1133;
 wire n_1134;
 wire n_1135;
 wire n_1136;
 wire n_1137;
 wire n_1138;
 wire n_1139;
 wire n_114;
 wire n_1140;
 wire n_1141;
 wire n_1142;
 wire n_1143;
 wire n_1144;
 wire n_1145;
 wire n_1146;
 wire n_1147;
 wire n_1148;
 wire n_1149;
 wire n_115;
 wire n_1150;
 wire n_1151;
 wire n_1152;
 wire n_1153;
 wire n_1154;
 wire n_1155;
 wire n_1156;
 wire n_1157;
 wire n_1158;
 wire n_1159;
 wire n_116;
 wire n_1160;
 wire n_1161;
 wire n_1162;
 wire n_1163;
 wire n_1164;
 wire n_1165;
 wire n_1166;
 wire n_1167;
 wire n_1168;
 wire n_1169;
 wire n_117;
 wire n_1170;
 wire n_1171;
 wire n_1172;
 wire n_1173;
 wire n_1174;
 wire n_1175;
 wire n_1176;
 wire n_1177;
 wire n_1178;
 wire n_1179;
 wire n_118;
 wire n_1180;
 wire n_1181;
 wire n_1182;
 wire n_1183;
 wire n_1184;
 wire n_1185;
 wire n_1186;
 wire n_1187;
 wire n_1188;
 wire n_1189;
 wire n_119;
 wire n_1190;
 wire n_1191;
 wire n_1192;
 wire n_1193;
 wire n_1194;
 wire n_1195;
 wire n_1196;
 wire n_1197;
 wire n_1198;
 wire n_1199;
 wire n_12;
 wire n_120;
 wire n_1200;
 wire n_1201;
 wire n_1202;
 wire n_1203;
 wire n_1204;
 wire n_1205;
 wire n_1206;
 wire n_1207;
 wire n_1208;
 wire n_1209;
 wire n_121;
 wire n_1210;
 wire n_1211;
 wire n_1212;
 wire n_1213;
 wire n_1214;
 wire n_1215;
 wire n_1216;
 wire n_1217;
 wire n_1218;
 wire n_1219;
 wire n_122;
 wire n_1220;
 wire n_1221;
 wire n_1222;
 wire n_1223;
 wire n_1224;
 wire n_1225;
 wire n_1226;
 wire n_1227;
 wire n_1228;
 wire n_1229;
 wire n_123;
 wire n_1230;
 wire n_1231;
 wire n_1232;
 wire n_1233;
 wire n_1234;
 wire n_1235;
 wire n_1236;
 wire n_1237;
 wire n_1238;
 wire n_1239;
 wire n_124;
 wire n_1240;
 wire n_1241;
 wire n_1242;
 wire n_1243;
 wire n_1244;
 wire n_1245;
 wire n_1246;
 wire n_1247;
 wire n_1248;
 wire n_1249;
 wire n_125;
 wire n_1250;
 wire n_1251;
 wire n_1252;
 wire n_1253;
 wire n_1254;
 wire n_1255;
 wire n_1256;
 wire n_1257;
 wire n_1258;
 wire n_1259;
 wire n_126;
 wire n_1260;
 wire n_1261;
 wire n_1262;
 wire n_1263;
 wire n_1264;
 wire n_1265;
 wire n_1266;
 wire n_1267;
 wire n_1268;
 wire n_1269;
 wire n_127;
 wire n_1270;
 wire n_1271;
 wire n_1272;
 wire n_1273;
 wire n_1274;
 wire n_1275;
 wire n_1276;
 wire n_1279;
 wire n_128;
 wire n_1281;
 wire n_1282;
 wire n_1283;
 wire n_1284;
 wire n_1285;
 wire n_1286;
 wire n_1287;
 wire n_1289;
 wire n_129;
 wire n_1290;
 wire n_1291;
 wire n_1292;
 wire n_1293;
 wire n_1294;
 wire n_1295;
 wire n_1296;
 wire n_1297;
 wire n_1298;
 wire n_1299;
 wire n_13;
 wire n_130;
 wire n_1300;
 wire n_1302;
 wire n_1303;
 wire n_1304;
 wire n_1305;
 wire n_1306;
 wire n_1307;
 wire n_1308;
 wire n_1309;
 wire n_131;
 wire n_1310;
 wire n_1311;
 wire n_1312;
 wire n_1313;
 wire n_1314;
 wire n_1315;
 wire n_1316;
 wire n_1317;
 wire n_1318;
 wire n_1319;
 wire n_132;
 wire n_1320;
 wire n_1321;
 wire n_1322;
 wire n_1323;
 wire n_1324;
 wire n_1325;
 wire n_1326;
 wire n_1327;
 wire n_1328;
 wire n_1329;
 wire n_133;
 wire n_1330;
 wire n_1331;
 wire n_1332;
 wire n_1333;
 wire n_1334;
 wire n_1335;
 wire n_1336;
 wire n_1337;
 wire n_1338;
 wire n_1339;
 wire n_134;
 wire n_1340;
 wire n_1341;
 wire n_1342;
 wire n_1343;
 wire n_1344;
 wire n_1345;
 wire n_1346;
 wire n_1347;
 wire n_1348;
 wire n_1349;
 wire n_135;
 wire n_1350;
 wire n_1351;
 wire n_1352;
 wire n_1353;
 wire n_1354;
 wire n_1355;
 wire n_1356;
 wire n_1357;
 wire n_1358;
 wire n_1359;
 wire n_136;
 wire n_1360;
 wire n_1361;
 wire n_1362;
 wire n_1363;
 wire n_1364;
 wire n_1365;
 wire n_1366;
 wire n_1367;
 wire n_1368;
 wire n_1369;
 wire n_137;
 wire n_1370;
 wire n_1371;
 wire n_1372;
 wire n_1373;
 wire n_1374;
 wire n_1375;
 wire n_1376;
 wire n_1377;
 wire n_1378;
 wire n_1379;
 wire n_138;
 wire n_1380;
 wire n_1381;
 wire n_1382;
 wire n_1383;
 wire n_13834;
 wire n_13835;
 wire n_13836;
 wire n_13837;
 wire n_13838;
 wire n_13839;
 wire n_1384;
 wire n_13840;
 wire n_13841;
 wire n_13842;
 wire n_13843;
 wire n_13844;
 wire n_13845;
 wire n_13846;
 wire n_13847;
 wire n_13848;
 wire n_13849;
 wire n_1385;
 wire n_13850;
 wire n_13851;
 wire n_13852;
 wire n_13856;
 wire n_13857;
 wire n_13858;
 wire n_13859;
 wire n_1386;
 wire n_13860;
 wire n_13861;
 wire n_13862;
 wire n_13863;
 wire n_13864;
 wire n_13865;
 wire n_13866;
 wire n_13867;
 wire n_13868;
 wire n_13869;
 wire n_1387;
 wire n_1388;
 wire n_13883;
 wire n_13884;
 wire n_1389;
 wire n_139;
 wire n_1390;
 wire n_1391;
 wire n_13919;
 wire n_1392;
 wire n_13920;
 wire n_1393;
 wire n_1394;
 wire n_13946;
 wire n_1395;
 wire n_1396;
 wire n_1397;
 wire n_13972;
 wire n_1398;
 wire n_13981;
 wire n_1399;
 wire n_14;
 wire n_140;
 wire n_1400;
 wire n_1401;
 wire n_14012;
 wire n_14014;
 wire n_14015;
 wire n_14017;
 wire n_14018;
 wire n_14019;
 wire n_1402;
 wire n_14020;
 wire n_14021;
 wire n_14022;
 wire n_14023;
 wire n_14024;
 wire n_14025;
 wire n_14026;
 wire n_14028;
 wire n_14029;
 wire n_1403;
 wire n_14030;
 wire n_14031;
 wire n_14032;
 wire n_14033;
 wire n_1404;
 wire n_1405;
 wire n_14054;
 wire n_14055;
 wire n_14056;
 wire n_14057;
 wire n_14058;
 wire n_14059;
 wire n_1406;
 wire n_14060;
 wire n_14061;
 wire n_14062;
 wire n_14063;
 wire n_14064;
 wire n_14065;
 wire n_14066;
 wire n_14067;
 wire n_14068;
 wire n_14069;
 wire n_1407;
 wire n_14070;
 wire n_14071;
 wire n_14072;
 wire n_14073;
 wire n_14074;
 wire n_14075;
 wire n_14076;
 wire n_14077;
 wire n_14078;
 wire n_14079;
 wire n_1408;
 wire n_14080;
 wire n_14081;
 wire n_14082;
 wire n_14085;
 wire n_14086;
 wire n_14087;
 wire n_14088;
 wire n_14089;
 wire n_1409;
 wire n_14090;
 wire n_14091;
 wire n_14092;
 wire n_14093;
 wire n_14094;
 wire n_14095;
 wire n_14096;
 wire n_14097;
 wire n_14098;
 wire n_14099;
 wire n_141;
 wire n_1410;
 wire n_14100;
 wire n_14101;
 wire n_14102;
 wire n_14103;
 wire n_14105;
 wire n_14106;
 wire n_14107;
 wire n_14108;
 wire n_14109;
 wire n_1411;
 wire n_14110;
 wire n_14111;
 wire n_14112;
 wire n_14113;
 wire n_14114;
 wire n_14115;
 wire n_14116;
 wire n_14117;
 wire n_14118;
 wire n_14119;
 wire n_1412;
 wire n_14120;
 wire n_14121;
 wire n_14123;
 wire n_14124;
 wire n_14125;
 wire n_14126;
 wire n_14127;
 wire n_14128;
 wire n_14129;
 wire n_1413;
 wire n_14130;
 wire n_14131;
 wire n_14132;
 wire n_14133;
 wire n_14134;
 wire n_14135;
 wire n_14136;
 wire n_14137;
 wire n_14139;
 wire n_14140;
 wire n_14141;
 wire n_14142;
 wire n_14143;
 wire n_14145;
 wire n_14146;
 wire n_14147;
 wire n_14148;
 wire n_14149;
 wire n_1415;
 wire n_14150;
 wire n_14151;
 wire n_14152;
 wire n_14153;
 wire n_14154;
 wire n_14155;
 wire n_14156;
 wire n_14157;
 wire n_14159;
 wire n_1416;
 wire n_14160;
 wire n_14161;
 wire n_14163;
 wire n_14164;
 wire n_14165;
 wire n_14166;
 wire n_14167;
 wire n_14168;
 wire n_14169;
 wire n_14170;
 wire n_14171;
 wire n_14172;
 wire n_14173;
 wire n_14174;
 wire n_14175;
 wire n_14176;
 wire n_14177;
 wire n_14178;
 wire n_14180;
 wire n_14181;
 wire n_14182;
 wire n_14183;
 wire n_14184;
 wire n_14185;
 wire n_14186;
 wire n_1419;
 wire n_14190;
 wire n_14191;
 wire n_14192;
 wire n_14193;
 wire n_14194;
 wire n_14196;
 wire n_14197;
 wire n_14199;
 wire n_142;
 wire n_1420;
 wire n_14200;
 wire n_14201;
 wire n_14203;
 wire n_14204;
 wire n_14205;
 wire n_14209;
 wire n_1421;
 wire n_14210;
 wire n_14212;
 wire n_14214;
 wire n_14215;
 wire n_14218;
 wire n_14219;
 wire n_1422;
 wire n_14220;
 wire n_14221;
 wire n_14222;
 wire n_14224;
 wire n_14225;
 wire n_14226;
 wire n_14228;
 wire n_14229;
 wire n_1423;
 wire n_14230;
 wire n_14231;
 wire n_14233;
 wire n_14234;
 wire n_14235;
 wire n_14236;
 wire n_14237;
 wire n_1424;
 wire n_14241;
 wire n_14243;
 wire n_14244;
 wire n_14245;
 wire n_14246;
 wire n_14247;
 wire n_14248;
 wire n_14249;
 wire n_1425;
 wire n_14250;
 wire n_14251;
 wire n_14252;
 wire n_14254;
 wire n_14255;
 wire n_14256;
 wire n_14257;
 wire n_14258;
 wire n_14259;
 wire n_1426;
 wire n_14261;
 wire n_14262;
 wire n_14263;
 wire n_14264;
 wire n_14266;
 wire n_14267;
 wire n_14268;
 wire n_14269;
 wire n_1427;
 wire n_14270;
 wire n_14271;
 wire n_14277;
 wire n_14278;
 wire n_14279;
 wire n_14280;
 wire n_14282;
 wire n_14283;
 wire n_14284;
 wire n_14285;
 wire n_14286;
 wire n_14287;
 wire n_14288;
 wire n_14289;
 wire n_1429;
 wire n_14290;
 wire n_14291;
 wire n_14292;
 wire n_14293;
 wire n_14294;
 wire n_14295;
 wire n_14296;
 wire n_14297;
 wire n_14298;
 wire n_14299;
 wire n_143;
 wire n_1430;
 wire n_14300;
 wire n_14301;
 wire n_14302;
 wire n_14303;
 wire n_14304;
 wire n_14305;
 wire n_14306;
 wire n_14307;
 wire n_14308;
 wire n_14309;
 wire n_1431;
 wire n_14310;
 wire n_14311;
 wire n_14312;
 wire n_14313;
 wire n_14314;
 wire n_14315;
 wire n_14316;
 wire n_14317;
 wire n_14318;
 wire n_14319;
 wire n_1432;
 wire n_14320;
 wire n_14321;
 wire n_14322;
 wire n_14323;
 wire n_14324;
 wire n_14325;
 wire n_14326;
 wire n_14327;
 wire n_14328;
 wire n_14329;
 wire n_1433;
 wire n_14330;
 wire n_14331;
 wire n_14332;
 wire n_14333;
 wire n_14334;
 wire n_14335;
 wire n_14336;
 wire n_14337;
 wire n_14338;
 wire n_14339;
 wire n_1434;
 wire n_14340;
 wire n_14341;
 wire n_14342;
 wire n_14343;
 wire n_14344;
 wire n_14345;
 wire n_14346;
 wire n_14347;
 wire n_14348;
 wire n_14349;
 wire n_1435;
 wire n_14350;
 wire n_14351;
 wire n_14352;
 wire n_14353;
 wire n_14354;
 wire n_14355;
 wire n_14356;
 wire n_14357;
 wire n_14358;
 wire n_14359;
 wire n_1436;
 wire n_14360;
 wire n_14361;
 wire n_14362;
 wire n_14363;
 wire n_14364;
 wire n_14365;
 wire n_14366;
 wire n_14367;
 wire n_14368;
 wire n_14369;
 wire n_1437;
 wire n_14370;
 wire n_14371;
 wire n_14372;
 wire n_14373;
 wire n_14374;
 wire n_14375;
 wire n_14376;
 wire n_14377;
 wire n_14378;
 wire n_14379;
 wire n_1438;
 wire n_14380;
 wire n_14381;
 wire n_14382;
 wire n_14383;
 wire n_14384;
 wire n_14385;
 wire n_14386;
 wire n_14387;
 wire n_14388;
 wire n_14389;
 wire n_1439;
 wire n_14390;
 wire n_14391;
 wire n_14392;
 wire n_14393;
 wire n_14394;
 wire n_14395;
 wire n_14396;
 wire n_14397;
 wire n_14398;
 wire n_14399;
 wire n_144;
 wire n_1440;
 wire n_14400;
 wire n_14401;
 wire n_14402;
 wire n_14403;
 wire n_14404;
 wire n_14405;
 wire n_14406;
 wire n_14407;
 wire n_14408;
 wire n_14409;
 wire n_1441;
 wire n_14410;
 wire n_14411;
 wire n_14412;
 wire n_14413;
 wire n_14414;
 wire n_14415;
 wire n_14416;
 wire n_14417;
 wire n_14418;
 wire n_14419;
 wire n_1442;
 wire n_14420;
 wire n_14421;
 wire n_14422;
 wire n_14423;
 wire n_14424;
 wire n_14425;
 wire n_14426;
 wire n_14427;
 wire n_14428;
 wire n_14429;
 wire n_1443;
 wire n_14430;
 wire n_14431;
 wire n_14432;
 wire n_14433;
 wire n_14434;
 wire n_14435;
 wire n_14436;
 wire n_14437;
 wire n_14438;
 wire n_14439;
 wire n_1444;
 wire n_14440;
 wire n_14441;
 wire n_14442;
 wire n_14443;
 wire n_14444;
 wire n_14445;
 wire n_14446;
 wire n_14447;
 wire n_14448;
 wire n_14449;
 wire n_1445;
 wire n_14450;
 wire n_14451;
 wire n_14452;
 wire n_14453;
 wire n_14454;
 wire n_14455;
 wire n_14456;
 wire n_14457;
 wire n_14458;
 wire n_14459;
 wire n_1446;
 wire n_14460;
 wire n_14461;
 wire n_14462;
 wire n_14463;
 wire n_14464;
 wire n_14465;
 wire n_14466;
 wire n_14467;
 wire n_14468;
 wire n_14469;
 wire n_1447;
 wire n_14471;
 wire n_14472;
 wire n_14473;
 wire n_14474;
 wire n_14475;
 wire n_14476;
 wire n_14477;
 wire n_14478;
 wire n_14479;
 wire n_1448;
 wire n_14480;
 wire n_14481;
 wire n_14482;
 wire n_14483;
 wire n_14484;
 wire n_14485;
 wire n_14486;
 wire n_14487;
 wire n_14488;
 wire n_14489;
 wire n_1449;
 wire n_14490;
 wire n_14491;
 wire n_14492;
 wire n_14493;
 wire n_14494;
 wire n_14495;
 wire n_14496;
 wire n_14497;
 wire n_14498;
 wire n_14499;
 wire n_145;
 wire n_1450;
 wire n_14500;
 wire n_14501;
 wire n_14502;
 wire n_14503;
 wire n_14504;
 wire n_14505;
 wire n_14506;
 wire n_14507;
 wire n_14508;
 wire n_14509;
 wire n_1451;
 wire n_14510;
 wire n_14511;
 wire n_14512;
 wire n_14513;
 wire n_14514;
 wire n_14515;
 wire n_14516;
 wire n_14517;
 wire n_14518;
 wire n_14519;
 wire n_1452;
 wire n_14520;
 wire n_14521;
 wire n_14522;
 wire n_14523;
 wire n_14524;
 wire n_14525;
 wire n_14526;
 wire n_14527;
 wire n_14528;
 wire n_14529;
 wire n_1453;
 wire n_14530;
 wire n_14531;
 wire n_14533;
 wire n_14534;
 wire n_14535;
 wire n_14536;
 wire n_1454;
 wire n_1455;
 wire n_1456;
 wire n_14564;
 wire n_1457;
 wire n_14575;
 wire n_1458;
 wire n_1459;
 wire n_1460;
 wire n_1461;
 wire n_1462;
 wire n_1463;
 wire n_1464;
 wire n_1465;
 wire n_1466;
 wire n_1467;
 wire n_1468;
 wire n_1469;
 wire n_147;
 wire n_1470;
 wire n_1471;
 wire n_1472;
 wire n_1473;
 wire n_1474;
 wire n_1475;
 wire n_1476;
 wire n_1477;
 wire n_1478;
 wire n_1479;
 wire n_148;
 wire n_1480;
 wire n_1481;
 wire n_1482;
 wire n_1483;
 wire n_1484;
 wire n_1485;
 wire n_1486;
 wire n_1487;
 wire n_1488;
 wire n_1489;
 wire n_149;
 wire n_1490;
 wire n_1491;
 wire n_1492;
 wire n_1493;
 wire n_1494;
 wire n_1495;
 wire n_1496;
 wire n_1497;
 wire n_1498;
 wire n_1499;
 wire n_15;
 wire n_150;
 wire n_1500;
 wire n_1501;
 wire n_1502;
 wire n_1503;
 wire n_1504;
 wire n_1505;
 wire n_1506;
 wire n_1507;
 wire n_1508;
 wire n_1509;
 wire n_151;
 wire n_1510;
 wire n_1511;
 wire n_1512;
 wire n_1513;
 wire n_1514;
 wire n_1515;
 wire n_1516;
 wire n_1517;
 wire n_1518;
 wire n_1519;
 wire n_152;
 wire n_1520;
 wire n_1521;
 wire n_1522;
 wire n_1523;
 wire n_1524;
 wire n_1525;
 wire n_1526;
 wire n_1527;
 wire n_1528;
 wire n_1529;
 wire n_1530;
 wire n_1531;
 wire n_1532;
 wire n_1533;
 wire n_1534;
 wire n_1535;
 wire n_1536;
 wire n_1537;
 wire n_1538;
 wire n_1539;
 wire n_154;
 wire n_1540;
 wire n_1541;
 wire n_1542;
 wire n_1543;
 wire n_1544;
 wire n_1545;
 wire n_1546;
 wire n_1547;
 wire n_1548;
 wire n_1549;
 wire n_155;
 wire n_1550;
 wire n_1551;
 wire n_1552;
 wire n_1553;
 wire n_1554;
 wire n_1555;
 wire n_1556;
 wire n_1557;
 wire n_1558;
 wire n_1559;
 wire n_156;
 wire n_1560;
 wire n_1561;
 wire n_1562;
 wire n_1563;
 wire n_1564;
 wire n_1565;
 wire n_1566;
 wire n_1567;
 wire n_1568;
 wire n_1569;
 wire n_15699_BAR;
 wire n_157;
 wire n_1570;
 wire n_1571;
 wire n_1572;
 wire n_1573;
 wire n_1574;
 wire n_1575;
 wire n_1576;
 wire n_1577;
 wire n_1578;
 wire n_1579;
 wire n_158;
 wire n_1580;
 wire n_1581;
 wire n_1582;
 wire n_1583;
 wire n_1584;
 wire n_1585;
 wire n_1586;
 wire n_1587;
 wire n_1588;
 wire n_1589;
 wire n_159;
 wire n_1590;
 wire n_1591;
 wire n_1592;
 wire n_1593;
 wire n_1594;
 wire n_1595;
 wire n_1596;
 wire n_1597;
 wire n_1598;
 wire n_1599;
 wire n_160;
 wire n_1600;
 wire n_1601;
 wire n_1602;
 wire n_1603;
 wire n_1604;
 wire n_1605;
 wire n_1606;
 wire n_1607;
 wire n_1608;
 wire n_1609;
 wire n_161;
 wire n_1610;
 wire n_1611;
 wire n_1612;
 wire n_1613;
 wire n_1614;
 wire n_1615;
 wire n_1616;
 wire n_1617;
 wire n_1618;
 wire n_1619;
 wire n_162;
 wire n_1620;
 wire n_1621;
 wire n_1622;
 wire n_1623;
 wire n_1624;
 wire n_1625;
 wire n_1626;
 wire n_1627;
 wire n_1628;
 wire n_1629;
 wire n_163;
 wire n_1630;
 wire n_1631;
 wire n_1632;
 wire n_1633;
 wire n_1634;
 wire n_1635;
 wire n_1636;
 wire n_1637;
 wire n_1638;
 wire n_1639;
 wire n_164;
 wire n_1640;
 wire n_1641;
 wire n_1643;
 wire n_1644;
 wire n_1645;
 wire n_1646;
 wire n_1647;
 wire n_1648;
 wire n_1649;
 wire n_165;
 wire n_1650;
 wire n_1651;
 wire n_1652;
 wire n_1653;
 wire n_1654;
 wire n_1655;
 wire n_1657;
 wire n_1658;
 wire n_1659;
 wire n_166;
 wire n_1660;
 wire n_1661;
 wire n_1662;
 wire n_1663;
 wire n_1664;
 wire n_1665;
 wire n_1666;
 wire n_1667;
 wire n_1668;
 wire n_1669;
 wire n_167;
 wire n_1670;
 wire n_1671;
 wire n_1672;
 wire n_1673;
 wire n_1674;
 wire n_1675;
 wire n_1676;
 wire n_1677;
 wire n_1678;
 wire n_1679;
 wire n_168;
 wire n_1680;
 wire n_1681;
 wire n_1682;
 wire n_1683;
 wire n_1684;
 wire n_1685;
 wire n_1686;
 wire n_1688;
 wire n_1689;
 wire n_169;
 wire n_1690;
 wire n_1691;
 wire n_1692;
 wire n_1693;
 wire n_1694;
 wire n_1695;
 wire n_1696;
 wire n_1697;
 wire n_1698;
 wire n_1699;
 wire n_17;
 wire n_170;
 wire n_1700;
 wire n_1701;
 wire n_1702;
 wire n_1703;
 wire n_1704;
 wire n_1705;
 wire n_1706;
 wire n_1707;
 wire n_1708;
 wire n_1709;
 wire n_171;
 wire n_1710;
 wire n_1711;
 wire n_1712;
 wire n_1713;
 wire n_1714;
 wire n_1715;
 wire n_1716;
 wire n_1717;
 wire n_1718;
 wire n_1719;
 wire n_172;
 wire n_1720;
 wire n_1721;
 wire n_1722;
 wire n_1723;
 wire n_1724;
 wire n_1725;
 wire n_1726;
 wire n_1727;
 wire n_1728;
 wire n_1729;
 wire n_173;
 wire n_1730;
 wire n_1731;
 wire n_1732;
 wire n_1733;
 wire n_1734;
 wire n_1735;
 wire n_1736;
 wire n_1737;
 wire n_1738;
 wire n_1739;
 wire n_174;
 wire n_1740;
 wire n_1741;
 wire n_1742;
 wire n_1743;
 wire n_1744;
 wire n_1745;
 wire n_1746;
 wire n_1747;
 wire n_1748;
 wire n_1749;
 wire n_175;
 wire n_1750;
 wire n_1751;
 wire n_1752;
 wire n_1753;
 wire n_1754;
 wire n_1755;
 wire n_1756;
 wire n_1757;
 wire n_1758;
 wire n_1759;
 wire n_176;
 wire n_1760;
 wire n_1761;
 wire n_1762;
 wire n_1763;
 wire n_1764;
 wire n_1765;
 wire n_1766;
 wire n_1767;
 wire n_1768;
 wire n_1769;
 wire n_177;
 wire n_1770;
 wire n_1771;
 wire n_1772;
 wire n_1773;
 wire n_1774;
 wire n_1775;
 wire n_1776;
 wire n_1777;
 wire n_1778;
 wire n_1779;
 wire n_178;
 wire n_1780;
 wire n_1781;
 wire n_1782;
 wire n_1783;
 wire n_1784;
 wire n_1785;
 wire n_1786;
 wire n_1787;
 wire n_1788;
 wire n_1789;
 wire n_179;
 wire n_1790;
 wire n_1791;
 wire n_1792;
 wire n_1793;
 wire n_1794;
 wire n_1795;
 wire n_1796;
 wire n_1797;
 wire n_1798;
 wire n_1799;
 wire n_180;
 wire n_1800;
 wire n_1801;
 wire n_1802;
 wire n_1803;
 wire n_1804;
 wire n_1805;
 wire n_1806;
 wire n_1807;
 wire n_1808;
 wire n_1809;
 wire n_181;
 wire n_1810;
 wire n_1811;
 wire n_1812;
 wire n_1813;
 wire n_1814;
 wire n_1815;
 wire n_1816;
 wire n_1817;
 wire n_1818;
 wire n_1819;
 wire n_182;
 wire n_1820;
 wire n_1821;
 wire n_1822;
 wire n_1823;
 wire n_1824;
 wire n_1825;
 wire n_1826;
 wire n_1827;
 wire n_1828;
 wire n_1829;
 wire n_183;
 wire n_1830;
 wire n_1831;
 wire n_1832;
 wire n_1833;
 wire n_1834;
 wire n_1835;
 wire n_1836;
 wire n_1837;
 wire n_1838;
 wire n_1839;
 wire n_184;
 wire n_1840;
 wire n_1841;
 wire n_1842;
 wire n_1843;
 wire n_1844;
 wire n_1845;
 wire n_1846;
 wire n_1847;
 wire n_1849;
 wire n_185;
 wire n_1850;
 wire n_1851;
 wire n_1852;
 wire n_1853;
 wire n_1854;
 wire n_1855;
 wire n_186;
 wire n_1860;
 wire n_1861;
 wire n_1863;
 wire n_1865;
 wire n_1866;
 wire n_1867;
 wire n_187;
 wire n_1871;
 wire n_1873;
 wire n_1875;
 wire n_1877;
 wire n_1879;
 wire n_188;
 wire n_1883;
 wire n_1884;
 wire n_1889;
 wire n_189;
 wire n_1891;
 wire n_1895;
 wire n_1896;
 wire n_190;
 wire n_1900;
 wire n_1903;
 wire n_191;
 wire n_1910;
 wire n_1911;
 wire n_1912;
 wire n_1913;
 wire n_1914;
 wire n_1915;
 wire n_1916;
 wire n_1917;
 wire n_1918;
 wire n_1919;
 wire n_192;
 wire n_1920;
 wire n_1922;
 wire n_1923;
 wire n_1925;
 wire n_193;
 wire n_1930;
 wire n_1931;
 wire n_1932;
 wire n_1933;
 wire n_1934;
 wire n_1935;
 wire n_1936;
 wire n_1937;
 wire n_1939;
 wire n_194;
 wire n_1940;
 wire n_1942;
 wire n_1943;
 wire n_1944;
 wire n_1945;
 wire n_1949;
 wire n_195;
 wire n_1950;
 wire n_1951;
 wire n_1952;
 wire n_1954;
 wire n_1955;
 wire n_1956;
 wire n_1957;
 wire n_196;
 wire n_1960;
 wire n_1961;
 wire n_1962;
 wire n_1963;
 wire n_1964;
 wire n_1965;
 wire n_1966;
 wire n_1967;
 wire n_1968;
 wire n_1969;
 wire n_197;
 wire n_1970;
 wire n_1971;
 wire n_1972;
 wire n_1974;
 wire n_1975;
 wire n_1976;
 wire n_1977;
 wire n_1978;
 wire n_1979;
 wire n_198;
 wire n_1980;
 wire n_1981;
 wire n_1982;
 wire n_1983;
 wire n_1984;
 wire n_1985;
 wire n_1986;
 wire n_1988;
 wire n_1989;
 wire n_199;
 wire n_1990;
 wire n_1991;
 wire n_1992;
 wire n_1993;
 wire n_1994;
 wire n_1995;
 wire n_1996;
 wire n_1997;
 wire n_1998;
 wire n_1999;
 wire n_2;
 wire n_20;
 wire n_200;
 wire n_2000;
 wire n_2001;
 wire n_2002;
 wire n_2003;
 wire n_2004;
 wire n_2005;
 wire n_2006;
 wire n_2007;
 wire n_2008;
 wire n_2009;
 wire n_201;
 wire n_2010;
 wire n_2011;
 wire n_2012;
 wire n_2013;
 wire n_2014;
 wire n_2015;
 wire n_2016;
 wire n_2017;
 wire n_2019;
 wire n_202;
 wire n_2020;
 wire n_2021;
 wire n_2022;
 wire n_2023;
 wire n_2024;
 wire n_2025;
 wire n_2026;
 wire n_2027;
 wire n_203;
 wire n_204;
 wire n_2043;
 wire n_205;
 wire n_2053;
 wire n_2054;
 wire n_2055;
 wire n_2056;
 wire n_2057;
 wire n_2058;
 wire n_2059;
 wire n_206;
 wire n_2060;
 wire n_2061;
 wire n_2062;
 wire n_2063;
 wire n_2064;
 wire n_2065;
 wire n_2066;
 wire n_2067;
 wire n_2068;
 wire n_2069;
 wire n_207;
 wire n_2070;
 wire n_2071;
 wire n_2072;
 wire n_2073;
 wire n_2074;
 wire n_2075;
 wire n_2076;
 wire n_2077;
 wire n_2078;
 wire n_2079;
 wire n_208;
 wire n_2080;
 wire n_2081;
 wire n_2082;
 wire n_2083;
 wire n_2084;
 wire n_2085;
 wire n_2086;
 wire n_2087;
 wire n_2088;
 wire n_2089;
 wire n_209;
 wire n_2090;
 wire n_2091;
 wire n_2092;
 wire n_2093;
 wire n_2094;
 wire n_2095;
 wire n_2096;
 wire n_2097;
 wire n_2098;
 wire n_2099;
 wire n_210;
 wire n_2100;
 wire n_2101;
 wire n_2102;
 wire n_2103;
 wire n_2104;
 wire n_2105;
 wire n_2106;
 wire n_2107;
 wire n_2108;
 wire n_2109;
 wire n_211;
 wire n_2110;
 wire n_2111;
 wire n_2112;
 wire n_2113;
 wire n_2114;
 wire n_2115;
 wire n_2116;
 wire n_2117;
 wire n_2118;
 wire n_2119;
 wire n_212;
 wire n_2120;
 wire n_2121;
 wire n_2122;
 wire n_2123;
 wire n_2124;
 wire n_2125;
 wire n_2126;
 wire n_2127;
 wire n_2128;
 wire n_2129;
 wire n_213;
 wire n_2130;
 wire n_2131;
 wire n_2132;
 wire n_2133;
 wire n_2134;
 wire n_2135;
 wire n_2136;
 wire n_2137;
 wire n_2138;
 wire n_2139;
 wire n_214;
 wire n_2140;
 wire n_2141;
 wire n_2142;
 wire n_2143;
 wire n_2144;
 wire n_2145;
 wire n_2146;
 wire n_2147;
 wire n_2148;
 wire n_2149;
 wire n_215;
 wire n_2150;
 wire n_2151;
 wire n_2152;
 wire n_2153;
 wire n_2154;
 wire n_2155;
 wire n_2156;
 wire n_2157;
 wire n_2158;
 wire n_2159;
 wire n_216;
 wire n_2160;
 wire n_2161;
 wire n_2162;
 wire n_2163;
 wire n_2164;
 wire n_2165;
 wire n_2166;
 wire n_2167;
 wire n_2168;
 wire n_2169;
 wire n_217;
 wire n_2170;
 wire n_2171;
 wire n_2173;
 wire n_2174;
 wire n_2175;
 wire n_2176;
 wire n_2177;
 wire n_2178;
 wire n_2179;
 wire n_218;
 wire n_2180;
 wire n_2181;
 wire n_2182;
 wire n_2183;
 wire n_2184;
 wire n_2185;
 wire n_2186;
 wire n_2187;
 wire n_2188;
 wire n_2189;
 wire n_219;
 wire n_2190;
 wire n_2191;
 wire n_2192;
 wire n_2193;
 wire n_2194;
 wire n_2195;
 wire n_2196;
 wire n_2197;
 wire n_2198;
 wire n_2199;
 wire n_22;
 wire n_220;
 wire n_2200;
 wire n_2201;
 wire n_2202;
 wire n_2203;
 wire n_2204;
 wire n_2205;
 wire n_2206;
 wire n_2207;
 wire n_2208;
 wire n_2209;
 wire n_221;
 wire n_2210;
 wire n_2211;
 wire n_2212;
 wire n_2213;
 wire n_2214;
 wire n_2215;
 wire n_2216;
 wire n_2217;
 wire n_2218;
 wire n_2219;
 wire n_222;
 wire n_2220;
 wire n_2221;
 wire n_2222;
 wire n_2223;
 wire n_2224;
 wire n_2225;
 wire n_2226;
 wire n_2227;
 wire n_2228;
 wire n_2229;
 wire n_223;
 wire n_2230;
 wire n_2231;
 wire n_2232;
 wire n_2233;
 wire n_2234;
 wire n_2235;
 wire n_2236;
 wire n_2237;
 wire n_2238;
 wire n_2239;
 wire n_224;
 wire n_2240;
 wire n_2241;
 wire n_2242;
 wire n_2243;
 wire n_2244;
 wire n_2245;
 wire n_2246;
 wire n_2247;
 wire n_2248;
 wire n_2249;
 wire n_225;
 wire n_2250;
 wire n_2251;
 wire n_2252;
 wire n_2253;
 wire n_2254;
 wire n_2255;
 wire n_2256;
 wire n_2257;
 wire n_2258;
 wire n_2259;
 wire n_226;
 wire n_2260;
 wire n_2261;
 wire n_2262;
 wire n_2263;
 wire n_2264;
 wire n_2265;
 wire n_2266;
 wire n_2267;
 wire n_2268;
 wire n_2269;
 wire n_227;
 wire n_2270;
 wire n_2271;
 wire n_2272;
 wire n_2273;
 wire n_2274;
 wire n_2275;
 wire n_2276;
 wire n_2277;
 wire n_2278;
 wire n_2279;
 wire n_228;
 wire n_2280;
 wire n_2281;
 wire n_2282;
 wire n_2283;
 wire n_2284;
 wire n_2285;
 wire n_2286;
 wire n_2287;
 wire n_2288;
 wire n_2289;
 wire n_229;
 wire n_2290;
 wire n_2291;
 wire n_2292;
 wire n_2293;
 wire n_2294;
 wire n_2295;
 wire n_2296;
 wire n_2297;
 wire n_2298;
 wire n_2299;
 wire n_23;
 wire n_230;
 wire n_2300;
 wire n_2301;
 wire n_2302;
 wire n_2303;
 wire n_2304;
 wire n_2305;
 wire n_2306;
 wire n_2307;
 wire n_2308;
 wire n_2309;
 wire n_231;
 wire n_2310;
 wire n_2311;
 wire n_2312;
 wire n_2313;
 wire n_2314;
 wire n_2315;
 wire n_2316;
 wire n_2317;
 wire n_2318;
 wire n_2319;
 wire n_232;
 wire n_2320;
 wire n_2321;
 wire n_2322;
 wire n_2323;
 wire n_2324;
 wire n_2325;
 wire n_2326;
 wire n_2327;
 wire n_2328;
 wire n_2329;
 wire n_233;
 wire n_2330;
 wire n_2331;
 wire n_2332;
 wire n_2333;
 wire n_2334;
 wire n_2335;
 wire n_2336;
 wire n_2337;
 wire n_2338;
 wire n_2339;
 wire n_234;
 wire n_2340;
 wire n_2341;
 wire n_2342;
 wire n_2343;
 wire n_2344;
 wire n_2345;
 wire n_2346;
 wire n_2347;
 wire n_2348;
 wire n_2349;
 wire n_235;
 wire n_2350;
 wire n_2351;
 wire n_2352;
 wire n_2353;
 wire n_2354;
 wire n_2355;
 wire n_2356;
 wire n_2357;
 wire n_2358;
 wire n_2359;
 wire n_236;
 wire n_2360;
 wire n_2361;
 wire n_2362;
 wire n_2363;
 wire n_2364;
 wire n_2365;
 wire n_2367;
 wire n_2368;
 wire n_2369;
 wire n_237;
 wire n_2370;
 wire n_2371;
 wire n_2372;
 wire n_2373;
 wire n_2374;
 wire n_2375;
 wire n_2376;
 wire n_2377;
 wire n_2378;
 wire n_2379;
 wire n_238;
 wire n_2380;
 wire n_2381;
 wire n_2382;
 wire n_2383;
 wire n_2384;
 wire n_2385;
 wire n_2386;
 wire n_2387;
 wire n_2388;
 wire n_2389;
 wire n_239;
 wire n_2390;
 wire n_2391;
 wire n_2392;
 wire n_2393;
 wire n_2394;
 wire n_2395;
 wire n_2396;
 wire n_2397;
 wire n_2398;
 wire n_2399;
 wire n_24;
 wire n_240;
 wire n_2400;
 wire n_2401;
 wire n_2402;
 wire n_2403;
 wire n_2404;
 wire n_2405;
 wire n_2406;
 wire n_2407;
 wire n_2408;
 wire n_2409;
 wire n_241;
 wire n_2410;
 wire n_2411;
 wire n_2412;
 wire n_2413;
 wire n_2414;
 wire n_2415;
 wire n_2416;
 wire n_2417;
 wire n_2418;
 wire n_2419;
 wire n_242;
 wire n_2420;
 wire n_2421;
 wire n_2422;
 wire n_2423;
 wire n_2424;
 wire n_2425;
 wire n_2426;
 wire n_2427;
 wire n_2428;
 wire n_2429;
 wire n_243;
 wire n_2430;
 wire n_2431;
 wire n_2432;
 wire n_2433;
 wire n_2434;
 wire n_2435;
 wire n_2436;
 wire n_2437;
 wire n_2438;
 wire n_2439;
 wire n_244;
 wire n_2440;
 wire n_2441;
 wire n_2442;
 wire n_2443;
 wire n_2444;
 wire n_2445;
 wire n_2446;
 wire n_2447;
 wire n_2448;
 wire n_2449;
 wire n_245;
 wire n_2450;
 wire n_2451;
 wire n_2452;
 wire n_2453;
 wire n_2454;
 wire n_2455;
 wire n_2456;
 wire n_2457;
 wire n_2458;
 wire n_2459;
 wire n_246;
 wire n_2460;
 wire n_2461;
 wire n_2462;
 wire n_2463;
 wire n_2464;
 wire n_2465;
 wire n_2466;
 wire n_2467;
 wire n_2468;
 wire n_2469;
 wire n_247;
 wire n_2470;
 wire n_2471;
 wire n_2472;
 wire n_2473;
 wire n_2474;
 wire n_2475;
 wire n_2476;
 wire n_2477;
 wire n_2478;
 wire n_2479;
 wire n_248;
 wire n_2480;
 wire n_2481;
 wire n_2482;
 wire n_2483;
 wire n_2484;
 wire n_2485;
 wire n_2486;
 wire n_2487;
 wire n_2488;
 wire n_2489;
 wire n_2490;
 wire n_2491;
 wire n_2492;
 wire n_2493;
 wire n_2494;
 wire n_2495;
 wire n_2496;
 wire n_2497;
 wire n_2498;
 wire n_2499;
 wire n_25;
 wire n_250;
 wire n_2500;
 wire n_2501;
 wire n_2502;
 wire n_2503;
 wire n_2504;
 wire n_2505;
 wire n_2506;
 wire n_2507;
 wire n_2508;
 wire n_2509;
 wire n_251;
 wire n_2510;
 wire n_2511;
 wire n_2512;
 wire n_2513;
 wire n_2514;
 wire n_2515;
 wire n_2516;
 wire n_2517;
 wire n_2518;
 wire n_2519;
 wire n_252;
 wire n_2520;
 wire n_2521;
 wire n_2522;
 wire n_2523;
 wire n_2524;
 wire n_2525;
 wire n_2526;
 wire n_2527;
 wire n_2528;
 wire n_2529;
 wire n_253;
 wire n_2530;
 wire n_2531;
 wire n_2532;
 wire n_2533;
 wire n_2534;
 wire n_2535;
 wire n_2536;
 wire n_2537;
 wire n_2538;
 wire n_2539;
 wire n_254;
 wire n_2540;
 wire n_2541;
 wire n_2542;
 wire n_2543;
 wire n_2544;
 wire n_2545;
 wire n_2546;
 wire n_2547;
 wire n_2548;
 wire n_2549;
 wire n_255;
 wire n_2550;
 wire n_2551;
 wire n_2552;
 wire n_2553;
 wire n_2554;
 wire n_2555;
 wire n_2556;
 wire n_2557;
 wire n_2558;
 wire n_2559;
 wire n_256;
 wire n_2560;
 wire n_2561;
 wire n_2562;
 wire n_2563;
 wire n_2564;
 wire n_2565;
 wire n_2566;
 wire n_2567;
 wire n_2568;
 wire n_2569;
 wire n_257;
 wire n_2570;
 wire n_2571;
 wire n_2572;
 wire n_2573;
 wire n_2574;
 wire n_2575;
 wire n_2576;
 wire n_2577;
 wire n_2578;
 wire n_2579;
 wire n_258;
 wire n_2580;
 wire n_2581;
 wire n_2582;
 wire n_2583;
 wire n_2584;
 wire n_2585;
 wire n_2586;
 wire n_2587;
 wire n_2588;
 wire n_2589;
 wire n_259;
 wire n_2590;
 wire n_2591;
 wire n_2592;
 wire n_2593;
 wire n_2594;
 wire n_2595;
 wire n_2596;
 wire n_2597;
 wire n_2598;
 wire n_2599;
 wire n_26;
 wire n_260;
 wire n_2600;
 wire n_2601;
 wire n_2602;
 wire n_2603;
 wire n_2604;
 wire n_2605;
 wire n_2606;
 wire n_2607;
 wire n_2608;
 wire n_2609;
 wire n_261;
 wire n_2610;
 wire n_2611;
 wire n_2612;
 wire n_2613;
 wire n_2614;
 wire n_2615;
 wire n_2616;
 wire n_2617;
 wire n_2618;
 wire n_2619;
 wire n_262;
 wire n_2620;
 wire n_2621;
 wire n_2622;
 wire n_2623;
 wire n_2624;
 wire n_2625;
 wire n_2626;
 wire n_2627;
 wire n_2628;
 wire n_2629;
 wire n_263;
 wire n_2630;
 wire n_2631;
 wire n_2632;
 wire n_2633;
 wire n_2634;
 wire n_2635;
 wire n_2636;
 wire n_2637;
 wire n_2638;
 wire n_2639;
 wire n_264;
 wire n_2640;
 wire n_2641;
 wire n_2642;
 wire n_2643;
 wire n_2644;
 wire n_2645;
 wire n_2646;
 wire n_2647;
 wire n_2648;
 wire n_2649;
 wire n_265;
 wire n_2650;
 wire n_2651;
 wire n_2652;
 wire n_2653;
 wire n_2654;
 wire n_2655;
 wire n_2656;
 wire n_2657;
 wire n_2658;
 wire n_2659;
 wire n_266;
 wire n_2660;
 wire n_2661;
 wire n_2662;
 wire n_2663;
 wire n_2664;
 wire n_2665;
 wire n_2666;
 wire n_2667;
 wire n_2668;
 wire n_2669;
 wire n_267;
 wire n_2670;
 wire n_2671;
 wire n_2672;
 wire n_2673;
 wire n_2674;
 wire n_2675;
 wire n_2676;
 wire n_2677;
 wire n_2678;
 wire n_2679;
 wire n_268;
 wire n_2680;
 wire n_2681;
 wire n_2682;
 wire n_2683;
 wire n_2684;
 wire n_2685;
 wire n_2686;
 wire n_2687;
 wire n_2688;
 wire n_2689;
 wire n_269;
 wire n_2690;
 wire n_2691;
 wire n_2692;
 wire n_2693;
 wire n_2694;
 wire n_2695;
 wire n_2696;
 wire n_2697;
 wire n_2698;
 wire n_2699;
 wire n_27;
 wire n_270;
 wire n_2700;
 wire n_2701;
 wire n_2702;
 wire n_2703;
 wire n_2704;
 wire n_2705;
 wire n_2706;
 wire n_2707;
 wire n_2708;
 wire n_2709;
 wire n_271;
 wire n_2710;
 wire n_2711;
 wire n_2712;
 wire n_2713;
 wire n_2714;
 wire n_2715;
 wire n_2716;
 wire n_2717;
 wire n_2718;
 wire n_2719;
 wire n_272;
 wire n_2720;
 wire n_2721;
 wire n_2722;
 wire n_2723;
 wire n_2724;
 wire n_2725;
 wire n_2726;
 wire n_2727;
 wire n_2728;
 wire n_2729;
 wire n_273;
 wire n_2730;
 wire n_2731;
 wire n_2732;
 wire n_2733;
 wire n_2734;
 wire n_2735;
 wire n_2736;
 wire n_2737;
 wire n_2738;
 wire n_2739;
 wire n_274;
 wire n_2740;
 wire n_2741;
 wire n_2742;
 wire n_2743;
 wire n_2744;
 wire n_2745;
 wire n_2746;
 wire n_2747;
 wire n_2748;
 wire n_2749;
 wire n_275;
 wire n_2750;
 wire n_2751;
 wire n_2752;
 wire n_2753;
 wire n_2754;
 wire n_2755;
 wire n_2756;
 wire n_2757;
 wire n_2758;
 wire n_2759;
 wire n_276;
 wire n_2760;
 wire n_2761;
 wire n_2762;
 wire n_2763;
 wire n_2764;
 wire n_2765;
 wire n_2766;
 wire n_2767;
 wire n_2768;
 wire n_2769;
 wire n_277;
 wire n_2770;
 wire n_2771;
 wire n_2772;
 wire n_2773;
 wire n_2774;
 wire n_2775;
 wire n_2776;
 wire n_2777;
 wire n_2778;
 wire n_2779;
 wire n_278;
 wire n_2780;
 wire n_2781;
 wire n_2782;
 wire n_2783;
 wire n_2784;
 wire n_2785;
 wire n_2786;
 wire n_2787;
 wire n_2788;
 wire n_2789;
 wire n_279;
 wire n_2790;
 wire n_2791;
 wire n_2792;
 wire n_2793;
 wire n_2794;
 wire n_2795;
 wire n_2796;
 wire n_2797;
 wire n_2798;
 wire n_2799;
 wire n_28;
 wire n_280;
 wire n_2800;
 wire n_2801;
 wire n_2802;
 wire n_2803;
 wire n_2804;
 wire n_2805;
 wire n_2806;
 wire n_2807;
 wire n_2808;
 wire n_2809;
 wire n_281;
 wire n_2810;
 wire n_2811;
 wire n_2812;
 wire n_2813;
 wire n_2814;
 wire n_2815;
 wire n_2816;
 wire n_2817;
 wire n_2818;
 wire n_2819;
 wire n_282;
 wire n_2820;
 wire n_2821;
 wire n_2822;
 wire n_2823;
 wire n_2824;
 wire n_2825;
 wire n_2826;
 wire n_2827;
 wire n_2828;
 wire n_2829;
 wire n_283;
 wire n_2830;
 wire n_2831;
 wire n_2832;
 wire n_2833;
 wire n_2834;
 wire n_2835;
 wire n_2836;
 wire n_2837;
 wire n_2838;
 wire n_2839;
 wire n_284;
 wire n_2840;
 wire n_2841;
 wire n_2842;
 wire n_2843;
 wire n_2844;
 wire n_2845;
 wire n_2846;
 wire n_2847;
 wire n_2848;
 wire n_2849;
 wire n_285;
 wire n_2850;
 wire n_2851;
 wire n_2852;
 wire n_2853;
 wire n_2854;
 wire n_2855;
 wire n_2856;
 wire n_2857;
 wire n_2858;
 wire n_2859;
 wire n_286;
 wire n_2860;
 wire n_2861;
 wire n_2862;
 wire n_2863;
 wire n_2864;
 wire n_2865;
 wire n_2866;
 wire n_2867;
 wire n_2868;
 wire n_2869;
 wire n_287;
 wire n_2870;
 wire n_2871;
 wire n_2872;
 wire n_2873;
 wire n_2874;
 wire n_2875;
 wire n_2877;
 wire n_2878;
 wire n_2879;
 wire n_288;
 wire n_2880;
 wire n_2882;
 wire n_2887;
 wire n_2888;
 wire n_289;
 wire n_2896;
 wire n_29;
 wire n_290;
 wire n_2907;
 wire n_2908;
 wire n_291;
 wire n_292;
 wire n_2928;
 wire n_2929;
 wire n_293;
 wire n_2930;
 wire n_2931;
 wire n_2932;
 wire n_2934;
 wire n_2935;
 wire n_2936;
 wire n_2937;
 wire n_2938;
 wire n_2939;
 wire n_294;
 wire n_2940;
 wire n_2941;
 wire n_2942;
 wire n_2943;
 wire n_2944;
 wire n_2945;
 wire n_2946;
 wire n_2947;
 wire n_2948;
 wire n_2949;
 wire n_295;
 wire n_2950;
 wire n_2951;
 wire n_2952;
 wire n_2953;
 wire n_2957;
 wire n_2958;
 wire n_2959;
 wire n_296;
 wire n_2960;
 wire n_2961;
 wire n_2962;
 wire n_2963;
 wire n_2964;
 wire n_297;
 wire n_2971;
 wire n_2972;
 wire n_2973;
 wire n_2974;
 wire n_2975;
 wire n_2976;
 wire n_2977;
 wire n_2978;
 wire n_2979;
 wire n_298;
 wire n_2980;
 wire n_2982;
 wire n_2983;
 wire n_2984;
 wire n_2986;
 wire n_2987;
 wire n_2988;
 wire n_2989;
 wire n_299;
 wire n_2990;
 wire n_2991;
 wire n_2992;
 wire n_2993;
 wire n_2994;
 wire n_2995;
 wire n_2996;
 wire n_2997;
 wire n_2998;
 wire n_2999;
 wire n_3;
 wire n_30;
 wire n_300;
 wire n_3000;
 wire n_3001;
 wire n_3002;
 wire n_3003;
 wire n_3005;
 wire n_3007;
 wire n_3008;
 wire n_3009;
 wire n_301;
 wire n_3010;
 wire n_3011;
 wire n_3012;
 wire n_3014;
 wire n_3016;
 wire n_3017;
 wire n_3018;
 wire n_3019;
 wire n_302;
 wire n_3020;
 wire n_3021;
 wire n_3022;
 wire n_3023;
 wire n_3024;
 wire n_3025;
 wire n_3026;
 wire n_3027;
 wire n_3028;
 wire n_3029;
 wire n_303;
 wire n_3030;
 wire n_3031;
 wire n_3034;
 wire n_3035;
 wire n_3037;
 wire n_3039;
 wire n_304;
 wire n_3040;
 wire n_3041;
 wire n_3042;
 wire n_3043;
 wire n_3045;
 wire n_3047;
 wire n_3049;
 wire n_305;
 wire n_3052;
 wire n_3053;
 wire n_3054;
 wire n_3055;
 wire n_3057;
 wire n_3058;
 wire n_3059;
 wire n_306;
 wire n_3060;
 wire n_3061;
 wire n_3062;
 wire n_3063;
 wire n_3064;
 wire n_3065;
 wire n_3066;
 wire n_3067;
 wire n_3068;
 wire n_3069;
 wire n_307;
 wire n_3070;
 wire n_3071;
 wire n_3074;
 wire n_3077;
 wire n_3078;
 wire n_3079;
 wire n_3080;
 wire n_3081;
 wire n_3082;
 wire n_3083;
 wire n_3084;
 wire n_3086;
 wire n_3087;
 wire n_3088;
 wire n_3089;
 wire n_309;
 wire n_3090;
 wire n_3091;
 wire n_3092;
 wire n_3093;
 wire n_3094;
 wire n_3095;
 wire n_3096;
 wire n_3097;
 wire n_3098;
 wire n_3099;
 wire n_31;
 wire n_310;
 wire n_3100;
 wire n_3101;
 wire n_3102;
 wire n_3103;
 wire n_3104;
 wire n_3105;
 wire n_3106;
 wire n_3107;
 wire n_3108;
 wire n_3109;
 wire n_3110;
 wire n_3111;
 wire n_3112;
 wire n_3113;
 wire n_3114;
 wire n_3115;
 wire n_3116;
 wire n_3117;
 wire n_3118;
 wire n_3119;
 wire n_312;
 wire n_3120;
 wire n_3121;
 wire n_3122;
 wire n_3123;
 wire n_3124;
 wire n_3125;
 wire n_3126;
 wire n_3127;
 wire n_3128;
 wire n_3129;
 wire n_313;
 wire n_3130;
 wire n_3132;
 wire n_3133;
 wire n_3135;
 wire n_3136;
 wire n_3137;
 wire n_3138;
 wire n_3139;
 wire n_314;
 wire n_3140;
 wire n_3141;
 wire n_3142;
 wire n_3143;
 wire n_3144;
 wire n_3145;
 wire n_3146;
 wire n_3147;
 wire n_3148;
 wire n_3149;
 wire n_315;
 wire n_3150;
 wire n_3151;
 wire n_3152;
 wire n_3153;
 wire n_3154;
 wire n_3155;
 wire n_3156;
 wire n_3157;
 wire n_3158;
 wire n_3159;
 wire n_316;
 wire n_3160;
 wire n_3161;
 wire n_3162;
 wire n_3163;
 wire n_3164;
 wire n_3165;
 wire n_3166;
 wire n_3167;
 wire n_3168;
 wire n_3169;
 wire n_317;
 wire n_3170;
 wire n_3171;
 wire n_3172;
 wire n_3173;
 wire n_3174;
 wire n_3175;
 wire n_3176;
 wire n_3177;
 wire n_3178;
 wire n_3179;
 wire n_318;
 wire n_3180;
 wire n_3181;
 wire n_3182;
 wire n_3183;
 wire n_3184;
 wire n_3185;
 wire n_3186;
 wire n_3187;
 wire n_3188;
 wire n_3189;
 wire n_319;
 wire n_3190;
 wire n_3191;
 wire n_3192;
 wire n_3193;
 wire n_3194;
 wire n_3196;
 wire n_3198;
 wire n_3199;
 wire n_32;
 wire n_320;
 wire n_3200;
 wire n_3201;
 wire n_3202;
 wire n_3203;
 wire n_3204;
 wire n_3206;
 wire n_3207;
 wire n_3208;
 wire n_3209;
 wire n_321;
 wire n_3210;
 wire n_3212;
 wire n_3213;
 wire n_3214;
 wire n_3215;
 wire n_3216;
 wire n_3217;
 wire n_3218;
 wire n_3219;
 wire n_322;
 wire n_3220;
 wire n_3221;
 wire n_3222;
 wire n_323;
 wire n_324;
 wire n_325;
 wire n_326;
 wire n_327;
 wire n_328;
 wire n_3287;
 wire n_329;
 wire n_3292;
 wire n_3294;
 wire n_3297;
 wire n_3299;
 wire n_33;
 wire n_330;
 wire n_3302;
 wire n_3303;
 wire n_3305;
 wire n_3306;
 wire n_331;
 wire n_3310;
 wire n_3311;
 wire n_332;
 wire n_333;
 wire n_3336;
 wire n_3337;
 wire n_334;
 wire n_3341;
 wire n_3344;
 wire n_3345;
 wire n_3347;
 wire n_3348;
 wire n_3349;
 wire n_335;
 wire n_3350;
 wire n_3351;
 wire n_3353;
 wire n_3354;
 wire n_3355;
 wire n_3358;
 wire n_336;
 wire n_337;
 wire n_3386;
 wire n_339;
 wire n_3395;
 wire n_34;
 wire n_340;
 wire n_3401;
 wire n_3409;
 wire n_341;
 wire n_3411;
 wire n_3415;
 wire n_342;
 wire n_3427;
 wire n_343;
 wire n_3432;
 wire n_3434;
 wire n_3436;
 wire n_3438;
 wire n_344;
 wire n_3440;
 wire n_3444;
 wire n_345;
 wire n_3452;
 wire n_3454;
 wire n_3456;
 wire n_3466;
 wire n_3468;
 wire n_347;
 wire n_3472;
 wire n_3474;
 wire n_3476;
 wire n_348;
 wire n_3480;
 wire n_3481;
 wire n_3483;
 wire n_3487;
 wire n_3488;
 wire n_3489;
 wire n_349;
 wire n_3490;
 wire n_3491;
 wire n_3494;
 wire n_3495;
 wire n_3496;
 wire n_3497;
 wire n_3498;
 wire n_3499;
 wire n_35;
 wire n_350;
 wire n_3500;
 wire n_3501;
 wire n_3502;
 wire n_3503;
 wire n_3504;
 wire n_3505;
 wire n_3506;
 wire n_3507;
 wire n_3508;
 wire n_3509;
 wire n_351;
 wire n_3510;
 wire n_3511;
 wire n_3512;
 wire n_3513;
 wire n_3514;
 wire n_3515;
 wire n_3516;
 wire n_3517;
 wire n_3518;
 wire n_3519;
 wire n_352;
 wire n_3520;
 wire n_3521;
 wire n_3522;
 wire n_3523;
 wire n_3524;
 wire n_3526;
 wire n_3527;
 wire n_3528;
 wire n_3529;
 wire n_353;
 wire n_3530;
 wire n_3531;
 wire n_3532;
 wire n_354;
 wire n_3541;
 wire n_3543;
 wire n_3544;
 wire n_3545;
 wire n_355;
 wire n_3555;
 wire n_3556;
 wire n_3557;
 wire n_3558;
 wire n_3559;
 wire n_356;
 wire n_3560;
 wire n_3561;
 wire n_3562;
 wire n_3563;
 wire n_3564;
 wire n_3565;
 wire n_3566;
 wire n_3567;
 wire n_3568;
 wire n_3569;
 wire n_357;
 wire n_3570;
 wire n_3571;
 wire n_3572;
 wire n_3573;
 wire n_3574;
 wire n_3575;
 wire n_3576;
 wire n_3577;
 wire n_3578;
 wire n_3579;
 wire n_358;
 wire n_3580;
 wire n_3581;
 wire n_3582;
 wire n_3583;
 wire n_3584;
 wire n_3585;
 wire n_3586;
 wire n_3587;
 wire n_3588;
 wire n_3589;
 wire n_3590;
 wire n_3591;
 wire n_3592;
 wire n_3593;
 wire n_3594;
 wire n_3595;
 wire n_3596;
 wire n_3597;
 wire n_3598;
 wire n_3599;
 wire n_36;
 wire n_360;
 wire n_361;
 wire n_362;
 wire n_3626;
 wire n_3627;
 wire n_3628;
 wire n_3629;
 wire n_363;
 wire n_3630;
 wire n_3631;
 wire n_3632;
 wire n_3633;
 wire n_3634;
 wire n_3635;
 wire n_3636;
 wire n_3637;
 wire n_3638;
 wire n_3639;
 wire n_364;
 wire n_3640;
 wire n_3641;
 wire n_3642;
 wire n_3643;
 wire n_3645;
 wire n_3646;
 wire n_3647;
 wire n_3648;
 wire n_3649;
 wire n_365;
 wire n_3650;
 wire n_3651;
 wire n_3652;
 wire n_3653;
 wire n_3654;
 wire n_3655;
 wire n_3656;
 wire n_3657;
 wire n_3658;
 wire n_3659;
 wire n_366;
 wire n_3660;
 wire n_3661;
 wire n_3662;
 wire n_3663;
 wire n_3664;
 wire n_3665;
 wire n_3666;
 wire n_367;
 wire n_368;
 wire n_369;
 wire n_37;
 wire n_370;
 wire n_371;
 wire n_3715;
 wire n_3716;
 wire n_3717;
 wire n_3718;
 wire n_3719;
 wire n_372;
 wire n_3720;
 wire n_3721;
 wire n_3722;
 wire n_3723;
 wire n_3724;
 wire n_3725;
 wire n_3726;
 wire n_3727;
 wire n_3728;
 wire n_3729;
 wire n_373;
 wire n_3730;
 wire n_3731;
 wire n_3732;
 wire n_3733;
 wire n_3734;
 wire n_3735;
 wire n_3736;
 wire n_3737;
 wire n_3738;
 wire n_3739;
 wire n_374;
 wire n_3740;
 wire n_3741;
 wire n_3742;
 wire n_3743;
 wire n_3744;
 wire n_3745;
 wire n_3746;
 wire n_3747;
 wire n_3748;
 wire n_3749;
 wire n_375;
 wire n_3750;
 wire n_3751;
 wire n_3752;
 wire n_3753;
 wire n_3754;
 wire n_3755;
 wire n_3756;
 wire n_3757;
 wire n_3758;
 wire n_3759;
 wire n_376;
 wire n_3760;
 wire n_3761;
 wire n_3762;
 wire n_3763;
 wire n_3764;
 wire n_3765;
 wire n_3766;
 wire n_3767;
 wire n_3768;
 wire n_3769;
 wire n_377;
 wire n_3770;
 wire n_3771;
 wire n_3772;
 wire n_3773;
 wire n_3774;
 wire n_3775;
 wire n_3776;
 wire n_3778;
 wire n_3779;
 wire n_378;
 wire n_3780;
 wire n_3781;
 wire n_3782;
 wire n_3783;
 wire n_3784;
 wire n_3785;
 wire n_3786;
 wire n_3787;
 wire n_3788;
 wire n_3789;
 wire n_379;
 wire n_3790;
 wire n_3791;
 wire n_3792;
 wire n_3793;
 wire n_3794;
 wire n_3795;
 wire n_3796;
 wire n_3797;
 wire n_3798;
 wire n_3799;
 wire n_38;
 wire n_380;
 wire n_3800;
 wire n_3801;
 wire n_3802;
 wire n_3803;
 wire n_3804;
 wire n_3805;
 wire n_3806;
 wire n_3807;
 wire n_3808;
 wire n_3809;
 wire n_381;
 wire n_3810;
 wire n_3811;
 wire n_3812;
 wire n_3813;
 wire n_3814;
 wire n_3815;
 wire n_3816;
 wire n_3817;
 wire n_3818;
 wire n_3819;
 wire n_382;
 wire n_3820;
 wire n_3821;
 wire n_3822;
 wire n_3823;
 wire n_3824;
 wire n_3825;
 wire n_3826;
 wire n_3827;
 wire n_3828;
 wire n_3829;
 wire n_383;
 wire n_3830;
 wire n_3831;
 wire n_3832;
 wire n_3833;
 wire n_3834;
 wire n_3835;
 wire n_3836;
 wire n_3837;
 wire n_3838;
 wire n_3839;
 wire n_384;
 wire n_3840;
 wire n_3844;
 wire n_3845;
 wire n_3846;
 wire n_3847;
 wire n_3848;
 wire n_3849;
 wire n_385;
 wire n_3850;
 wire n_386;
 wire n_387;
 wire n_388;
 wire n_389;
 wire n_39;
 wire n_390;
 wire n_391;
 wire n_392;
 wire n_393;
 wire n_394;
 wire n_395;
 wire n_396;
 wire n_397;
 wire n_398;
 wire n_399;
 wire n_4;
 wire n_40;
 wire n_400;
 wire n_401;
 wire n_402;
 wire n_403;
 wire n_404;
 wire n_405;
 wire n_406;
 wire n_407;
 wire n_408;
 wire n_409;
 wire n_41;
 wire n_410;
 wire n_411;
 wire n_412;
 wire n_413;
 wire n_414;
 wire n_415;
 wire n_416;
 wire n_417;
 wire n_418;
 wire n_419;
 wire n_42;
 wire n_420;
 wire n_421;
 wire n_422;
 wire n_423;
 wire n_424;
 wire n_425;
 wire n_426;
 wire n_427;
 wire n_428;
 wire n_429;
 wire n_43;
 wire n_430;
 wire n_431;
 wire n_432;
 wire n_433;
 wire n_434;
 wire n_435;
 wire n_436;
 wire n_437;
 wire n_438;
 wire n_439;
 wire n_44;
 wire n_440;
 wire n_441;
 wire n_442;
 wire n_443;
 wire n_444;
 wire n_445;
 wire n_446;
 wire n_447;
 wire n_448;
 wire n_449;
 wire n_45;
 wire n_450;
 wire n_451;
 wire n_452;
 wire n_453;
 wire n_454;
 wire n_455;
 wire n_456;
 wire n_457;
 wire n_458;
 wire n_459;
 wire n_46;
 wire n_460;
 wire n_461;
 wire n_462;
 wire n_463;
 wire n_464;
 wire n_465;
 wire n_466;
 wire n_467;
 wire n_468;
 wire n_469;
 wire n_47;
 wire n_470;
 wire n_471;
 wire n_472;
 wire n_473;
 wire n_474;
 wire n_475;
 wire n_476;
 wire n_477;
 wire n_478;
 wire n_479;
 wire n_48;
 wire n_480;
 wire n_481;
 wire n_483;
 wire n_484;
 wire n_485;
 wire n_486;
 wire n_487;
 wire n_489;
 wire n_49;
 wire n_490;
 wire n_491;
 wire n_492;
 wire n_493;
 wire n_494;
 wire n_495;
 wire n_496;
 wire n_497;
 wire n_498;
 wire n_499;
 wire n_5;
 wire n_50;
 wire n_500;
 wire n_501;
 wire n_502;
 wire n_503;
 wire n_504;
 wire n_505;
 wire n_506;
 wire n_507;
 wire n_508;
 wire n_509;
 wire n_51;
 wire n_510;
 wire n_511;
 wire n_512;
 wire n_513;
 wire n_514;
 wire n_515;
 wire n_516;
 wire n_517;
 wire n_518;
 wire n_519;
 wire n_520;
 wire n_521;
 wire n_522;
 wire n_523;
 wire n_524;
 wire n_525;
 wire n_526;
 wire n_527;
 wire n_528;
 wire n_529;
 wire n_53;
 wire n_530;
 wire n_531;
 wire n_532;
 wire n_533;
 wire n_534;
 wire n_535;
 wire n_536;
 wire n_537;
 wire n_538;
 wire n_539;
 wire n_54;
 wire n_540;
 wire n_541;
 wire n_542;
 wire n_543;
 wire n_544;
 wire n_545;
 wire n_546;
 wire n_547;
 wire n_548;
 wire n_549;
 wire n_55;
 wire n_550;
 wire n_551;
 wire n_552;
 wire n_553;
 wire n_554;
 wire n_555;
 wire n_556;
 wire n_557;
 wire n_558;
 wire n_559;
 wire n_56;
 wire n_560;
 wire n_561;
 wire n_562;
 wire n_563;
 wire n_564;
 wire n_565;
 wire n_566;
 wire n_567;
 wire n_568;
 wire n_569;
 wire n_57;
 wire n_570;
 wire n_571;
 wire n_572;
 wire n_573;
 wire n_574;
 wire n_575;
 wire n_576;
 wire n_577;
 wire n_578;
 wire n_579;
 wire n_58;
 wire n_580;
 wire n_581;
 wire n_582;
 wire n_583;
 wire n_584;
 wire n_585;
 wire n_586;
 wire n_587;
 wire n_588;
 wire n_589;
 wire n_59;
 wire n_590;
 wire n_591;
 wire n_592;
 wire n_593;
 wire n_594;
 wire n_595;
 wire n_596;
 wire n_597;
 wire n_598;
 wire n_599;
 wire n_600;
 wire n_601;
 wire n_602;
 wire n_603;
 wire n_604;
 wire n_605;
 wire n_606;
 wire n_607;
 wire n_608;
 wire n_609;
 wire n_61;
 wire n_610;
 wire n_611;
 wire n_612;
 wire n_613;
 wire n_614;
 wire n_615;
 wire n_616;
 wire n_617;
 wire n_618;
 wire n_619;
 wire n_62;
 wire n_620;
 wire n_621;
 wire n_622;
 wire n_623;
 wire n_624;
 wire n_625;
 wire n_626;
 wire n_627;
 wire n_628;
 wire n_629;
 wire n_63;
 wire n_630;
 wire n_631;
 wire n_632;
 wire n_633;
 wire n_634;
 wire n_635;
 wire n_636;
 wire n_637;
 wire n_638;
 wire n_639;
 wire n_64;
 wire n_640;
 wire n_642;
 wire n_643;
 wire n_644;
 wire n_645;
 wire n_646;
 wire n_647;
 wire n_648;
 wire n_649;
 wire n_65;
 wire n_650;
 wire n_651;
 wire n_652;
 wire n_653;
 wire n_654;
 wire n_655;
 wire n_656;
 wire n_657;
 wire n_658;
 wire n_659;
 wire n_66;
 wire n_660;
 wire n_661;
 wire n_662;
 wire n_663;
 wire n_664;
 wire n_665;
 wire n_666;
 wire n_667;
 wire n_668;
 wire n_669;
 wire n_67;
 wire n_670;
 wire n_671;
 wire n_672;
 wire n_674;
 wire n_675;
 wire n_676;
 wire n_677;
 wire n_678;
 wire n_679;
 wire n_68;
 wire n_680;
 wire n_681;
 wire n_682;
 wire n_683;
 wire n_686;
 wire n_687;
 wire n_688;
 wire n_689;
 wire n_69;
 wire n_690;
 wire n_691;
 wire n_692;
 wire n_693;
 wire n_694;
 wire n_695;
 wire n_696;
 wire n_697;
 wire n_699;
 wire n_7;
 wire n_70;
 wire n_700;
 wire n_702;
 wire n_706;
 wire n_71;
 wire n_712;
 wire n_713;
 wire n_714;
 wire n_715;
 wire n_716;
 wire n_717;
 wire n_718;
 wire n_719;
 wire n_72;
 wire n_720;
 wire n_721;
 wire n_722;
 wire n_723;
 wire n_724;
 wire n_725;
 wire n_726;
 wire n_727;
 wire n_728;
 wire n_73;
 wire n_733;
 wire n_737;
 wire n_74;
 wire n_740;
 wire n_742;
 wire n_743;
 wire n_746;
 wire n_75;
 wire n_751;
 wire n_76;
 wire n_761;
 wire n_763;
 wire n_769;
 wire n_77;
 wire n_771;
 wire n_774;
 wire n_78;
 wire n_79;
 wire n_790;
 wire n_792;
 wire n_795;
 wire n_796;
 wire n_797;
 wire n_798;
 wire n_799;
 wire n_8;
 wire n_80;
 wire n_800;
 wire n_801;
 wire n_802;
 wire n_805;
 wire n_809;
 wire n_81;
 wire n_810;
 wire n_817;
 wire n_82;
 wire n_822;
 wire n_83;
 wire n_830;
 wire n_833;
 wire n_834;
 wire n_838;
 wire n_839;
 wire n_84;
 wire n_844;
 wire n_847;
 wire n_848;
 wire n_849;
 wire n_85;
 wire n_851;
 wire n_852;
 wire n_853;
 wire n_854;
 wire n_856;
 wire n_86;
 wire n_866;
 wire n_87;
 wire n_870;
 wire n_872;
 wire n_875;
 wire n_876;
 wire n_877;
 wire n_878;
 wire n_879;
 wire n_88;
 wire n_880;
 wire n_881;
 wire n_882;
 wire n_883;
 wire n_884;
 wire n_885;
 wire n_886;
 wire n_887;
 wire n_888;
 wire n_889;
 wire n_89;
 wire n_890;
 wire n_891;
 wire n_892;
 wire n_893;
 wire n_894;
 wire n_895;
 wire n_896;
 wire n_897;
 wire n_898;
 wire n_9;
 wire n_90;
 wire n_900;
 wire n_901;
 wire n_902;
 wire n_903;
 wire n_904;
 wire n_905;
 wire n_906;
 wire n_907;
 wire n_908;
 wire n_909;
 wire n_91;
 wire n_910;
 wire n_911;
 wire n_912;
 wire n_913;
 wire n_914;
 wire n_915;
 wire n_916;
 wire n_917;
 wire n_918;
 wire n_919;
 wire n_92;
 wire n_920;
 wire n_921;
 wire n_922;
 wire n_923;
 wire n_925;
 wire n_927;
 wire n_928;
 wire n_929;
 wire n_93;
 wire n_930;
 wire n_931;
 wire n_932;
 wire n_933;
 wire n_934;
 wire n_935;
 wire n_936;
 wire n_937;
 wire n_938;
 wire n_94;
 wire n_940;
 wire n_941;
 wire n_942;
 wire n_943;
 wire n_944;
 wire n_945;
 wire n_946;
 wire n_947;
 wire n_948;
 wire n_949;
 wire n_95;
 wire n_950;
 wire n_951;
 wire n_952;
 wire n_953;
 wire n_954;
 wire n_955;
 wire n_956;
 wire n_957;
 wire n_958;
 wire n_959;
 wire n_96;
 wire n_960;
 wire n_961;
 wire n_962;
 wire n_963;
 wire n_964;
 wire n_965;
 wire n_966;
 wire n_967;
 wire n_968;
 wire n_969;
 wire n_97;
 wire n_970;
 wire n_971;
 wire n_972;
 wire n_973;
 wire n_974;
 wire n_975;
 wire n_976;
 wire n_977;
 wire n_978;
 wire n_979;
 wire n_98;
 wire n_980;
 wire n_981;
 wire n_982;
 wire n_983;
 wire n_984;
 wire n_985;
 wire n_986;
 wire n_987;
 wire n_988;
 wire n_989;
 wire n_99;
 wire n_991;
 wire n_992;
 wire n_994;
 wire n_995;
 wire n_996;
 wire n_997;
 wire n_998;
 wire n_999;
 wire nan_sign_d;
 wire opa_00;
 wire opa_dn;
 wire opa_inf;
 wire opa_nan;
 wire opa_nan_r;
 wire opas_r1;
 wire opas_r2;
 wire opb_00;
 wire opb_dn;
 wire opb_inf;
 wire opb_nan;
 wire qnan_d;
 wire result_zero_sign_d;
 wire sign;
 wire sign_exe;
 wire sign_exe_r;
 wire sign_fasu;
 wire sign_fasu_r;
 wire sign_mul;
 wire sign_mul_r;
 wire snan_d;
 wire sub_327_16_n_450;
 wire sub_327_16_n_454;
 wire sub_327_16_n_455;
 wire sub_327_16_n_459;
 wire sub_327_16_n_460;
 wire sub_327_16_n_464;
 wire sub_327_16_n_465;
 wire sub_327_16_n_469;
 wire sub_327_16_n_470;
 wire sub_327_16_n_474;
 wire sub_327_16_n_475;
 wire sub_327_16_n_479;
 wire sub_327_16_n_480;
 wire sub_327_16_n_484;
 wire sub_327_16_n_485;
 wire sub_327_16_n_489;
 wire sub_327_16_n_490;
 wire sub_327_16_n_494;
 wire sub_327_16_n_495;
 wire sub_327_16_n_499;
 wire sub_327_16_n_500;
 wire sub_327_16_n_504;
 wire sub_327_16_n_505;
 wire sub_327_16_n_509;
 wire sub_327_16_n_510;
 wire sub_327_16_n_514;
 wire sub_327_16_n_515;
 wire sub_327_16_n_519;
 wire sub_327_16_n_520;
 wire sub_327_16_n_524;
 wire sub_327_16_n_525;
 wire sub_327_16_n_529;
 wire sub_327_16_n_530;
 wire sub_327_16_n_534;
 wire sub_327_16_n_535;
 wire sub_327_16_n_539;
 wire sub_327_16_n_540;
 wire sub_327_16_n_544;
 wire sub_327_16_n_545;
 wire sub_327_16_n_549;
 wire sub_327_16_n_550;
 wire sub_327_16_n_554;
 wire sub_327_16_n_555;
 wire sub_327_16_n_559;
 wire sub_327_16_n_560;
 wire sub_327_16_n_564;
 wire sub_327_16_n_565;
 wire sub_327_16_n_569;
 wire sub_327_16_n_570;
 wire sub_327_16_n_574;
 wire sub_327_16_n_575;
 wire sub_327_16_n_579;
 wire sub_327_16_n_580;
 wire sub_327_16_n_584;
 wire sub_327_16_n_589;
 wire u0_expa_00;
 wire u0_expa_ff;
 wire u0_expb_00;
 wire u0_expb_ff;
 wire u0_fracta_00;
 wire u0_fractb_00;
 wire u0_infa_f_r;
 wire u0_infb_f_r;
 wire u0_n_321;
 wire u0_qnan_r_a;
 wire u0_qnan_r_b;
 wire u0_snan_r_a;
 wire u0_snan_r_b;
 wire u1_add_r;
 wire u1_fracta_eq_fractb;
 wire u1_fracta_lt_fractb;
 wire u1_n_1012;
 wire u1_n_1013;
 wire u1_n_1014;
 wire u1_n_1015;
 wire u1_n_1016;
 wire u1_n_1017;
 wire u1_n_1018;
 wire u1_n_1019;
 wire u1_n_1020;
 wire u1_n_1021;
 wire u1_n_1022;
 wire u1_n_1023;
 wire u1_n_1024;
 wire u1_n_1025;
 wire u1_n_1026;
 wire u1_n_1027;
 wire u1_n_1028;
 wire u1_n_1029;
 wire u1_n_1030;
 wire u1_n_1031;
 wire u1_n_1032;
 wire u1_n_1033;
 wire u1_n_1034;
 wire u1_n_1039;
 wire u1_n_1040;
 wire u1_n_1041;
 wire u1_n_1042;
 wire u1_n_1043;
 wire u1_n_1044;
 wire u1_n_1045;
 wire u1_n_1046;
 wire u1_n_1047;
 wire u1_n_1048;
 wire u1_n_1049;
 wire u1_n_1050;
 wire u1_n_1051;
 wire u1_n_1052;
 wire u1_n_1053;
 wire u1_n_1054;
 wire u1_n_1055;
 wire u1_n_1056;
 wire u1_n_1057;
 wire u1_n_1058;
 wire u1_n_1059;
 wire u1_n_1060;
 wire u1_n_1061;
 wire u1_n_1066;
 wire u1_n_1592;
 wire u1_n_1593;
 wire u1_n_1594;
 wire u1_n_2218;
 wire u1_n_3397;
 wire u1_n_4702;
 wire u1_n_4761;
 wire u1_n_4917;
 wire u1_n_4919;
 wire u1_n_4993;
 wire u1_n_5054;
 wire u1_n_5382;
 wire u1_n_5489;
 wire u1_n_590;
 wire u1_n_68;
 wire u1_n_8071;
 wire u1_n_840;
 wire u1_n_850;
 wire u1_n_852;
 wire u1_n_853;
 wire u1_n_867;
 wire u1_n_873;
 wire u1_n_880;
 wire u1_n_886;
 wire u1_n_909;
 wire u1_n_915;
 wire u1_n_917;
 wire u1_n_921;
 wire u1_n_923;
 wire u1_n_937;
 wire u1_n_941;
 wire u1_n_947;
 wire u1_n_966;
 wire u1_n_969;
 wire u1_n_972;
 wire u1_n_978;
 wire u1_n_980;
 wire u1_n_984;
 wire u1_n_986;
 wire u1_n_990;
 wire u1_n_992;
 wire u1_n_996;
 wire u1_n_997;
 wire u1_signa_r;
 wire u1_signb_r;
 wire u2_n_1384;
 wire u2_n_1392;
 wire u2_n_1398;
 wire u2_n_1399;
 wire u2_n_140;
 wire u2_n_1444;
 wire u2_n_1448;
 wire u2_n_1475;
 wire u2_n_1487;
 wire u2_n_1489;
 wire u2_n_1493;
 wire u2_n_1494;
 wire u2_n_1756;
 wire u2_n_1777;
 wire u2_n_1792;
 wire u2_n_1831;
 wire u2_n_606;
 wire u2_n_710;
 wire u2_n_772;
 wire u2_n_775;
 wire u3_sub_52_45_Y_add_52_31_n_630;
 wire u3_sub_52_45_Y_add_52_31_n_633;
 wire u3_sub_52_45_Y_add_52_31_n_636;
 wire u3_sub_52_45_Y_add_52_31_n_639;
 wire u3_sub_52_45_Y_add_52_31_n_642;
 wire u3_sub_52_45_Y_add_52_31_n_645;
 wire u3_sub_52_45_Y_add_52_31_n_648;
 wire u3_sub_52_45_Y_add_52_31_n_651;
 wire u3_sub_52_45_Y_add_52_31_n_654;
 wire u3_sub_52_45_Y_add_52_31_n_657;
 wire u3_sub_52_45_Y_add_52_31_n_660;
 wire u3_sub_52_45_Y_add_52_31_n_663;
 wire u3_sub_52_45_Y_add_52_31_n_666;
 wire u3_sub_52_45_Y_add_52_31_n_669;
 wire u3_sub_52_45_Y_add_52_31_n_672;
 wire u3_sub_52_45_Y_add_52_31_n_675;
 wire u3_sub_52_45_Y_add_52_31_n_678;
 wire u3_sub_52_45_Y_add_52_31_n_681;
 wire u3_sub_52_45_Y_add_52_31_n_684;
 wire u3_sub_52_45_Y_add_52_31_n_687;
 wire u3_sub_52_45_Y_add_52_31_n_690;
 wire u3_sub_52_45_Y_add_52_31_n_693;
 wire u3_sub_52_45_Y_add_52_31_n_696;
 wire u3_sub_52_45_Y_add_52_31_n_698;
 wire u3_sub_52_45_Y_add_52_31_n_699;
 wire u3_sub_52_45_Y_add_52_31_n_702;
 wire u3_sub_52_45_Y_add_52_31_n_762;
 wire u3_sub_52_45_Y_add_52_31_n_767;
 wire u3_sub_52_45_Y_add_52_31_n_770;
 wire u3_sub_52_45_Y_add_52_31_n_771;
 wire u3_sub_52_45_Y_add_52_31_n_772;
 wire u3_sub_52_45_Y_add_52_31_n_773;
 wire u3_sub_52_45_Y_add_52_31_n_774;
 wire u3_sub_52_45_Y_add_52_31_n_775;
 wire u3_sub_52_45_Y_add_52_31_n_776;
 wire u3_sub_52_45_Y_add_52_31_n_777;
 wire u3_sub_52_45_Y_add_52_31_n_778;
 wire u3_sub_52_45_Y_add_52_31_n_779;
 wire u3_sub_52_45_Y_add_52_31_n_780;
 wire u3_sub_52_45_Y_add_52_31_n_781;
 wire u3_sub_52_45_Y_add_52_31_n_782;
 wire u3_sub_52_45_Y_add_52_31_n_784;
 wire u3_sub_52_45_Y_add_52_31_n_785;
 wire u3_sub_52_45_Y_add_52_31_n_786;
 wire u3_sub_52_45_Y_add_52_31_n_787;
 wire u3_sub_52_45_Y_add_52_31_n_788;
 wire u3_sub_52_45_Y_add_52_31_n_789;
 wire u3_sub_52_45_Y_add_52_31_n_790;
 wire u3_sub_52_45_Y_add_52_31_n_791;
 wire u3_sub_52_45_Y_add_52_31_n_792;
 wire u3_sub_52_45_Y_add_52_31_n_793;
 wire u3_sub_52_45_Y_add_52_31_n_794;
 wire u3_sub_52_45_Y_add_52_31_n_795;
 wire u3_sub_52_45_Y_add_52_31_n_796;
 wire u3_sub_52_45_Y_add_52_31_n_797;
 wire u3_sub_52_45_Y_add_52_31_n_798;
 wire u3_sub_52_45_Y_add_52_31_n_803;
 wire u3_sub_52_45_Y_add_52_31_n_807;
 wire u3_sub_52_45_Y_add_52_31_n_809;
 wire u3_sub_52_45_Y_add_52_31_n_812;
 wire u3_sub_52_45_Y_add_52_31_n_817;
 wire u3_sub_52_45_Y_add_52_31_n_819;
 wire u3_sub_52_45_Y_add_52_31_n_821;
 wire u3_sub_52_45_Y_add_52_31_n_824;
 wire u3_sub_52_45_Y_add_52_31_n_829;
 wire u3_sub_52_45_Y_add_52_31_n_831;
 wire u3_sub_52_45_Y_add_52_31_n_841;
 wire u3_sub_52_45_Y_add_52_31_n_842;
 wire u4_exp_out1_co;
 wire u4_exp_zero;
 wire u4_f2i_zero;
 wire u4_g;
 wire u4_n_1091;
 wire u4_n_1248;
 wire u4_n_1266;
 wire u4_n_1362;
 wire u4_n_1438;
 wire u4_n_1439;
 wire u4_n_1442;
 wire u4_n_1446;
 wire u4_n_1454;
 wire u4_n_1722;
 wire u4_n_1792;
 wire u4_n_1793;
 wire u4_n_1794;
 wire u4_n_1795;
 wire u4_n_1796;
 wire u4_n_1797;
 wire u4_n_1798;
 wire u4_n_1799;
 wire u4_n_1800;
 wire u4_n_1801;
 wire u4_n_1802;
 wire u4_n_1803;
 wire u4_n_1804;
 wire u4_n_1805;
 wire u4_n_1806;
 wire u4_n_1807;
 wire u4_n_1808;
 wire u4_n_1809;
 wire u4_n_1810;
 wire u4_n_1811;
 wire u4_n_1812;
 wire u4_n_1813;
 wire u4_n_1814;
 wire u4_n_1815;
 wire u4_n_1816;
 wire u4_n_1817;
 wire u4_n_1818;
 wire u4_n_1819;
 wire u4_n_1820;
 wire u4_n_1821;
 wire u4_n_1822;
 wire u4_n_1823;
 wire u4_n_1824;
 wire u4_n_1825;
 wire u4_n_1826;
 wire u4_n_1827;
 wire u4_n_1828;
 wire u4_n_1829;
 wire u4_n_1830;
 wire u4_n_1831;
 wire u4_n_1832;
 wire u4_n_1833;
 wire u4_n_1834;
 wire u4_n_1835;
 wire u4_n_1836;
 wire u4_n_1837;
 wire u4_n_1838;
 wire u4_n_1839;
 wire u4_n_1840;
 wire u4_n_1841;
 wire u4_n_1842;
 wire u4_n_1843;
 wire u4_n_1844;
 wire u4_n_1845;
 wire u4_n_1846;
 wire u4_n_1847;
 wire u4_n_1848;
 wire u4_n_1849;
 wire u4_n_1850;
 wire u4_n_1851;
 wire u4_n_1852;
 wire u4_n_1934;
 wire u4_n_1938;
 wire u4_n_1942;
 wire u4_n_1944;
 wire u4_n_1946;
 wire u4_n_1948;
 wire u4_op_dn;
 wire u4_round2a_BAR;
 wire u4_sll_315_50_n_0;
 wire u4_sll_315_50_n_1;
 wire u4_sll_315_50_n_10;
 wire u4_sll_315_50_n_100;
 wire u4_sll_315_50_n_101;
 wire u4_sll_315_50_n_102;
 wire u4_sll_315_50_n_103;
 wire u4_sll_315_50_n_104;
 wire u4_sll_315_50_n_105;
 wire u4_sll_315_50_n_106;
 wire u4_sll_315_50_n_107;
 wire u4_sll_315_50_n_108;
 wire u4_sll_315_50_n_109;
 wire u4_sll_315_50_n_11;
 wire u4_sll_315_50_n_110;
 wire u4_sll_315_50_n_111;
 wire u4_sll_315_50_n_112;
 wire u4_sll_315_50_n_113;
 wire u4_sll_315_50_n_114;
 wire u4_sll_315_50_n_115;
 wire u4_sll_315_50_n_116;
 wire u4_sll_315_50_n_117;
 wire u4_sll_315_50_n_118;
 wire u4_sll_315_50_n_119;
 wire u4_sll_315_50_n_120;
 wire u4_sll_315_50_n_121;
 wire u4_sll_315_50_n_122;
 wire u4_sll_315_50_n_123;
 wire u4_sll_315_50_n_124;
 wire u4_sll_315_50_n_125;
 wire u4_sll_315_50_n_126;
 wire u4_sll_315_50_n_127;
 wire u4_sll_315_50_n_128;
 wire u4_sll_315_50_n_129;
 wire u4_sll_315_50_n_13;
 wire u4_sll_315_50_n_130;
 wire u4_sll_315_50_n_131;
 wire u4_sll_315_50_n_132;
 wire u4_sll_315_50_n_133;
 wire u4_sll_315_50_n_134;
 wire u4_sll_315_50_n_135;
 wire u4_sll_315_50_n_136;
 wire u4_sll_315_50_n_137;
 wire u4_sll_315_50_n_138;
 wire u4_sll_315_50_n_139;
 wire u4_sll_315_50_n_14;
 wire u4_sll_315_50_n_140;
 wire u4_sll_315_50_n_141;
 wire u4_sll_315_50_n_142;
 wire u4_sll_315_50_n_143;
 wire u4_sll_315_50_n_144;
 wire u4_sll_315_50_n_145;
 wire u4_sll_315_50_n_146;
 wire u4_sll_315_50_n_147;
 wire u4_sll_315_50_n_148;
 wire u4_sll_315_50_n_149;
 wire u4_sll_315_50_n_150;
 wire u4_sll_315_50_n_151;
 wire u4_sll_315_50_n_152;
 wire u4_sll_315_50_n_153;
 wire u4_sll_315_50_n_154;
 wire u4_sll_315_50_n_155;
 wire u4_sll_315_50_n_156;
 wire u4_sll_315_50_n_157;
 wire u4_sll_315_50_n_158;
 wire u4_sll_315_50_n_159;
 wire u4_sll_315_50_n_16;
 wire u4_sll_315_50_n_160;
 wire u4_sll_315_50_n_161;
 wire u4_sll_315_50_n_162;
 wire u4_sll_315_50_n_163;
 wire u4_sll_315_50_n_164;
 wire u4_sll_315_50_n_165;
 wire u4_sll_315_50_n_166;
 wire u4_sll_315_50_n_167;
 wire u4_sll_315_50_n_168;
 wire u4_sll_315_50_n_169;
 wire u4_sll_315_50_n_17;
 wire u4_sll_315_50_n_170;
 wire u4_sll_315_50_n_171;
 wire u4_sll_315_50_n_172;
 wire u4_sll_315_50_n_173;
 wire u4_sll_315_50_n_174;
 wire u4_sll_315_50_n_175;
 wire u4_sll_315_50_n_176;
 wire u4_sll_315_50_n_177;
 wire u4_sll_315_50_n_178;
 wire u4_sll_315_50_n_179;
 wire u4_sll_315_50_n_18;
 wire u4_sll_315_50_n_180;
 wire u4_sll_315_50_n_181;
 wire u4_sll_315_50_n_182;
 wire u4_sll_315_50_n_183;
 wire u4_sll_315_50_n_184;
 wire u4_sll_315_50_n_185;
 wire u4_sll_315_50_n_186;
 wire u4_sll_315_50_n_187;
 wire u4_sll_315_50_n_188;
 wire u4_sll_315_50_n_189;
 wire u4_sll_315_50_n_19;
 wire u4_sll_315_50_n_190;
 wire u4_sll_315_50_n_191;
 wire u4_sll_315_50_n_192;
 wire u4_sll_315_50_n_193;
 wire u4_sll_315_50_n_194;
 wire u4_sll_315_50_n_195;
 wire u4_sll_315_50_n_196;
 wire u4_sll_315_50_n_197;
 wire u4_sll_315_50_n_198;
 wire u4_sll_315_50_n_199;
 wire u4_sll_315_50_n_2;
 wire u4_sll_315_50_n_200;
 wire u4_sll_315_50_n_201;
 wire u4_sll_315_50_n_202;
 wire u4_sll_315_50_n_203;
 wire u4_sll_315_50_n_204;
 wire u4_sll_315_50_n_205;
 wire u4_sll_315_50_n_206;
 wire u4_sll_315_50_n_207;
 wire u4_sll_315_50_n_208;
 wire u4_sll_315_50_n_209;
 wire u4_sll_315_50_n_210;
 wire u4_sll_315_50_n_211;
 wire u4_sll_315_50_n_212;
 wire u4_sll_315_50_n_213;
 wire u4_sll_315_50_n_214;
 wire u4_sll_315_50_n_215;
 wire u4_sll_315_50_n_216;
 wire u4_sll_315_50_n_217;
 wire u4_sll_315_50_n_218;
 wire u4_sll_315_50_n_219;
 wire u4_sll_315_50_n_29;
 wire u4_sll_315_50_n_3;
 wire u4_sll_315_50_n_30;
 wire u4_sll_315_50_n_31;
 wire u4_sll_315_50_n_32;
 wire u4_sll_315_50_n_33;
 wire u4_sll_315_50_n_34;
 wire u4_sll_315_50_n_35;
 wire u4_sll_315_50_n_36;
 wire u4_sll_315_50_n_37;
 wire u4_sll_315_50_n_38;
 wire u4_sll_315_50_n_39;
 wire u4_sll_315_50_n_4;
 wire u4_sll_315_50_n_40;
 wire u4_sll_315_50_n_41;
 wire u4_sll_315_50_n_42;
 wire u4_sll_315_50_n_43;
 wire u4_sll_315_50_n_44;
 wire u4_sll_315_50_n_45;
 wire u4_sll_315_50_n_46;
 wire u4_sll_315_50_n_47;
 wire u4_sll_315_50_n_48;
 wire u4_sll_315_50_n_49;
 wire u4_sll_315_50_n_5;
 wire u4_sll_315_50_n_50;
 wire u4_sll_315_50_n_51;
 wire u4_sll_315_50_n_52;
 wire u4_sll_315_50_n_53;
 wire u4_sll_315_50_n_54;
 wire u4_sll_315_50_n_55;
 wire u4_sll_315_50_n_56;
 wire u4_sll_315_50_n_57;
 wire u4_sll_315_50_n_58;
 wire u4_sll_315_50_n_59;
 wire u4_sll_315_50_n_6;
 wire u4_sll_315_50_n_60;
 wire u4_sll_315_50_n_61;
 wire u4_sll_315_50_n_62;
 wire u4_sll_315_50_n_63;
 wire u4_sll_315_50_n_64;
 wire u4_sll_315_50_n_65;
 wire u4_sll_315_50_n_66;
 wire u4_sll_315_50_n_67;
 wire u4_sll_315_50_n_68;
 wire u4_sll_315_50_n_69;
 wire u4_sll_315_50_n_7;
 wire u4_sll_315_50_n_70;
 wire u4_sll_315_50_n_71;
 wire u4_sll_315_50_n_72;
 wire u4_sll_315_50_n_73;
 wire u4_sll_315_50_n_74;
 wire u4_sll_315_50_n_75;
 wire u4_sll_315_50_n_76;
 wire u4_sll_315_50_n_77;
 wire u4_sll_315_50_n_78;
 wire u4_sll_315_50_n_79;
 wire u4_sll_315_50_n_8;
 wire u4_sll_315_50_n_80;
 wire u4_sll_315_50_n_81;
 wire u4_sll_315_50_n_82;
 wire u4_sll_315_50_n_83;
 wire u4_sll_315_50_n_84;
 wire u4_sll_315_50_n_85;
 wire u4_sll_315_50_n_86;
 wire u4_sll_315_50_n_87;
 wire u4_sll_315_50_n_88;
 wire u4_sll_315_50_n_89;
 wire u4_sll_315_50_n_9;
 wire u4_sll_315_50_n_90;
 wire u4_sll_315_50_n_91;
 wire u4_sll_315_50_n_92;
 wire u4_sll_315_50_n_93;
 wire u4_sll_315_50_n_94;
 wire u4_sll_315_50_n_95;
 wire u4_sll_315_50_n_96;
 wire u4_sll_315_50_n_97;
 wire u4_sll_315_50_n_98;
 wire u4_sll_315_50_n_99;
 wire u5_mul_69_18_n_0;
 wire u5_mul_69_18_n_1;
 wire u5_mul_69_18_n_10;
 wire u5_mul_69_18_n_100;
 wire u5_mul_69_18_n_1000;
 wire u5_mul_69_18_n_1001;
 wire u5_mul_69_18_n_1002;
 wire u5_mul_69_18_n_1003;
 wire u5_mul_69_18_n_1008;
 wire u5_mul_69_18_n_1009;
 wire u5_mul_69_18_n_101;
 wire u5_mul_69_18_n_1012;
 wire u5_mul_69_18_n_1014;
 wire u5_mul_69_18_n_102;
 wire u5_mul_69_18_n_1020;
 wire u5_mul_69_18_n_1023;
 wire u5_mul_69_18_n_1024;
 wire u5_mul_69_18_n_1026;
 wire u5_mul_69_18_n_1027;
 wire u5_mul_69_18_n_1029;
 wire u5_mul_69_18_n_103;
 wire u5_mul_69_18_n_1032;
 wire u5_mul_69_18_n_1034;
 wire u5_mul_69_18_n_1035;
 wire u5_mul_69_18_n_1036;
 wire u5_mul_69_18_n_1037;
 wire u5_mul_69_18_n_104;
 wire u5_mul_69_18_n_1040;
 wire u5_mul_69_18_n_1041;
 wire u5_mul_69_18_n_1042;
 wire u5_mul_69_18_n_1044;
 wire u5_mul_69_18_n_1048;
 wire u5_mul_69_18_n_105;
 wire u5_mul_69_18_n_1050;
 wire u5_mul_69_18_n_1051;
 wire u5_mul_69_18_n_1057;
 wire u5_mul_69_18_n_1059;
 wire u5_mul_69_18_n_106;
 wire u5_mul_69_18_n_1060;
 wire u5_mul_69_18_n_1061;
 wire u5_mul_69_18_n_1062;
 wire u5_mul_69_18_n_1063;
 wire u5_mul_69_18_n_1065;
 wire u5_mul_69_18_n_1067;
 wire u5_mul_69_18_n_107;
 wire u5_mul_69_18_n_1071;
 wire u5_mul_69_18_n_1078;
 wire u5_mul_69_18_n_1079;
 wire u5_mul_69_18_n_108;
 wire u5_mul_69_18_n_1080;
 wire u5_mul_69_18_n_1084;
 wire u5_mul_69_18_n_1085;
 wire u5_mul_69_18_n_1088;
 wire u5_mul_69_18_n_1089;
 wire u5_mul_69_18_n_109;
 wire u5_mul_69_18_n_1093;
 wire u5_mul_69_18_n_1094;
 wire u5_mul_69_18_n_1095;
 wire u5_mul_69_18_n_1096;
 wire u5_mul_69_18_n_1097;
 wire u5_mul_69_18_n_11;
 wire u5_mul_69_18_n_110;
 wire u5_mul_69_18_n_1100;
 wire u5_mul_69_18_n_1103;
 wire u5_mul_69_18_n_1104;
 wire u5_mul_69_18_n_1106;
 wire u5_mul_69_18_n_1109;
 wire u5_mul_69_18_n_111;
 wire u5_mul_69_18_n_1114;
 wire u5_mul_69_18_n_1115;
 wire u5_mul_69_18_n_1116;
 wire u5_mul_69_18_n_1117;
 wire u5_mul_69_18_n_1118;
 wire u5_mul_69_18_n_1119;
 wire u5_mul_69_18_n_112;
 wire u5_mul_69_18_n_1120;
 wire u5_mul_69_18_n_1121;
 wire u5_mul_69_18_n_1122;
 wire u5_mul_69_18_n_1123;
 wire u5_mul_69_18_n_1124;
 wire u5_mul_69_18_n_1125;
 wire u5_mul_69_18_n_1126;
 wire u5_mul_69_18_n_1127;
 wire u5_mul_69_18_n_1128;
 wire u5_mul_69_18_n_1129;
 wire u5_mul_69_18_n_113;
 wire u5_mul_69_18_n_1130;
 wire u5_mul_69_18_n_1131;
 wire u5_mul_69_18_n_1132;
 wire u5_mul_69_18_n_1133;
 wire u5_mul_69_18_n_1134;
 wire u5_mul_69_18_n_1135;
 wire u5_mul_69_18_n_1136;
 wire u5_mul_69_18_n_1137;
 wire u5_mul_69_18_n_1138;
 wire u5_mul_69_18_n_1139;
 wire u5_mul_69_18_n_1140;
 wire u5_mul_69_18_n_1141;
 wire u5_mul_69_18_n_1142;
 wire u5_mul_69_18_n_1143;
 wire u5_mul_69_18_n_1144;
 wire u5_mul_69_18_n_1145;
 wire u5_mul_69_18_n_1146;
 wire u5_mul_69_18_n_1147;
 wire u5_mul_69_18_n_1148;
 wire u5_mul_69_18_n_1149;
 wire u5_mul_69_18_n_115;
 wire u5_mul_69_18_n_1150;
 wire u5_mul_69_18_n_1151;
 wire u5_mul_69_18_n_1152;
 wire u5_mul_69_18_n_1153;
 wire u5_mul_69_18_n_1154;
 wire u5_mul_69_18_n_1155;
 wire u5_mul_69_18_n_1156;
 wire u5_mul_69_18_n_1157;
 wire u5_mul_69_18_n_1158;
 wire u5_mul_69_18_n_1159;
 wire u5_mul_69_18_n_116;
 wire u5_mul_69_18_n_1160;
 wire u5_mul_69_18_n_1161;
 wire u5_mul_69_18_n_1162;
 wire u5_mul_69_18_n_1163;
 wire u5_mul_69_18_n_1164;
 wire u5_mul_69_18_n_1165;
 wire u5_mul_69_18_n_1166;
 wire u5_mul_69_18_n_1167;
 wire u5_mul_69_18_n_1168;
 wire u5_mul_69_18_n_1169;
 wire u5_mul_69_18_n_117;
 wire u5_mul_69_18_n_1170;
 wire u5_mul_69_18_n_1171;
 wire u5_mul_69_18_n_1172;
 wire u5_mul_69_18_n_1173;
 wire u5_mul_69_18_n_1174;
 wire u5_mul_69_18_n_1175;
 wire u5_mul_69_18_n_1176;
 wire u5_mul_69_18_n_118;
 wire u5_mul_69_18_n_1181;
 wire u5_mul_69_18_n_1186;
 wire u5_mul_69_18_n_1187;
 wire u5_mul_69_18_n_1188;
 wire u5_mul_69_18_n_1189;
 wire u5_mul_69_18_n_1190;
 wire u5_mul_69_18_n_1191;
 wire u5_mul_69_18_n_1192;
 wire u5_mul_69_18_n_1193;
 wire u5_mul_69_18_n_1194;
 wire u5_mul_69_18_n_1195;
 wire u5_mul_69_18_n_1196;
 wire u5_mul_69_18_n_1197;
 wire u5_mul_69_18_n_1198;
 wire u5_mul_69_18_n_1199;
 wire u5_mul_69_18_n_12;
 wire u5_mul_69_18_n_1200;
 wire u5_mul_69_18_n_1201;
 wire u5_mul_69_18_n_1202;
 wire u5_mul_69_18_n_1203;
 wire u5_mul_69_18_n_1204;
 wire u5_mul_69_18_n_1205;
 wire u5_mul_69_18_n_1206;
 wire u5_mul_69_18_n_1207;
 wire u5_mul_69_18_n_1208;
 wire u5_mul_69_18_n_1209;
 wire u5_mul_69_18_n_121;
 wire u5_mul_69_18_n_1210;
 wire u5_mul_69_18_n_1211;
 wire u5_mul_69_18_n_1212;
 wire u5_mul_69_18_n_1213;
 wire u5_mul_69_18_n_1214;
 wire u5_mul_69_18_n_1215;
 wire u5_mul_69_18_n_1216;
 wire u5_mul_69_18_n_1217;
 wire u5_mul_69_18_n_1218;
 wire u5_mul_69_18_n_1219;
 wire u5_mul_69_18_n_122;
 wire u5_mul_69_18_n_1220;
 wire u5_mul_69_18_n_1221;
 wire u5_mul_69_18_n_1222;
 wire u5_mul_69_18_n_1223;
 wire u5_mul_69_18_n_1224;
 wire u5_mul_69_18_n_1225;
 wire u5_mul_69_18_n_1226;
 wire u5_mul_69_18_n_1227;
 wire u5_mul_69_18_n_1228;
 wire u5_mul_69_18_n_1229;
 wire u5_mul_69_18_n_123;
 wire u5_mul_69_18_n_1232;
 wire u5_mul_69_18_n_1234;
 wire u5_mul_69_18_n_1236;
 wire u5_mul_69_18_n_1239;
 wire u5_mul_69_18_n_1241;
 wire u5_mul_69_18_n_1246;
 wire u5_mul_69_18_n_1247;
 wire u5_mul_69_18_n_1249;
 wire u5_mul_69_18_n_125;
 wire u5_mul_69_18_n_1256;
 wire u5_mul_69_18_n_1257;
 wire u5_mul_69_18_n_1258;
 wire u5_mul_69_18_n_1260;
 wire u5_mul_69_18_n_1265;
 wire u5_mul_69_18_n_1266;
 wire u5_mul_69_18_n_1267;
 wire u5_mul_69_18_n_1268;
 wire u5_mul_69_18_n_127;
 wire u5_mul_69_18_n_1270;
 wire u5_mul_69_18_n_1277;
 wire u5_mul_69_18_n_1278;
 wire u5_mul_69_18_n_1279;
 wire u5_mul_69_18_n_128;
 wire u5_mul_69_18_n_1284;
 wire u5_mul_69_18_n_1285;
 wire u5_mul_69_18_n_129;
 wire u5_mul_69_18_n_1291;
 wire u5_mul_69_18_n_1295;
 wire u5_mul_69_18_n_1298;
 wire u5_mul_69_18_n_13;
 wire u5_mul_69_18_n_130;
 wire u5_mul_69_18_n_1301;
 wire u5_mul_69_18_n_1303;
 wire u5_mul_69_18_n_1305;
 wire u5_mul_69_18_n_1306;
 wire u5_mul_69_18_n_1310;
 wire u5_mul_69_18_n_1311;
 wire u5_mul_69_18_n_1312;
 wire u5_mul_69_18_n_1313;
 wire u5_mul_69_18_n_1316;
 wire u5_mul_69_18_n_1319;
 wire u5_mul_69_18_n_132;
 wire u5_mul_69_18_n_1320;
 wire u5_mul_69_18_n_1322;
 wire u5_mul_69_18_n_1323;
 wire u5_mul_69_18_n_1324;
 wire u5_mul_69_18_n_1326;
 wire u5_mul_69_18_n_1327;
 wire u5_mul_69_18_n_1329;
 wire u5_mul_69_18_n_133;
 wire u5_mul_69_18_n_1330;
 wire u5_mul_69_18_n_1331;
 wire u5_mul_69_18_n_1332;
 wire u5_mul_69_18_n_1335;
 wire u5_mul_69_18_n_1339;
 wire u5_mul_69_18_n_134;
 wire u5_mul_69_18_n_1343;
 wire u5_mul_69_18_n_1344;
 wire u5_mul_69_18_n_1346;
 wire u5_mul_69_18_n_1352;
 wire u5_mul_69_18_n_1353;
 wire u5_mul_69_18_n_1354;
 wire u5_mul_69_18_n_1356;
 wire u5_mul_69_18_n_1357;
 wire u5_mul_69_18_n_1358;
 wire u5_mul_69_18_n_1359;
 wire u5_mul_69_18_n_1360;
 wire u5_mul_69_18_n_1361;
 wire u5_mul_69_18_n_1362;
 wire u5_mul_69_18_n_1363;
 wire u5_mul_69_18_n_1364;
 wire u5_mul_69_18_n_1365;
 wire u5_mul_69_18_n_1366;
 wire u5_mul_69_18_n_1367;
 wire u5_mul_69_18_n_1368;
 wire u5_mul_69_18_n_137;
 wire u5_mul_69_18_n_1371;
 wire u5_mul_69_18_n_1372;
 wire u5_mul_69_18_n_1375;
 wire u5_mul_69_18_n_1378;
 wire u5_mul_69_18_n_1379;
 wire u5_mul_69_18_n_138;
 wire u5_mul_69_18_n_1382;
 wire u5_mul_69_18_n_1383;
 wire u5_mul_69_18_n_1384;
 wire u5_mul_69_18_n_1386;
 wire u5_mul_69_18_n_1389;
 wire u5_mul_69_18_n_139;
 wire u5_mul_69_18_n_1391;
 wire u5_mul_69_18_n_1392;
 wire u5_mul_69_18_n_1393;
 wire u5_mul_69_18_n_1395;
 wire u5_mul_69_18_n_14;
 wire u5_mul_69_18_n_1402;
 wire u5_mul_69_18_n_1404;
 wire u5_mul_69_18_n_1405;
 wire u5_mul_69_18_n_1407;
 wire u5_mul_69_18_n_1409;
 wire u5_mul_69_18_n_141;
 wire u5_mul_69_18_n_1410;
 wire u5_mul_69_18_n_1411;
 wire u5_mul_69_18_n_1412;
 wire u5_mul_69_18_n_1413;
 wire u5_mul_69_18_n_1415;
 wire u5_mul_69_18_n_1416;
 wire u5_mul_69_18_n_1417;
 wire u5_mul_69_18_n_1418;
 wire u5_mul_69_18_n_1419;
 wire u5_mul_69_18_n_142;
 wire u5_mul_69_18_n_1420;
 wire u5_mul_69_18_n_1421;
 wire u5_mul_69_18_n_1422;
 wire u5_mul_69_18_n_1423;
 wire u5_mul_69_18_n_1424;
 wire u5_mul_69_18_n_1425;
 wire u5_mul_69_18_n_1426;
 wire u5_mul_69_18_n_1427;
 wire u5_mul_69_18_n_1429;
 wire u5_mul_69_18_n_143;
 wire u5_mul_69_18_n_1437;
 wire u5_mul_69_18_n_1439;
 wire u5_mul_69_18_n_144;
 wire u5_mul_69_18_n_1441;
 wire u5_mul_69_18_n_1444;
 wire u5_mul_69_18_n_1445;
 wire u5_mul_69_18_n_1446;
 wire u5_mul_69_18_n_1447;
 wire u5_mul_69_18_n_1448;
 wire u5_mul_69_18_n_1449;
 wire u5_mul_69_18_n_1452;
 wire u5_mul_69_18_n_1453;
 wire u5_mul_69_18_n_1455;
 wire u5_mul_69_18_n_1457;
 wire u5_mul_69_18_n_1458;
 wire u5_mul_69_18_n_146;
 wire u5_mul_69_18_n_1460;
 wire u5_mul_69_18_n_1461;
 wire u5_mul_69_18_n_1462;
 wire u5_mul_69_18_n_1463;
 wire u5_mul_69_18_n_1464;
 wire u5_mul_69_18_n_1465;
 wire u5_mul_69_18_n_1466;
 wire u5_mul_69_18_n_1467;
 wire u5_mul_69_18_n_1468;
 wire u5_mul_69_18_n_1469;
 wire u5_mul_69_18_n_1470;
 wire u5_mul_69_18_n_1471;
 wire u5_mul_69_18_n_1472;
 wire u5_mul_69_18_n_1473;
 wire u5_mul_69_18_n_1474;
 wire u5_mul_69_18_n_1475;
 wire u5_mul_69_18_n_1476;
 wire u5_mul_69_18_n_1477;
 wire u5_mul_69_18_n_1478;
 wire u5_mul_69_18_n_1479;
 wire u5_mul_69_18_n_148;
 wire u5_mul_69_18_n_1480;
 wire u5_mul_69_18_n_1481;
 wire u5_mul_69_18_n_1482;
 wire u5_mul_69_18_n_1483;
 wire u5_mul_69_18_n_1484;
 wire u5_mul_69_18_n_1485;
 wire u5_mul_69_18_n_1486;
 wire u5_mul_69_18_n_1487;
 wire u5_mul_69_18_n_1488;
 wire u5_mul_69_18_n_1489;
 wire u5_mul_69_18_n_149;
 wire u5_mul_69_18_n_1490;
 wire u5_mul_69_18_n_1491;
 wire u5_mul_69_18_n_1492;
 wire u5_mul_69_18_n_1493;
 wire u5_mul_69_18_n_1494;
 wire u5_mul_69_18_n_1495;
 wire u5_mul_69_18_n_1496;
 wire u5_mul_69_18_n_1497;
 wire u5_mul_69_18_n_1498;
 wire u5_mul_69_18_n_1499;
 wire u5_mul_69_18_n_150;
 wire u5_mul_69_18_n_1500;
 wire u5_mul_69_18_n_1501;
 wire u5_mul_69_18_n_1503;
 wire u5_mul_69_18_n_151;
 wire u5_mul_69_18_n_1510;
 wire u5_mul_69_18_n_1511;
 wire u5_mul_69_18_n_1514;
 wire u5_mul_69_18_n_1517;
 wire u5_mul_69_18_n_1518;
 wire u5_mul_69_18_n_152;
 wire u5_mul_69_18_n_1520;
 wire u5_mul_69_18_n_1523;
 wire u5_mul_69_18_n_1524;
 wire u5_mul_69_18_n_1527;
 wire u5_mul_69_18_n_1528;
 wire u5_mul_69_18_n_153;
 wire u5_mul_69_18_n_1531;
 wire u5_mul_69_18_n_1532;
 wire u5_mul_69_18_n_1534;
 wire u5_mul_69_18_n_1535;
 wire u5_mul_69_18_n_1537;
 wire u5_mul_69_18_n_1538;
 wire u5_mul_69_18_n_154;
 wire u5_mul_69_18_n_1540;
 wire u5_mul_69_18_n_1541;
 wire u5_mul_69_18_n_1546;
 wire u5_mul_69_18_n_1548;
 wire u5_mul_69_18_n_1549;
 wire u5_mul_69_18_n_155;
 wire u5_mul_69_18_n_1550;
 wire u5_mul_69_18_n_1551;
 wire u5_mul_69_18_n_1552;
 wire u5_mul_69_18_n_1554;
 wire u5_mul_69_18_n_1558;
 wire u5_mul_69_18_n_156;
 wire u5_mul_69_18_n_1560;
 wire u5_mul_69_18_n_1561;
 wire u5_mul_69_18_n_1563;
 wire u5_mul_69_18_n_1564;
 wire u5_mul_69_18_n_1565;
 wire u5_mul_69_18_n_1566;
 wire u5_mul_69_18_n_1567;
 wire u5_mul_69_18_n_1568;
 wire u5_mul_69_18_n_1569;
 wire u5_mul_69_18_n_157;
 wire u5_mul_69_18_n_1570;
 wire u5_mul_69_18_n_1572;
 wire u5_mul_69_18_n_1574;
 wire u5_mul_69_18_n_1575;
 wire u5_mul_69_18_n_1577;
 wire u5_mul_69_18_n_1578;
 wire u5_mul_69_18_n_1579;
 wire u5_mul_69_18_n_158;
 wire u5_mul_69_18_n_1581;
 wire u5_mul_69_18_n_1583;
 wire u5_mul_69_18_n_1587;
 wire u5_mul_69_18_n_159;
 wire u5_mul_69_18_n_1591;
 wire u5_mul_69_18_n_1594;
 wire u5_mul_69_18_n_1597;
 wire u5_mul_69_18_n_1598;
 wire u5_mul_69_18_n_1599;
 wire u5_mul_69_18_n_160;
 wire u5_mul_69_18_n_1600;
 wire u5_mul_69_18_n_1601;
 wire u5_mul_69_18_n_1602;
 wire u5_mul_69_18_n_1604;
 wire u5_mul_69_18_n_1606;
 wire u5_mul_69_18_n_161;
 wire u5_mul_69_18_n_1612;
 wire u5_mul_69_18_n_1614;
 wire u5_mul_69_18_n_1616;
 wire u5_mul_69_18_n_1617;
 wire u5_mul_69_18_n_1618;
 wire u5_mul_69_18_n_1619;
 wire u5_mul_69_18_n_162;
 wire u5_mul_69_18_n_1620;
 wire u5_mul_69_18_n_1621;
 wire u5_mul_69_18_n_1622;
 wire u5_mul_69_18_n_1624;
 wire u5_mul_69_18_n_1625;
 wire u5_mul_69_18_n_1626;
 wire u5_mul_69_18_n_1627;
 wire u5_mul_69_18_n_1628;
 wire u5_mul_69_18_n_163;
 wire u5_mul_69_18_n_1632;
 wire u5_mul_69_18_n_1633;
 wire u5_mul_69_18_n_1634;
 wire u5_mul_69_18_n_1638;
 wire u5_mul_69_18_n_1639;
 wire u5_mul_69_18_n_164;
 wire u5_mul_69_18_n_1641;
 wire u5_mul_69_18_n_1642;
 wire u5_mul_69_18_n_1643;
 wire u5_mul_69_18_n_1647;
 wire u5_mul_69_18_n_1649;
 wire u5_mul_69_18_n_165;
 wire u5_mul_69_18_n_1652;
 wire u5_mul_69_18_n_1653;
 wire u5_mul_69_18_n_1654;
 wire u5_mul_69_18_n_1655;
 wire u5_mul_69_18_n_1656;
 wire u5_mul_69_18_n_1657;
 wire u5_mul_69_18_n_1658;
 wire u5_mul_69_18_n_1659;
 wire u5_mul_69_18_n_166;
 wire u5_mul_69_18_n_1660;
 wire u5_mul_69_18_n_1661;
 wire u5_mul_69_18_n_1662;
 wire u5_mul_69_18_n_1663;
 wire u5_mul_69_18_n_1664;
 wire u5_mul_69_18_n_1665;
 wire u5_mul_69_18_n_1668;
 wire u5_mul_69_18_n_1669;
 wire u5_mul_69_18_n_167;
 wire u5_mul_69_18_n_1673;
 wire u5_mul_69_18_n_1677;
 wire u5_mul_69_18_n_1678;
 wire u5_mul_69_18_n_1679;
 wire u5_mul_69_18_n_168;
 wire u5_mul_69_18_n_1680;
 wire u5_mul_69_18_n_1682;
 wire u5_mul_69_18_n_1684;
 wire u5_mul_69_18_n_1686;
 wire u5_mul_69_18_n_1687;
 wire u5_mul_69_18_n_1688;
 wire u5_mul_69_18_n_1689;
 wire u5_mul_69_18_n_169;
 wire u5_mul_69_18_n_1691;
 wire u5_mul_69_18_n_1692;
 wire u5_mul_69_18_n_1693;
 wire u5_mul_69_18_n_1694;
 wire u5_mul_69_18_n_1695;
 wire u5_mul_69_18_n_1696;
 wire u5_mul_69_18_n_1697;
 wire u5_mul_69_18_n_1698;
 wire u5_mul_69_18_n_1699;
 wire u5_mul_69_18_n_170;
 wire u5_mul_69_18_n_1700;
 wire u5_mul_69_18_n_1701;
 wire u5_mul_69_18_n_1702;
 wire u5_mul_69_18_n_1703;
 wire u5_mul_69_18_n_1704;
 wire u5_mul_69_18_n_1705;
 wire u5_mul_69_18_n_1706;
 wire u5_mul_69_18_n_1707;
 wire u5_mul_69_18_n_1708;
 wire u5_mul_69_18_n_1709;
 wire u5_mul_69_18_n_171;
 wire u5_mul_69_18_n_1710;
 wire u5_mul_69_18_n_1711;
 wire u5_mul_69_18_n_1712;
 wire u5_mul_69_18_n_1713;
 wire u5_mul_69_18_n_1714;
 wire u5_mul_69_18_n_1716;
 wire u5_mul_69_18_n_1719;
 wire u5_mul_69_18_n_172;
 wire u5_mul_69_18_n_1721;
 wire u5_mul_69_18_n_1722;
 wire u5_mul_69_18_n_173;
 wire u5_mul_69_18_n_1731;
 wire u5_mul_69_18_n_1732;
 wire u5_mul_69_18_n_1733;
 wire u5_mul_69_18_n_1735;
 wire u5_mul_69_18_n_1737;
 wire u5_mul_69_18_n_1738;
 wire u5_mul_69_18_n_1739;
 wire u5_mul_69_18_n_174;
 wire u5_mul_69_18_n_1743;
 wire u5_mul_69_18_n_1745;
 wire u5_mul_69_18_n_1746;
 wire u5_mul_69_18_n_1748;
 wire u5_mul_69_18_n_1749;
 wire u5_mul_69_18_n_175;
 wire u5_mul_69_18_n_1750;
 wire u5_mul_69_18_n_1752;
 wire u5_mul_69_18_n_1753;
 wire u5_mul_69_18_n_1754;
 wire u5_mul_69_18_n_1756;
 wire u5_mul_69_18_n_1758;
 wire u5_mul_69_18_n_1759;
 wire u5_mul_69_18_n_176;
 wire u5_mul_69_18_n_1760;
 wire u5_mul_69_18_n_177;
 wire u5_mul_69_18_n_1770;
 wire u5_mul_69_18_n_1771;
 wire u5_mul_69_18_n_1772;
 wire u5_mul_69_18_n_1773;
 wire u5_mul_69_18_n_1774;
 wire u5_mul_69_18_n_1775;
 wire u5_mul_69_18_n_178;
 wire u5_mul_69_18_n_1780;
 wire u5_mul_69_18_n_1782;
 wire u5_mul_69_18_n_1783;
 wire u5_mul_69_18_n_1784;
 wire u5_mul_69_18_n_1785;
 wire u5_mul_69_18_n_1786;
 wire u5_mul_69_18_n_1787;
 wire u5_mul_69_18_n_1788;
 wire u5_mul_69_18_n_1789;
 wire u5_mul_69_18_n_179;
 wire u5_mul_69_18_n_1790;
 wire u5_mul_69_18_n_1794;
 wire u5_mul_69_18_n_1797;
 wire u5_mul_69_18_n_1798;
 wire u5_mul_69_18_n_1799;
 wire u5_mul_69_18_n_180;
 wire u5_mul_69_18_n_1800;
 wire u5_mul_69_18_n_1801;
 wire u5_mul_69_18_n_1802;
 wire u5_mul_69_18_n_1803;
 wire u5_mul_69_18_n_1804;
 wire u5_mul_69_18_n_1806;
 wire u5_mul_69_18_n_1807;
 wire u5_mul_69_18_n_1808;
 wire u5_mul_69_18_n_1809;
 wire u5_mul_69_18_n_181;
 wire u5_mul_69_18_n_1810;
 wire u5_mul_69_18_n_1811;
 wire u5_mul_69_18_n_1812;
 wire u5_mul_69_18_n_1817;
 wire u5_mul_69_18_n_1818;
 wire u5_mul_69_18_n_1819;
 wire u5_mul_69_18_n_182;
 wire u5_mul_69_18_n_1820;
 wire u5_mul_69_18_n_1821;
 wire u5_mul_69_18_n_1822;
 wire u5_mul_69_18_n_1823;
 wire u5_mul_69_18_n_1826;
 wire u5_mul_69_18_n_1828;
 wire u5_mul_69_18_n_1829;
 wire u5_mul_69_18_n_183;
 wire u5_mul_69_18_n_1830;
 wire u5_mul_69_18_n_1831;
 wire u5_mul_69_18_n_1832;
 wire u5_mul_69_18_n_1833;
 wire u5_mul_69_18_n_1835;
 wire u5_mul_69_18_n_1836;
 wire u5_mul_69_18_n_1837;
 wire u5_mul_69_18_n_1838;
 wire u5_mul_69_18_n_1839;
 wire u5_mul_69_18_n_184;
 wire u5_mul_69_18_n_1840;
 wire u5_mul_69_18_n_1841;
 wire u5_mul_69_18_n_1842;
 wire u5_mul_69_18_n_1843;
 wire u5_mul_69_18_n_1844;
 wire u5_mul_69_18_n_1846;
 wire u5_mul_69_18_n_1847;
 wire u5_mul_69_18_n_1848;
 wire u5_mul_69_18_n_1849;
 wire u5_mul_69_18_n_185;
 wire u5_mul_69_18_n_1850;
 wire u5_mul_69_18_n_1851;
 wire u5_mul_69_18_n_1852;
 wire u5_mul_69_18_n_1854;
 wire u5_mul_69_18_n_1856;
 wire u5_mul_69_18_n_1857;
 wire u5_mul_69_18_n_1858;
 wire u5_mul_69_18_n_1859;
 wire u5_mul_69_18_n_186;
 wire u5_mul_69_18_n_1860;
 wire u5_mul_69_18_n_1864;
 wire u5_mul_69_18_n_1866;
 wire u5_mul_69_18_n_1867;
 wire u5_mul_69_18_n_1868;
 wire u5_mul_69_18_n_1869;
 wire u5_mul_69_18_n_187;
 wire u5_mul_69_18_n_1872;
 wire u5_mul_69_18_n_1873;
 wire u5_mul_69_18_n_1874;
 wire u5_mul_69_18_n_1875;
 wire u5_mul_69_18_n_1876;
 wire u5_mul_69_18_n_188;
 wire u5_mul_69_18_n_1881;
 wire u5_mul_69_18_n_1882;
 wire u5_mul_69_18_n_1883;
 wire u5_mul_69_18_n_1884;
 wire u5_mul_69_18_n_1885;
 wire u5_mul_69_18_n_1887;
 wire u5_mul_69_18_n_1888;
 wire u5_mul_69_18_n_1889;
 wire u5_mul_69_18_n_189;
 wire u5_mul_69_18_n_1890;
 wire u5_mul_69_18_n_1891;
 wire u5_mul_69_18_n_1893;
 wire u5_mul_69_18_n_1894;
 wire u5_mul_69_18_n_1895;
 wire u5_mul_69_18_n_1896;
 wire u5_mul_69_18_n_1897;
 wire u5_mul_69_18_n_1898;
 wire u5_mul_69_18_n_1899;
 wire u5_mul_69_18_n_19;
 wire u5_mul_69_18_n_190;
 wire u5_mul_69_18_n_1900;
 wire u5_mul_69_18_n_1901;
 wire u5_mul_69_18_n_1902;
 wire u5_mul_69_18_n_1903;
 wire u5_mul_69_18_n_1905;
 wire u5_mul_69_18_n_1906;
 wire u5_mul_69_18_n_1907;
 wire u5_mul_69_18_n_1908;
 wire u5_mul_69_18_n_1909;
 wire u5_mul_69_18_n_191;
 wire u5_mul_69_18_n_1910;
 wire u5_mul_69_18_n_1911;
 wire u5_mul_69_18_n_1912;
 wire u5_mul_69_18_n_1913;
 wire u5_mul_69_18_n_1914;
 wire u5_mul_69_18_n_1915;
 wire u5_mul_69_18_n_1916;
 wire u5_mul_69_18_n_1917;
 wire u5_mul_69_18_n_1918;
 wire u5_mul_69_18_n_1919;
 wire u5_mul_69_18_n_192;
 wire u5_mul_69_18_n_1920;
 wire u5_mul_69_18_n_1921;
 wire u5_mul_69_18_n_1922;
 wire u5_mul_69_18_n_1923;
 wire u5_mul_69_18_n_1924;
 wire u5_mul_69_18_n_1925;
 wire u5_mul_69_18_n_1926;
 wire u5_mul_69_18_n_1929;
 wire u5_mul_69_18_n_193;
 wire u5_mul_69_18_n_1930;
 wire u5_mul_69_18_n_1931;
 wire u5_mul_69_18_n_1932;
 wire u5_mul_69_18_n_1933;
 wire u5_mul_69_18_n_1934;
 wire u5_mul_69_18_n_1935;
 wire u5_mul_69_18_n_1936;
 wire u5_mul_69_18_n_1937;
 wire u5_mul_69_18_n_1938;
 wire u5_mul_69_18_n_1939;
 wire u5_mul_69_18_n_194;
 wire u5_mul_69_18_n_1940;
 wire u5_mul_69_18_n_1941;
 wire u5_mul_69_18_n_1942;
 wire u5_mul_69_18_n_1943;
 wire u5_mul_69_18_n_1944;
 wire u5_mul_69_18_n_1945;
 wire u5_mul_69_18_n_1946;
 wire u5_mul_69_18_n_1947;
 wire u5_mul_69_18_n_1949;
 wire u5_mul_69_18_n_195;
 wire u5_mul_69_18_n_1950;
 wire u5_mul_69_18_n_1951;
 wire u5_mul_69_18_n_1952;
 wire u5_mul_69_18_n_1953;
 wire u5_mul_69_18_n_1954;
 wire u5_mul_69_18_n_1955;
 wire u5_mul_69_18_n_1956;
 wire u5_mul_69_18_n_1957;
 wire u5_mul_69_18_n_1958;
 wire u5_mul_69_18_n_1959;
 wire u5_mul_69_18_n_196;
 wire u5_mul_69_18_n_1960;
 wire u5_mul_69_18_n_1961;
 wire u5_mul_69_18_n_1962;
 wire u5_mul_69_18_n_1963;
 wire u5_mul_69_18_n_1965;
 wire u5_mul_69_18_n_1966;
 wire u5_mul_69_18_n_1968;
 wire u5_mul_69_18_n_197;
 wire u5_mul_69_18_n_1970;
 wire u5_mul_69_18_n_1972;
 wire u5_mul_69_18_n_1974;
 wire u5_mul_69_18_n_1976;
 wire u5_mul_69_18_n_1978;
 wire u5_mul_69_18_n_198;
 wire u5_mul_69_18_n_1980;
 wire u5_mul_69_18_n_1982;
 wire u5_mul_69_18_n_1984;
 wire u5_mul_69_18_n_1986;
 wire u5_mul_69_18_n_1988;
 wire u5_mul_69_18_n_199;
 wire u5_mul_69_18_n_1990;
 wire u5_mul_69_18_n_1992;
 wire u5_mul_69_18_n_1994;
 wire u5_mul_69_18_n_1996;
 wire u5_mul_69_18_n_1998;
 wire u5_mul_69_18_n_2;
 wire u5_mul_69_18_n_20;
 wire u5_mul_69_18_n_200;
 wire u5_mul_69_18_n_2000;
 wire u5_mul_69_18_n_2002;
 wire u5_mul_69_18_n_2004;
 wire u5_mul_69_18_n_2006;
 wire u5_mul_69_18_n_2008;
 wire u5_mul_69_18_n_201;
 wire u5_mul_69_18_n_2010;
 wire u5_mul_69_18_n_2012;
 wire u5_mul_69_18_n_2014;
 wire u5_mul_69_18_n_2016;
 wire u5_mul_69_18_n_2018;
 wire u5_mul_69_18_n_202;
 wire u5_mul_69_18_n_2020;
 wire u5_mul_69_18_n_2022;
 wire u5_mul_69_18_n_2024;
 wire u5_mul_69_18_n_2026;
 wire u5_mul_69_18_n_2028;
 wire u5_mul_69_18_n_203;
 wire u5_mul_69_18_n_2030;
 wire u5_mul_69_18_n_2032;
 wire u5_mul_69_18_n_2034;
 wire u5_mul_69_18_n_2036;
 wire u5_mul_69_18_n_204;
 wire u5_mul_69_18_n_205;
 wire u5_mul_69_18_n_206;
 wire u5_mul_69_18_n_207;
 wire u5_mul_69_18_n_208;
 wire u5_mul_69_18_n_209;
 wire u5_mul_69_18_n_210;
 wire u5_mul_69_18_n_211;
 wire u5_mul_69_18_n_212;
 wire u5_mul_69_18_n_213;
 wire u5_mul_69_18_n_214;
 wire u5_mul_69_18_n_215;
 wire u5_mul_69_18_n_216;
 wire u5_mul_69_18_n_217;
 wire u5_mul_69_18_n_218;
 wire u5_mul_69_18_n_219;
 wire u5_mul_69_18_n_22;
 wire u5_mul_69_18_n_220;
 wire u5_mul_69_18_n_221;
 wire u5_mul_69_18_n_222;
 wire u5_mul_69_18_n_223;
 wire u5_mul_69_18_n_225;
 wire u5_mul_69_18_n_226;
 wire u5_mul_69_18_n_227;
 wire u5_mul_69_18_n_228;
 wire u5_mul_69_18_n_229;
 wire u5_mul_69_18_n_23;
 wire u5_mul_69_18_n_230;
 wire u5_mul_69_18_n_231;
 wire u5_mul_69_18_n_232;
 wire u5_mul_69_18_n_233;
 wire u5_mul_69_18_n_234;
 wire u5_mul_69_18_n_235;
 wire u5_mul_69_18_n_236;
 wire u5_mul_69_18_n_237;
 wire u5_mul_69_18_n_238;
 wire u5_mul_69_18_n_239;
 wire u5_mul_69_18_n_24;
 wire u5_mul_69_18_n_240;
 wire u5_mul_69_18_n_241;
 wire u5_mul_69_18_n_242;
 wire u5_mul_69_18_n_243;
 wire u5_mul_69_18_n_244;
 wire u5_mul_69_18_n_245;
 wire u5_mul_69_18_n_246;
 wire u5_mul_69_18_n_247;
 wire u5_mul_69_18_n_248;
 wire u5_mul_69_18_n_249;
 wire u5_mul_69_18_n_25;
 wire u5_mul_69_18_n_250;
 wire u5_mul_69_18_n_251;
 wire u5_mul_69_18_n_252;
 wire u5_mul_69_18_n_253;
 wire u5_mul_69_18_n_254;
 wire u5_mul_69_18_n_255;
 wire u5_mul_69_18_n_256;
 wire u5_mul_69_18_n_257;
 wire u5_mul_69_18_n_258;
 wire u5_mul_69_18_n_259;
 wire u5_mul_69_18_n_26;
 wire u5_mul_69_18_n_260;
 wire u5_mul_69_18_n_261;
 wire u5_mul_69_18_n_262;
 wire u5_mul_69_18_n_263;
 wire u5_mul_69_18_n_264;
 wire u5_mul_69_18_n_265;
 wire u5_mul_69_18_n_266;
 wire u5_mul_69_18_n_267;
 wire u5_mul_69_18_n_268;
 wire u5_mul_69_18_n_269;
 wire u5_mul_69_18_n_27;
 wire u5_mul_69_18_n_270;
 wire u5_mul_69_18_n_271;
 wire u5_mul_69_18_n_272;
 wire u5_mul_69_18_n_273;
 wire u5_mul_69_18_n_274;
 wire u5_mul_69_18_n_275;
 wire u5_mul_69_18_n_276;
 wire u5_mul_69_18_n_277;
 wire u5_mul_69_18_n_278;
 wire u5_mul_69_18_n_279;
 wire u5_mul_69_18_n_28;
 wire u5_mul_69_18_n_280;
 wire u5_mul_69_18_n_281;
 wire u5_mul_69_18_n_282;
 wire u5_mul_69_18_n_283;
 wire u5_mul_69_18_n_284;
 wire u5_mul_69_18_n_285;
 wire u5_mul_69_18_n_286;
 wire u5_mul_69_18_n_287;
 wire u5_mul_69_18_n_288;
 wire u5_mul_69_18_n_289;
 wire u5_mul_69_18_n_29;
 wire u5_mul_69_18_n_290;
 wire u5_mul_69_18_n_291;
 wire u5_mul_69_18_n_292;
 wire u5_mul_69_18_n_293;
 wire u5_mul_69_18_n_294;
 wire u5_mul_69_18_n_295;
 wire u5_mul_69_18_n_296;
 wire u5_mul_69_18_n_297;
 wire u5_mul_69_18_n_298;
 wire u5_mul_69_18_n_299;
 wire u5_mul_69_18_n_3;
 wire u5_mul_69_18_n_30;
 wire u5_mul_69_18_n_300;
 wire u5_mul_69_18_n_301;
 wire u5_mul_69_18_n_302;
 wire u5_mul_69_18_n_303;
 wire u5_mul_69_18_n_304;
 wire u5_mul_69_18_n_305;
 wire u5_mul_69_18_n_306;
 wire u5_mul_69_18_n_307;
 wire u5_mul_69_18_n_308;
 wire u5_mul_69_18_n_309;
 wire u5_mul_69_18_n_31;
 wire u5_mul_69_18_n_310;
 wire u5_mul_69_18_n_311;
 wire u5_mul_69_18_n_312;
 wire u5_mul_69_18_n_313;
 wire u5_mul_69_18_n_314;
 wire u5_mul_69_18_n_315;
 wire u5_mul_69_18_n_316;
 wire u5_mul_69_18_n_317;
 wire u5_mul_69_18_n_318;
 wire u5_mul_69_18_n_319;
 wire u5_mul_69_18_n_32;
 wire u5_mul_69_18_n_320;
 wire u5_mul_69_18_n_321;
 wire u5_mul_69_18_n_322;
 wire u5_mul_69_18_n_323;
 wire u5_mul_69_18_n_324;
 wire u5_mul_69_18_n_325;
 wire u5_mul_69_18_n_326;
 wire u5_mul_69_18_n_327;
 wire u5_mul_69_18_n_328;
 wire u5_mul_69_18_n_329;
 wire u5_mul_69_18_n_33;
 wire u5_mul_69_18_n_330;
 wire u5_mul_69_18_n_331;
 wire u5_mul_69_18_n_332;
 wire u5_mul_69_18_n_333;
 wire u5_mul_69_18_n_334;
 wire u5_mul_69_18_n_335;
 wire u5_mul_69_18_n_336;
 wire u5_mul_69_18_n_337;
 wire u5_mul_69_18_n_338;
 wire u5_mul_69_18_n_339;
 wire u5_mul_69_18_n_34;
 wire u5_mul_69_18_n_340;
 wire u5_mul_69_18_n_341;
 wire u5_mul_69_18_n_342;
 wire u5_mul_69_18_n_343;
 wire u5_mul_69_18_n_344;
 wire u5_mul_69_18_n_345;
 wire u5_mul_69_18_n_346;
 wire u5_mul_69_18_n_347;
 wire u5_mul_69_18_n_348;
 wire u5_mul_69_18_n_349;
 wire u5_mul_69_18_n_35;
 wire u5_mul_69_18_n_350;
 wire u5_mul_69_18_n_351;
 wire u5_mul_69_18_n_352;
 wire u5_mul_69_18_n_353;
 wire u5_mul_69_18_n_354;
 wire u5_mul_69_18_n_355;
 wire u5_mul_69_18_n_356;
 wire u5_mul_69_18_n_357;
 wire u5_mul_69_18_n_358;
 wire u5_mul_69_18_n_359;
 wire u5_mul_69_18_n_36;
 wire u5_mul_69_18_n_360;
 wire u5_mul_69_18_n_361;
 wire u5_mul_69_18_n_362;
 wire u5_mul_69_18_n_363;
 wire u5_mul_69_18_n_364;
 wire u5_mul_69_18_n_365;
 wire u5_mul_69_18_n_366;
 wire u5_mul_69_18_n_367;
 wire u5_mul_69_18_n_368;
 wire u5_mul_69_18_n_369;
 wire u5_mul_69_18_n_37;
 wire u5_mul_69_18_n_370;
 wire u5_mul_69_18_n_371;
 wire u5_mul_69_18_n_372;
 wire u5_mul_69_18_n_373;
 wire u5_mul_69_18_n_374;
 wire u5_mul_69_18_n_375;
 wire u5_mul_69_18_n_376;
 wire u5_mul_69_18_n_377;
 wire u5_mul_69_18_n_378;
 wire u5_mul_69_18_n_379;
 wire u5_mul_69_18_n_38;
 wire u5_mul_69_18_n_380;
 wire u5_mul_69_18_n_381;
 wire u5_mul_69_18_n_382;
 wire u5_mul_69_18_n_383;
 wire u5_mul_69_18_n_384;
 wire u5_mul_69_18_n_385;
 wire u5_mul_69_18_n_386;
 wire u5_mul_69_18_n_387;
 wire u5_mul_69_18_n_388;
 wire u5_mul_69_18_n_389;
 wire u5_mul_69_18_n_39;
 wire u5_mul_69_18_n_390;
 wire u5_mul_69_18_n_391;
 wire u5_mul_69_18_n_392;
 wire u5_mul_69_18_n_393;
 wire u5_mul_69_18_n_394;
 wire u5_mul_69_18_n_395;
 wire u5_mul_69_18_n_396;
 wire u5_mul_69_18_n_397;
 wire u5_mul_69_18_n_398;
 wire u5_mul_69_18_n_399;
 wire u5_mul_69_18_n_40;
 wire u5_mul_69_18_n_400;
 wire u5_mul_69_18_n_401;
 wire u5_mul_69_18_n_402;
 wire u5_mul_69_18_n_403;
 wire u5_mul_69_18_n_404;
 wire u5_mul_69_18_n_405;
 wire u5_mul_69_18_n_406;
 wire u5_mul_69_18_n_407;
 wire u5_mul_69_18_n_408;
 wire u5_mul_69_18_n_409;
 wire u5_mul_69_18_n_41;
 wire u5_mul_69_18_n_410;
 wire u5_mul_69_18_n_411;
 wire u5_mul_69_18_n_412;
 wire u5_mul_69_18_n_413;
 wire u5_mul_69_18_n_414;
 wire u5_mul_69_18_n_415;
 wire u5_mul_69_18_n_416;
 wire u5_mul_69_18_n_417;
 wire u5_mul_69_18_n_418;
 wire u5_mul_69_18_n_419;
 wire u5_mul_69_18_n_42;
 wire u5_mul_69_18_n_420;
 wire u5_mul_69_18_n_421;
 wire u5_mul_69_18_n_422;
 wire u5_mul_69_18_n_423;
 wire u5_mul_69_18_n_424;
 wire u5_mul_69_18_n_425;
 wire u5_mul_69_18_n_426;
 wire u5_mul_69_18_n_427;
 wire u5_mul_69_18_n_428;
 wire u5_mul_69_18_n_429;
 wire u5_mul_69_18_n_43;
 wire u5_mul_69_18_n_430;
 wire u5_mul_69_18_n_431;
 wire u5_mul_69_18_n_432;
 wire u5_mul_69_18_n_433;
 wire u5_mul_69_18_n_434;
 wire u5_mul_69_18_n_435;
 wire u5_mul_69_18_n_436;
 wire u5_mul_69_18_n_437;
 wire u5_mul_69_18_n_438;
 wire u5_mul_69_18_n_439;
 wire u5_mul_69_18_n_44;
 wire u5_mul_69_18_n_440;
 wire u5_mul_69_18_n_441;
 wire u5_mul_69_18_n_442;
 wire u5_mul_69_18_n_443;
 wire u5_mul_69_18_n_444;
 wire u5_mul_69_18_n_445;
 wire u5_mul_69_18_n_446;
 wire u5_mul_69_18_n_447;
 wire u5_mul_69_18_n_448;
 wire u5_mul_69_18_n_449;
 wire u5_mul_69_18_n_45;
 wire u5_mul_69_18_n_450;
 wire u5_mul_69_18_n_451;
 wire u5_mul_69_18_n_452;
 wire u5_mul_69_18_n_453;
 wire u5_mul_69_18_n_454;
 wire u5_mul_69_18_n_455;
 wire u5_mul_69_18_n_456;
 wire u5_mul_69_18_n_457;
 wire u5_mul_69_18_n_458;
 wire u5_mul_69_18_n_459;
 wire u5_mul_69_18_n_46;
 wire u5_mul_69_18_n_460;
 wire u5_mul_69_18_n_461;
 wire u5_mul_69_18_n_462;
 wire u5_mul_69_18_n_463;
 wire u5_mul_69_18_n_464;
 wire u5_mul_69_18_n_465;
 wire u5_mul_69_18_n_466;
 wire u5_mul_69_18_n_467;
 wire u5_mul_69_18_n_468;
 wire u5_mul_69_18_n_469;
 wire u5_mul_69_18_n_47;
 wire u5_mul_69_18_n_470;
 wire u5_mul_69_18_n_471;
 wire u5_mul_69_18_n_472;
 wire u5_mul_69_18_n_473;
 wire u5_mul_69_18_n_474;
 wire u5_mul_69_18_n_475;
 wire u5_mul_69_18_n_476;
 wire u5_mul_69_18_n_477;
 wire u5_mul_69_18_n_478;
 wire u5_mul_69_18_n_479;
 wire u5_mul_69_18_n_48;
 wire u5_mul_69_18_n_480;
 wire u5_mul_69_18_n_481;
 wire u5_mul_69_18_n_482;
 wire u5_mul_69_18_n_483;
 wire u5_mul_69_18_n_484;
 wire u5_mul_69_18_n_485;
 wire u5_mul_69_18_n_486;
 wire u5_mul_69_18_n_487;
 wire u5_mul_69_18_n_488;
 wire u5_mul_69_18_n_489;
 wire u5_mul_69_18_n_49;
 wire u5_mul_69_18_n_490;
 wire u5_mul_69_18_n_491;
 wire u5_mul_69_18_n_492;
 wire u5_mul_69_18_n_493;
 wire u5_mul_69_18_n_494;
 wire u5_mul_69_18_n_495;
 wire u5_mul_69_18_n_496;
 wire u5_mul_69_18_n_497;
 wire u5_mul_69_18_n_498;
 wire u5_mul_69_18_n_499;
 wire u5_mul_69_18_n_5;
 wire u5_mul_69_18_n_50;
 wire u5_mul_69_18_n_500;
 wire u5_mul_69_18_n_501;
 wire u5_mul_69_18_n_502;
 wire u5_mul_69_18_n_503;
 wire u5_mul_69_18_n_504;
 wire u5_mul_69_18_n_505;
 wire u5_mul_69_18_n_506;
 wire u5_mul_69_18_n_507;
 wire u5_mul_69_18_n_508;
 wire u5_mul_69_18_n_509;
 wire u5_mul_69_18_n_51;
 wire u5_mul_69_18_n_510;
 wire u5_mul_69_18_n_511;
 wire u5_mul_69_18_n_512;
 wire u5_mul_69_18_n_513;
 wire u5_mul_69_18_n_514;
 wire u5_mul_69_18_n_515;
 wire u5_mul_69_18_n_516;
 wire u5_mul_69_18_n_517;
 wire u5_mul_69_18_n_518;
 wire u5_mul_69_18_n_519;
 wire u5_mul_69_18_n_52;
 wire u5_mul_69_18_n_520;
 wire u5_mul_69_18_n_521;
 wire u5_mul_69_18_n_522;
 wire u5_mul_69_18_n_523;
 wire u5_mul_69_18_n_524;
 wire u5_mul_69_18_n_525;
 wire u5_mul_69_18_n_526;
 wire u5_mul_69_18_n_527;
 wire u5_mul_69_18_n_528;
 wire u5_mul_69_18_n_529;
 wire u5_mul_69_18_n_53;
 wire u5_mul_69_18_n_530;
 wire u5_mul_69_18_n_531;
 wire u5_mul_69_18_n_532;
 wire u5_mul_69_18_n_533;
 wire u5_mul_69_18_n_534;
 wire u5_mul_69_18_n_535;
 wire u5_mul_69_18_n_536;
 wire u5_mul_69_18_n_537;
 wire u5_mul_69_18_n_538;
 wire u5_mul_69_18_n_539;
 wire u5_mul_69_18_n_54;
 wire u5_mul_69_18_n_540;
 wire u5_mul_69_18_n_541;
 wire u5_mul_69_18_n_542;
 wire u5_mul_69_18_n_543;
 wire u5_mul_69_18_n_544;
 wire u5_mul_69_18_n_545;
 wire u5_mul_69_18_n_546;
 wire u5_mul_69_18_n_547;
 wire u5_mul_69_18_n_548;
 wire u5_mul_69_18_n_549;
 wire u5_mul_69_18_n_55;
 wire u5_mul_69_18_n_550;
 wire u5_mul_69_18_n_551;
 wire u5_mul_69_18_n_552;
 wire u5_mul_69_18_n_553;
 wire u5_mul_69_18_n_554;
 wire u5_mul_69_18_n_555;
 wire u5_mul_69_18_n_556;
 wire u5_mul_69_18_n_557;
 wire u5_mul_69_18_n_558;
 wire u5_mul_69_18_n_559;
 wire u5_mul_69_18_n_56;
 wire u5_mul_69_18_n_560;
 wire u5_mul_69_18_n_561;
 wire u5_mul_69_18_n_562;
 wire u5_mul_69_18_n_563;
 wire u5_mul_69_18_n_564;
 wire u5_mul_69_18_n_565;
 wire u5_mul_69_18_n_566;
 wire u5_mul_69_18_n_567;
 wire u5_mul_69_18_n_568;
 wire u5_mul_69_18_n_569;
 wire u5_mul_69_18_n_57;
 wire u5_mul_69_18_n_570;
 wire u5_mul_69_18_n_571;
 wire u5_mul_69_18_n_572;
 wire u5_mul_69_18_n_573;
 wire u5_mul_69_18_n_574;
 wire u5_mul_69_18_n_575;
 wire u5_mul_69_18_n_576;
 wire u5_mul_69_18_n_577;
 wire u5_mul_69_18_n_578;
 wire u5_mul_69_18_n_579;
 wire u5_mul_69_18_n_58;
 wire u5_mul_69_18_n_580;
 wire u5_mul_69_18_n_581;
 wire u5_mul_69_18_n_582;
 wire u5_mul_69_18_n_583;
 wire u5_mul_69_18_n_584;
 wire u5_mul_69_18_n_585;
 wire u5_mul_69_18_n_586;
 wire u5_mul_69_18_n_587;
 wire u5_mul_69_18_n_588;
 wire u5_mul_69_18_n_589;
 wire u5_mul_69_18_n_59;
 wire u5_mul_69_18_n_590;
 wire u5_mul_69_18_n_591;
 wire u5_mul_69_18_n_592;
 wire u5_mul_69_18_n_593;
 wire u5_mul_69_18_n_594;
 wire u5_mul_69_18_n_595;
 wire u5_mul_69_18_n_596;
 wire u5_mul_69_18_n_597;
 wire u5_mul_69_18_n_598;
 wire u5_mul_69_18_n_599;
 wire u5_mul_69_18_n_6;
 wire u5_mul_69_18_n_60;
 wire u5_mul_69_18_n_600;
 wire u5_mul_69_18_n_601;
 wire u5_mul_69_18_n_602;
 wire u5_mul_69_18_n_603;
 wire u5_mul_69_18_n_604;
 wire u5_mul_69_18_n_605;
 wire u5_mul_69_18_n_606;
 wire u5_mul_69_18_n_607;
 wire u5_mul_69_18_n_608;
 wire u5_mul_69_18_n_609;
 wire u5_mul_69_18_n_61;
 wire u5_mul_69_18_n_610;
 wire u5_mul_69_18_n_611;
 wire u5_mul_69_18_n_612;
 wire u5_mul_69_18_n_613;
 wire u5_mul_69_18_n_614;
 wire u5_mul_69_18_n_615;
 wire u5_mul_69_18_n_616;
 wire u5_mul_69_18_n_617;
 wire u5_mul_69_18_n_618;
 wire u5_mul_69_18_n_619;
 wire u5_mul_69_18_n_62;
 wire u5_mul_69_18_n_620;
 wire u5_mul_69_18_n_621;
 wire u5_mul_69_18_n_622;
 wire u5_mul_69_18_n_623;
 wire u5_mul_69_18_n_624;
 wire u5_mul_69_18_n_625;
 wire u5_mul_69_18_n_626;
 wire u5_mul_69_18_n_627;
 wire u5_mul_69_18_n_628;
 wire u5_mul_69_18_n_629;
 wire u5_mul_69_18_n_63;
 wire u5_mul_69_18_n_630;
 wire u5_mul_69_18_n_631;
 wire u5_mul_69_18_n_632;
 wire u5_mul_69_18_n_633;
 wire u5_mul_69_18_n_634;
 wire u5_mul_69_18_n_635;
 wire u5_mul_69_18_n_636;
 wire u5_mul_69_18_n_637;
 wire u5_mul_69_18_n_638;
 wire u5_mul_69_18_n_639;
 wire u5_mul_69_18_n_64;
 wire u5_mul_69_18_n_640;
 wire u5_mul_69_18_n_641;
 wire u5_mul_69_18_n_642;
 wire u5_mul_69_18_n_643;
 wire u5_mul_69_18_n_644;
 wire u5_mul_69_18_n_645;
 wire u5_mul_69_18_n_646;
 wire u5_mul_69_18_n_647;
 wire u5_mul_69_18_n_648;
 wire u5_mul_69_18_n_649;
 wire u5_mul_69_18_n_65;
 wire u5_mul_69_18_n_650;
 wire u5_mul_69_18_n_651;
 wire u5_mul_69_18_n_652;
 wire u5_mul_69_18_n_653;
 wire u5_mul_69_18_n_654;
 wire u5_mul_69_18_n_655;
 wire u5_mul_69_18_n_656;
 wire u5_mul_69_18_n_657;
 wire u5_mul_69_18_n_658;
 wire u5_mul_69_18_n_659;
 wire u5_mul_69_18_n_66;
 wire u5_mul_69_18_n_660;
 wire u5_mul_69_18_n_661;
 wire u5_mul_69_18_n_662;
 wire u5_mul_69_18_n_663;
 wire u5_mul_69_18_n_664;
 wire u5_mul_69_18_n_665;
 wire u5_mul_69_18_n_666;
 wire u5_mul_69_18_n_667;
 wire u5_mul_69_18_n_668;
 wire u5_mul_69_18_n_669;
 wire u5_mul_69_18_n_67;
 wire u5_mul_69_18_n_670;
 wire u5_mul_69_18_n_671;
 wire u5_mul_69_18_n_672;
 wire u5_mul_69_18_n_673;
 wire u5_mul_69_18_n_674;
 wire u5_mul_69_18_n_675;
 wire u5_mul_69_18_n_676;
 wire u5_mul_69_18_n_677;
 wire u5_mul_69_18_n_678;
 wire u5_mul_69_18_n_679;
 wire u5_mul_69_18_n_68;
 wire u5_mul_69_18_n_680;
 wire u5_mul_69_18_n_681;
 wire u5_mul_69_18_n_682;
 wire u5_mul_69_18_n_683;
 wire u5_mul_69_18_n_684;
 wire u5_mul_69_18_n_685;
 wire u5_mul_69_18_n_686;
 wire u5_mul_69_18_n_687;
 wire u5_mul_69_18_n_688;
 wire u5_mul_69_18_n_689;
 wire u5_mul_69_18_n_69;
 wire u5_mul_69_18_n_690;
 wire u5_mul_69_18_n_691;
 wire u5_mul_69_18_n_692;
 wire u5_mul_69_18_n_693;
 wire u5_mul_69_18_n_694;
 wire u5_mul_69_18_n_695;
 wire u5_mul_69_18_n_696;
 wire u5_mul_69_18_n_697;
 wire u5_mul_69_18_n_698;
 wire u5_mul_69_18_n_699;
 wire u5_mul_69_18_n_7;
 wire u5_mul_69_18_n_70;
 wire u5_mul_69_18_n_700;
 wire u5_mul_69_18_n_701;
 wire u5_mul_69_18_n_702;
 wire u5_mul_69_18_n_703;
 wire u5_mul_69_18_n_704;
 wire u5_mul_69_18_n_705;
 wire u5_mul_69_18_n_706;
 wire u5_mul_69_18_n_707;
 wire u5_mul_69_18_n_708;
 wire u5_mul_69_18_n_709;
 wire u5_mul_69_18_n_71;
 wire u5_mul_69_18_n_710;
 wire u5_mul_69_18_n_711;
 wire u5_mul_69_18_n_712;
 wire u5_mul_69_18_n_713;
 wire u5_mul_69_18_n_714;
 wire u5_mul_69_18_n_715;
 wire u5_mul_69_18_n_716;
 wire u5_mul_69_18_n_717;
 wire u5_mul_69_18_n_718;
 wire u5_mul_69_18_n_719;
 wire u5_mul_69_18_n_72;
 wire u5_mul_69_18_n_720;
 wire u5_mul_69_18_n_721;
 wire u5_mul_69_18_n_722;
 wire u5_mul_69_18_n_723;
 wire u5_mul_69_18_n_724;
 wire u5_mul_69_18_n_725;
 wire u5_mul_69_18_n_726;
 wire u5_mul_69_18_n_727;
 wire u5_mul_69_18_n_728;
 wire u5_mul_69_18_n_729;
 wire u5_mul_69_18_n_73;
 wire u5_mul_69_18_n_730;
 wire u5_mul_69_18_n_731;
 wire u5_mul_69_18_n_732;
 wire u5_mul_69_18_n_733;
 wire u5_mul_69_18_n_734;
 wire u5_mul_69_18_n_735;
 wire u5_mul_69_18_n_736;
 wire u5_mul_69_18_n_737;
 wire u5_mul_69_18_n_738;
 wire u5_mul_69_18_n_739;
 wire u5_mul_69_18_n_74;
 wire u5_mul_69_18_n_740;
 wire u5_mul_69_18_n_741;
 wire u5_mul_69_18_n_742;
 wire u5_mul_69_18_n_743;
 wire u5_mul_69_18_n_744;
 wire u5_mul_69_18_n_745;
 wire u5_mul_69_18_n_746;
 wire u5_mul_69_18_n_747;
 wire u5_mul_69_18_n_748;
 wire u5_mul_69_18_n_749;
 wire u5_mul_69_18_n_750;
 wire u5_mul_69_18_n_751;
 wire u5_mul_69_18_n_752;
 wire u5_mul_69_18_n_753;
 wire u5_mul_69_18_n_754;
 wire u5_mul_69_18_n_755;
 wire u5_mul_69_18_n_756;
 wire u5_mul_69_18_n_757;
 wire u5_mul_69_18_n_758;
 wire u5_mul_69_18_n_759;
 wire u5_mul_69_18_n_760;
 wire u5_mul_69_18_n_761;
 wire u5_mul_69_18_n_762;
 wire u5_mul_69_18_n_763;
 wire u5_mul_69_18_n_764;
 wire u5_mul_69_18_n_765;
 wire u5_mul_69_18_n_766;
 wire u5_mul_69_18_n_767;
 wire u5_mul_69_18_n_768;
 wire u5_mul_69_18_n_769;
 wire u5_mul_69_18_n_77;
 wire u5_mul_69_18_n_770;
 wire u5_mul_69_18_n_771;
 wire u5_mul_69_18_n_772;
 wire u5_mul_69_18_n_773;
 wire u5_mul_69_18_n_774;
 wire u5_mul_69_18_n_775;
 wire u5_mul_69_18_n_776;
 wire u5_mul_69_18_n_777;
 wire u5_mul_69_18_n_778;
 wire u5_mul_69_18_n_779;
 wire u5_mul_69_18_n_78;
 wire u5_mul_69_18_n_780;
 wire u5_mul_69_18_n_781;
 wire u5_mul_69_18_n_782;
 wire u5_mul_69_18_n_783;
 wire u5_mul_69_18_n_784;
 wire u5_mul_69_18_n_785;
 wire u5_mul_69_18_n_786;
 wire u5_mul_69_18_n_787;
 wire u5_mul_69_18_n_788;
 wire u5_mul_69_18_n_789;
 wire u5_mul_69_18_n_79;
 wire u5_mul_69_18_n_790;
 wire u5_mul_69_18_n_791;
 wire u5_mul_69_18_n_792;
 wire u5_mul_69_18_n_793;
 wire u5_mul_69_18_n_794;
 wire u5_mul_69_18_n_795;
 wire u5_mul_69_18_n_796;
 wire u5_mul_69_18_n_797;
 wire u5_mul_69_18_n_798;
 wire u5_mul_69_18_n_799;
 wire u5_mul_69_18_n_8;
 wire u5_mul_69_18_n_800;
 wire u5_mul_69_18_n_801;
 wire u5_mul_69_18_n_802;
 wire u5_mul_69_18_n_803;
 wire u5_mul_69_18_n_804;
 wire u5_mul_69_18_n_805;
 wire u5_mul_69_18_n_806;
 wire u5_mul_69_18_n_807;
 wire u5_mul_69_18_n_808;
 wire u5_mul_69_18_n_809;
 wire u5_mul_69_18_n_810;
 wire u5_mul_69_18_n_811;
 wire u5_mul_69_18_n_812;
 wire u5_mul_69_18_n_813;
 wire u5_mul_69_18_n_814;
 wire u5_mul_69_18_n_815;
 wire u5_mul_69_18_n_816;
 wire u5_mul_69_18_n_817;
 wire u5_mul_69_18_n_818;
 wire u5_mul_69_18_n_819;
 wire u5_mul_69_18_n_82;
 wire u5_mul_69_18_n_820;
 wire u5_mul_69_18_n_821;
 wire u5_mul_69_18_n_822;
 wire u5_mul_69_18_n_823;
 wire u5_mul_69_18_n_824;
 wire u5_mul_69_18_n_825;
 wire u5_mul_69_18_n_826;
 wire u5_mul_69_18_n_827;
 wire u5_mul_69_18_n_828;
 wire u5_mul_69_18_n_829;
 wire u5_mul_69_18_n_83;
 wire u5_mul_69_18_n_830;
 wire u5_mul_69_18_n_831;
 wire u5_mul_69_18_n_832;
 wire u5_mul_69_18_n_833;
 wire u5_mul_69_18_n_834;
 wire u5_mul_69_18_n_835;
 wire u5_mul_69_18_n_836;
 wire u5_mul_69_18_n_837;
 wire u5_mul_69_18_n_838;
 wire u5_mul_69_18_n_839;
 wire u5_mul_69_18_n_84;
 wire u5_mul_69_18_n_840;
 wire u5_mul_69_18_n_841;
 wire u5_mul_69_18_n_842;
 wire u5_mul_69_18_n_843;
 wire u5_mul_69_18_n_844;
 wire u5_mul_69_18_n_845;
 wire u5_mul_69_18_n_846;
 wire u5_mul_69_18_n_847;
 wire u5_mul_69_18_n_848;
 wire u5_mul_69_18_n_849;
 wire u5_mul_69_18_n_85;
 wire u5_mul_69_18_n_850;
 wire u5_mul_69_18_n_851;
 wire u5_mul_69_18_n_852;
 wire u5_mul_69_18_n_853;
 wire u5_mul_69_18_n_854;
 wire u5_mul_69_18_n_855;
 wire u5_mul_69_18_n_856;
 wire u5_mul_69_18_n_857;
 wire u5_mul_69_18_n_858;
 wire u5_mul_69_18_n_859;
 wire u5_mul_69_18_n_860;
 wire u5_mul_69_18_n_861;
 wire u5_mul_69_18_n_862;
 wire u5_mul_69_18_n_863;
 wire u5_mul_69_18_n_864;
 wire u5_mul_69_18_n_865;
 wire u5_mul_69_18_n_866;
 wire u5_mul_69_18_n_867;
 wire u5_mul_69_18_n_868;
 wire u5_mul_69_18_n_869;
 wire u5_mul_69_18_n_87;
 wire u5_mul_69_18_n_870;
 wire u5_mul_69_18_n_871;
 wire u5_mul_69_18_n_872;
 wire u5_mul_69_18_n_873;
 wire u5_mul_69_18_n_874;
 wire u5_mul_69_18_n_875;
 wire u5_mul_69_18_n_876;
 wire u5_mul_69_18_n_877;
 wire u5_mul_69_18_n_878;
 wire u5_mul_69_18_n_879;
 wire u5_mul_69_18_n_88;
 wire u5_mul_69_18_n_880;
 wire u5_mul_69_18_n_881;
 wire u5_mul_69_18_n_882;
 wire u5_mul_69_18_n_883;
 wire u5_mul_69_18_n_884;
 wire u5_mul_69_18_n_885;
 wire u5_mul_69_18_n_886;
 wire u5_mul_69_18_n_887;
 wire u5_mul_69_18_n_888;
 wire u5_mul_69_18_n_889;
 wire u5_mul_69_18_n_89;
 wire u5_mul_69_18_n_890;
 wire u5_mul_69_18_n_891;
 wire u5_mul_69_18_n_892;
 wire u5_mul_69_18_n_893;
 wire u5_mul_69_18_n_894;
 wire u5_mul_69_18_n_895;
 wire u5_mul_69_18_n_896;
 wire u5_mul_69_18_n_897;
 wire u5_mul_69_18_n_898;
 wire u5_mul_69_18_n_899;
 wire u5_mul_69_18_n_9;
 wire u5_mul_69_18_n_900;
 wire u5_mul_69_18_n_901;
 wire u5_mul_69_18_n_902;
 wire u5_mul_69_18_n_903;
 wire u5_mul_69_18_n_904;
 wire u5_mul_69_18_n_905;
 wire u5_mul_69_18_n_906;
 wire u5_mul_69_18_n_907;
 wire u5_mul_69_18_n_908;
 wire u5_mul_69_18_n_909;
 wire u5_mul_69_18_n_91;
 wire u5_mul_69_18_n_910;
 wire u5_mul_69_18_n_911;
 wire u5_mul_69_18_n_912;
 wire u5_mul_69_18_n_913;
 wire u5_mul_69_18_n_914;
 wire u5_mul_69_18_n_915;
 wire u5_mul_69_18_n_916;
 wire u5_mul_69_18_n_917;
 wire u5_mul_69_18_n_918;
 wire u5_mul_69_18_n_919;
 wire u5_mul_69_18_n_92;
 wire u5_mul_69_18_n_920;
 wire u5_mul_69_18_n_921;
 wire u5_mul_69_18_n_922;
 wire u5_mul_69_18_n_923;
 wire u5_mul_69_18_n_924;
 wire u5_mul_69_18_n_925;
 wire u5_mul_69_18_n_926;
 wire u5_mul_69_18_n_927;
 wire u5_mul_69_18_n_928;
 wire u5_mul_69_18_n_929;
 wire u5_mul_69_18_n_93;
 wire u5_mul_69_18_n_930;
 wire u5_mul_69_18_n_931;
 wire u5_mul_69_18_n_932;
 wire u5_mul_69_18_n_933;
 wire u5_mul_69_18_n_934;
 wire u5_mul_69_18_n_935;
 wire u5_mul_69_18_n_936;
 wire u5_mul_69_18_n_937;
 wire u5_mul_69_18_n_938;
 wire u5_mul_69_18_n_939;
 wire u5_mul_69_18_n_94;
 wire u5_mul_69_18_n_940;
 wire u5_mul_69_18_n_941;
 wire u5_mul_69_18_n_942;
 wire u5_mul_69_18_n_943;
 wire u5_mul_69_18_n_944;
 wire u5_mul_69_18_n_945;
 wire u5_mul_69_18_n_946;
 wire u5_mul_69_18_n_947;
 wire u5_mul_69_18_n_948;
 wire u5_mul_69_18_n_949;
 wire u5_mul_69_18_n_95;
 wire u5_mul_69_18_n_950;
 wire u5_mul_69_18_n_951;
 wire u5_mul_69_18_n_952;
 wire u5_mul_69_18_n_953;
 wire u5_mul_69_18_n_954;
 wire u5_mul_69_18_n_955;
 wire u5_mul_69_18_n_956;
 wire u5_mul_69_18_n_957;
 wire u5_mul_69_18_n_958;
 wire u5_mul_69_18_n_959;
 wire u5_mul_69_18_n_96;
 wire u5_mul_69_18_n_960;
 wire u5_mul_69_18_n_961;
 wire u5_mul_69_18_n_962;
 wire u5_mul_69_18_n_963;
 wire u5_mul_69_18_n_964;
 wire u5_mul_69_18_n_965;
 wire u5_mul_69_18_n_966;
 wire u5_mul_69_18_n_967;
 wire u5_mul_69_18_n_968;
 wire u5_mul_69_18_n_969;
 wire u5_mul_69_18_n_97;
 wire u5_mul_69_18_n_970;
 wire u5_mul_69_18_n_971;
 wire u5_mul_69_18_n_972;
 wire u5_mul_69_18_n_973;
 wire u5_mul_69_18_n_974;
 wire u5_mul_69_18_n_975;
 wire u5_mul_69_18_n_976;
 wire u5_mul_69_18_n_977;
 wire u5_mul_69_18_n_978;
 wire u5_mul_69_18_n_979;
 wire u5_mul_69_18_n_98;
 wire u5_mul_69_18_n_980;
 wire u5_mul_69_18_n_981;
 wire u5_mul_69_18_n_982;
 wire u5_mul_69_18_n_983;
 wire u5_mul_69_18_n_984;
 wire u5_mul_69_18_n_985;
 wire u5_mul_69_18_n_986;
 wire u5_mul_69_18_n_99;
 wire u5_mul_69_18_n_991;
 wire u5_mul_69_18_n_992;
 wire u5_mul_69_18_n_993;
 wire u5_mul_69_18_n_994;
 wire u5_mul_69_18_n_995;
 wire u5_mul_69_18_n_996;
 wire u5_mul_69_18_n_998;
 wire u5_mul_69_18_n_999;
 wire u5_n_2;
 wire u6_n_101;
 wire u6_n_102;
 wire u6_n_104;
 wire u6_n_105;
 wire u6_n_108;
 wire u6_n_109;
 wire u6_n_111;
 wire u6_n_112;
 wire u6_n_113;
 wire u6_n_115;
 wire u6_n_116;
 wire u6_n_117;
 wire u6_n_118;
 wire u6_n_119;
 wire u6_n_120;
 wire u6_n_122;
 wire u6_n_123;
 wire u6_n_124;
 wire u6_n_126;
 wire u6_n_127;
 wire u6_n_128;
 wire u6_n_129;
 wire u6_n_130;
 wire u6_n_131;
 wire u6_n_132;
 wire u6_n_133;
 wire u6_n_134;
 wire u6_n_135;
 wire u6_n_136;
 wire u6_n_137;
 wire u6_n_138;
 wire u6_n_139;
 wire u6_n_140;
 wire u6_n_141;
 wire u6_n_142;
 wire u6_n_143;
 wire u6_n_144;
 wire u6_n_145;
 wire u6_n_146;
 wire u6_n_147;
 wire u6_n_148;
 wire u6_n_149;
 wire u6_n_76;
 wire u6_n_77;
 wire u6_n_79;
 wire u6_n_81;
 wire u6_n_82;
 wire u6_n_83;
 wire u6_n_84;
 wire u6_n_87;
 wire u6_n_89;
 wire u6_n_91;
 wire u6_n_93;
 wire u6_n_95;
 wire u6_n_96;
 wire u6_n_99;
 wire u6_rem_96_22_Y_u6_div_90_17_n_0;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10;
 wire u6_rem_96_22_Y_u6_div_90_17_n_100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_10999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11;
 wire u6_rem_96_22_Y_u6_div_90_17_n_110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_11999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12;
 wire u6_rem_96_22_Y_u6_div_90_17_n_120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_12999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13;
 wire u6_rem_96_22_Y_u6_div_90_17_n_130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_13743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_14;
 wire u6_rem_96_22_Y_u6_div_90_17_n_140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_15;
 wire u6_rem_96_22_Y_u6_div_90_17_n_150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_16;
 wire u6_rem_96_22_Y_u6_div_90_17_n_160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_17;
 wire u6_rem_96_22_Y_u6_div_90_17_n_170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_18;
 wire u6_rem_96_22_Y_u6_div_90_17_n_180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_19;
 wire u6_rem_96_22_Y_u6_div_90_17_n_190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_1999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2;
 wire u6_rem_96_22_Y_u6_div_90_17_n_20;
 wire u6_rem_96_22_Y_u6_div_90_17_n_200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_21;
 wire u6_rem_96_22_Y_u6_div_90_17_n_210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_22;
 wire u6_rem_96_22_Y_u6_div_90_17_n_220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_23;
 wire u6_rem_96_22_Y_u6_div_90_17_n_230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_24;
 wire u6_rem_96_22_Y_u6_div_90_17_n_240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_25;
 wire u6_rem_96_22_Y_u6_div_90_17_n_250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_26;
 wire u6_rem_96_22_Y_u6_div_90_17_n_260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_27;
 wire u6_rem_96_22_Y_u6_div_90_17_n_270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_28;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_29;
 wire u6_rem_96_22_Y_u6_div_90_17_n_290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_2999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3;
 wire u6_rem_96_22_Y_u6_div_90_17_n_30;
 wire u6_rem_96_22_Y_u6_div_90_17_n_300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_31;
 wire u6_rem_96_22_Y_u6_div_90_17_n_310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_32;
 wire u6_rem_96_22_Y_u6_div_90_17_n_320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_33;
 wire u6_rem_96_22_Y_u6_div_90_17_n_330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_34;
 wire u6_rem_96_22_Y_u6_div_90_17_n_340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_35;
 wire u6_rem_96_22_Y_u6_div_90_17_n_350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_36;
 wire u6_rem_96_22_Y_u6_div_90_17_n_360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_37;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_38;
 wire u6_rem_96_22_Y_u6_div_90_17_n_380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_3999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4;
 wire u6_rem_96_22_Y_u6_div_90_17_n_40;
 wire u6_rem_96_22_Y_u6_div_90_17_n_400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_41;
 wire u6_rem_96_22_Y_u6_div_90_17_n_410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_42;
 wire u6_rem_96_22_Y_u6_div_90_17_n_420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_43;
 wire u6_rem_96_22_Y_u6_div_90_17_n_430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_44;
 wire u6_rem_96_22_Y_u6_div_90_17_n_440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_45;
 wire u6_rem_96_22_Y_u6_div_90_17_n_450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_46;
 wire u6_rem_96_22_Y_u6_div_90_17_n_460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_47;
 wire u6_rem_96_22_Y_u6_div_90_17_n_470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_48;
 wire u6_rem_96_22_Y_u6_div_90_17_n_480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_49;
 wire u6_rem_96_22_Y_u6_div_90_17_n_490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_4999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5;
 wire u6_rem_96_22_Y_u6_div_90_17_n_50;
 wire u6_rem_96_22_Y_u6_div_90_17_n_500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_51;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_53;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_54;
 wire u6_rem_96_22_Y_u6_div_90_17_n_540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_55;
 wire u6_rem_96_22_Y_u6_div_90_17_n_550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_56;
 wire u6_rem_96_22_Y_u6_div_90_17_n_560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_57;
 wire u6_rem_96_22_Y_u6_div_90_17_n_570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_58;
 wire u6_rem_96_22_Y_u6_div_90_17_n_580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_59;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_5998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6;
 wire u6_rem_96_22_Y_u6_div_90_17_n_60;
 wire u6_rem_96_22_Y_u6_div_90_17_n_600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_61;
 wire u6_rem_96_22_Y_u6_div_90_17_n_610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_62;
 wire u6_rem_96_22_Y_u6_div_90_17_n_620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_63;
 wire u6_rem_96_22_Y_u6_div_90_17_n_630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_65;
 wire u6_rem_96_22_Y_u6_div_90_17_n_650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_67;
 wire u6_rem_96_22_Y_u6_div_90_17_n_670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_68;
 wire u6_rem_96_22_Y_u6_div_90_17_n_680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_69;
 wire u6_rem_96_22_Y_u6_div_90_17_n_690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_6999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7;
 wire u6_rem_96_22_Y_u6_div_90_17_n_70;
 wire u6_rem_96_22_Y_u6_div_90_17_n_700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_72;
 wire u6_rem_96_22_Y_u6_div_90_17_n_720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_73;
 wire u6_rem_96_22_Y_u6_div_90_17_n_730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_74;
 wire u6_rem_96_22_Y_u6_div_90_17_n_740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_75;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_76;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_77;
 wire u6_rem_96_22_Y_u6_div_90_17_n_770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_78;
 wire u6_rem_96_22_Y_u6_div_90_17_n_780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_79;
 wire u6_rem_96_22_Y_u6_div_90_17_n_790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_7999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8;
 wire u6_rem_96_22_Y_u6_div_90_17_n_80;
 wire u6_rem_96_22_Y_u6_div_90_17_n_800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8052;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8085;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8088;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8121;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_82;
 wire u6_rem_96_22_Y_u6_div_90_17_n_820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8232;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_84;
 wire u6_rem_96_22_Y_u6_div_90_17_n_840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_85;
 wire u6_rem_96_22_Y_u6_div_90_17_n_850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8508;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_86;
 wire u6_rem_96_22_Y_u6_div_90_17_n_860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8646;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8682;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_87;
 wire u6_rem_96_22_Y_u6_div_90_17_n_870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8738;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8767;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_88;
 wire u6_rem_96_22_Y_u6_div_90_17_n_880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8800;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_8999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9;
 wire u6_rem_96_22_Y_u6_div_90_17_n_90;
 wire u6_rem_96_22_Y_u6_div_90_17_n_900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9000;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9001;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9002;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9003;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9004;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9005;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9006;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9007;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9008;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9009;
 wire u6_rem_96_22_Y_u6_div_90_17_n_901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9010;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9011;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9012;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9013;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9014;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9015;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9016;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9017;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9018;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9019;
 wire u6_rem_96_22_Y_u6_div_90_17_n_902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9020;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9021;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9022;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9023;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9024;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9025;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9026;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9027;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9028;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9029;
 wire u6_rem_96_22_Y_u6_div_90_17_n_903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9030;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9031;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9032;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9033;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9034;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9035;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9036;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9037;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9038;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9039;
 wire u6_rem_96_22_Y_u6_div_90_17_n_904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9040;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9041;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9042;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9043;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9044;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9045;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9046;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9047;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9048;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9049;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9050;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9051;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9053;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9054;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9055;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9056;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9057;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9058;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9059;
 wire u6_rem_96_22_Y_u6_div_90_17_n_906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9060;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9061;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9062;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9063;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9064;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9065;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9066;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9067;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9068;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9069;
 wire u6_rem_96_22_Y_u6_div_90_17_n_907;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9070;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9071;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9072;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9073;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9074;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9075;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9076;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9077;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9078;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9079;
 wire u6_rem_96_22_Y_u6_div_90_17_n_908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9080;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9081;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9082;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9083;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9084;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9086;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9087;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9089;
 wire u6_rem_96_22_Y_u6_div_90_17_n_909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9090;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9091;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9092;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9093;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9094;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9095;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9096;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9097;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9098;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9099;
 wire u6_rem_96_22_Y_u6_div_90_17_n_91;
 wire u6_rem_96_22_Y_u6_div_90_17_n_910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9100;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9101;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9102;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9103;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9104;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9105;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9106;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9107;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9108;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9109;
 wire u6_rem_96_22_Y_u6_div_90_17_n_911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9110;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9111;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9112;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9113;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9114;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9115;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9116;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9117;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9118;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9119;
 wire u6_rem_96_22_Y_u6_div_90_17_n_912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9120;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9122;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9123;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9124;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9125;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9126;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9127;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9128;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9129;
 wire u6_rem_96_22_Y_u6_div_90_17_n_913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9130;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9131;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9132;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9133;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9134;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9135;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9136;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9137;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9138;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9139;
 wire u6_rem_96_22_Y_u6_div_90_17_n_914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9140;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9141;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9142;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9143;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9144;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9145;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9146;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9147;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9148;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9149;
 wire u6_rem_96_22_Y_u6_div_90_17_n_915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9150;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9151;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9152;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9153;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9154;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9155;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9156;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9157;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9158;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9159;
 wire u6_rem_96_22_Y_u6_div_90_17_n_916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9160;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9161;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9162;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9163;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9164;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9165;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9166;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9167;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9168;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9169;
 wire u6_rem_96_22_Y_u6_div_90_17_n_917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9170;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9171;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9172;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9173;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9174;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9175;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9176;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9177;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9178;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9179;
 wire u6_rem_96_22_Y_u6_div_90_17_n_918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9180;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9181;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9182;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9183;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9184;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9185;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9186;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9187;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9188;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9189;
 wire u6_rem_96_22_Y_u6_div_90_17_n_919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9190;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9191;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9192;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9193;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9194;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9195;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9196;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9197;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9198;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9199;
 wire u6_rem_96_22_Y_u6_div_90_17_n_92;
 wire u6_rem_96_22_Y_u6_div_90_17_n_920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9200;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9201;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9202;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9203;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9204;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9205;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9206;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9207;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9208;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9209;
 wire u6_rem_96_22_Y_u6_div_90_17_n_921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9210;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9211;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9212;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9213;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9214;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9215;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9216;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9217;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9218;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9219;
 wire u6_rem_96_22_Y_u6_div_90_17_n_922;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9220;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9221;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9222;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9223;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9224;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9225;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9226;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9227;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9228;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9229;
 wire u6_rem_96_22_Y_u6_div_90_17_n_923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9230;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9231;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9233;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9234;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9235;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9236;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9237;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9238;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9239;
 wire u6_rem_96_22_Y_u6_div_90_17_n_924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9240;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9241;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9242;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9243;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9244;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9245;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9246;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9247;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9248;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9249;
 wire u6_rem_96_22_Y_u6_div_90_17_n_925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9250;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9251;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9252;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9253;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9254;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9255;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9256;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9257;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9258;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9259;
 wire u6_rem_96_22_Y_u6_div_90_17_n_926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9260;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9261;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9262;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9263;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9264;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9265;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9266;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9267;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9268;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9269;
 wire u6_rem_96_22_Y_u6_div_90_17_n_927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9270;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9271;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9272;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9273;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9274;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9275;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9276;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9277;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9278;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9279;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9280;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9281;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9282;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9283;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9284;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9285;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9286;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9287;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9288;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9289;
 wire u6_rem_96_22_Y_u6_div_90_17_n_929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9290;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9291;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9292;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9293;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9294;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9295;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9296;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9297;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9298;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9299;
 wire u6_rem_96_22_Y_u6_div_90_17_n_93;
 wire u6_rem_96_22_Y_u6_div_90_17_n_930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9300;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9301;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9302;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9303;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9304;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9305;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9306;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9307;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9308;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9309;
 wire u6_rem_96_22_Y_u6_div_90_17_n_931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9310;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9311;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9312;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9313;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9314;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9315;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9316;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9317;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9318;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9319;
 wire u6_rem_96_22_Y_u6_div_90_17_n_932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9320;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9321;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9322;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9323;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9324;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9325;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9326;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9327;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9328;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9329;
 wire u6_rem_96_22_Y_u6_div_90_17_n_933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9330;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9331;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9332;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9333;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9334;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9335;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9336;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9337;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9338;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9339;
 wire u6_rem_96_22_Y_u6_div_90_17_n_934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9340;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9341;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9342;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9343;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9344;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9345;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9346;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9347;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9348;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9349;
 wire u6_rem_96_22_Y_u6_div_90_17_n_935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9350;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9351;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9352;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9353;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9354;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9355;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9356;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9357;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9358;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9359;
 wire u6_rem_96_22_Y_u6_div_90_17_n_936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9360;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9361;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9362;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9363;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9364;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9365;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9366;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9367;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9368;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9369;
 wire u6_rem_96_22_Y_u6_div_90_17_n_937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9370;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9371;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9372;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9373;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9374;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9375;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9376;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9377;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9378;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9379;
 wire u6_rem_96_22_Y_u6_div_90_17_n_938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9380;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9381;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9382;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9383;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9384;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9385;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9386;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9387;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9388;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9389;
 wire u6_rem_96_22_Y_u6_div_90_17_n_939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9390;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9391;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9392;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9393;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9394;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9395;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9396;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9397;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9398;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9399;
 wire u6_rem_96_22_Y_u6_div_90_17_n_94;
 wire u6_rem_96_22_Y_u6_div_90_17_n_940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9400;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9401;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9402;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9403;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9404;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9405;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9406;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9407;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9408;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9409;
 wire u6_rem_96_22_Y_u6_div_90_17_n_941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9410;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9411;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9412;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9413;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9414;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9415;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9416;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9417;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9418;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9419;
 wire u6_rem_96_22_Y_u6_div_90_17_n_942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9420;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9421;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9422;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9423;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9424;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9425;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9426;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9427;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9428;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9429;
 wire u6_rem_96_22_Y_u6_div_90_17_n_943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9430;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9431;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9432;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9433;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9434;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9435;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9436;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9437;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9438;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9439;
 wire u6_rem_96_22_Y_u6_div_90_17_n_944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9440;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9441;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9442;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9443;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9444;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9445;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9446;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9447;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9448;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9449;
 wire u6_rem_96_22_Y_u6_div_90_17_n_945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9450;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9451;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9452;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9453;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9454;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9455;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9456;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9457;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9458;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9459;
 wire u6_rem_96_22_Y_u6_div_90_17_n_946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9460;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9461;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9462;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9463;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9464;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9465;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9466;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9467;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9468;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9469;
 wire u6_rem_96_22_Y_u6_div_90_17_n_947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9470;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9471;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9472;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9473;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9474;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9475;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9476;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9477;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9478;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9479;
 wire u6_rem_96_22_Y_u6_div_90_17_n_948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9480;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9481;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9482;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9483;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9484;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9485;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9486;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9487;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9488;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9489;
 wire u6_rem_96_22_Y_u6_div_90_17_n_949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9490;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9491;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9492;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9493;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9494;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9495;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9496;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9497;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9498;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9499;
 wire u6_rem_96_22_Y_u6_div_90_17_n_95;
 wire u6_rem_96_22_Y_u6_div_90_17_n_950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9500;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9501;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9502;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9503;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9504;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9505;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9506;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9507;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9509;
 wire u6_rem_96_22_Y_u6_div_90_17_n_951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9510;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9511;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9512;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9513;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9514;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9515;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9516;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9517;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9518;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9519;
 wire u6_rem_96_22_Y_u6_div_90_17_n_952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9520;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9521;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9522;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9523;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9524;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9525;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9526;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9527;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9528;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9529;
 wire u6_rem_96_22_Y_u6_div_90_17_n_953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9530;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9531;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9532;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9533;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9534;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9535;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9536;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9537;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9538;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9539;
 wire u6_rem_96_22_Y_u6_div_90_17_n_954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9540;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9541;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9542;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9543;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9544;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9545;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9546;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9547;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9548;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9549;
 wire u6_rem_96_22_Y_u6_div_90_17_n_955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9550;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9551;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9552;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9553;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9554;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9555;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9556;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9557;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9558;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9559;
 wire u6_rem_96_22_Y_u6_div_90_17_n_956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9560;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9561;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9562;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9563;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9564;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9565;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9566;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9567;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9568;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9569;
 wire u6_rem_96_22_Y_u6_div_90_17_n_957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9570;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9571;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9572;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9573;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9574;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9575;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9576;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9577;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9578;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9579;
 wire u6_rem_96_22_Y_u6_div_90_17_n_958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9580;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9581;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9582;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9583;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9584;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9585;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9586;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9587;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9588;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9589;
 wire u6_rem_96_22_Y_u6_div_90_17_n_959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9590;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9591;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9592;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9593;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9594;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9595;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9596;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9597;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9598;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9599;
 wire u6_rem_96_22_Y_u6_div_90_17_n_96;
 wire u6_rem_96_22_Y_u6_div_90_17_n_960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9600;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9601;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9602;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9603;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9604;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9605;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9606;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9607;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9608;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9609;
 wire u6_rem_96_22_Y_u6_div_90_17_n_961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9610;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9611;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9612;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9613;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9614;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9615;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9616;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9617;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9618;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9619;
 wire u6_rem_96_22_Y_u6_div_90_17_n_962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9620;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9621;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9622;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9623;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9624;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9625;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9626;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9627;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9628;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9629;
 wire u6_rem_96_22_Y_u6_div_90_17_n_963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9630;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9631;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9632;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9633;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9634;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9635;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9636;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9637;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9638;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9639;
 wire u6_rem_96_22_Y_u6_div_90_17_n_964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9640;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9641;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9642;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9643;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9644;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9645;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9647;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9648;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9649;
 wire u6_rem_96_22_Y_u6_div_90_17_n_965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9650;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9651;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9652;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9653;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9654;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9655;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9656;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9657;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9658;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9659;
 wire u6_rem_96_22_Y_u6_div_90_17_n_966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9660;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9661;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9662;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9663;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9664;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9665;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9666;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9667;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9668;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9669;
 wire u6_rem_96_22_Y_u6_div_90_17_n_967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9670;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9671;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9672;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9673;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9674;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9675;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9676;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9677;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9678;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9679;
 wire u6_rem_96_22_Y_u6_div_90_17_n_968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9680;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9681;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9683;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9684;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9685;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9686;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9687;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9688;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9689;
 wire u6_rem_96_22_Y_u6_div_90_17_n_969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9690;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9691;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9692;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9693;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9694;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9695;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9696;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9697;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9698;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9699;
 wire u6_rem_96_22_Y_u6_div_90_17_n_970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9700;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9701;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9702;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9703;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9704;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9705;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9706;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9707;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9708;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9709;
 wire u6_rem_96_22_Y_u6_div_90_17_n_971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9710;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9711;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9712;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9713;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9714;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9715;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9716;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9717;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9718;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9719;
 wire u6_rem_96_22_Y_u6_div_90_17_n_972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9720;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9721;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9722;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9723;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9724;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9725;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9726;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9727;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9728;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9729;
 wire u6_rem_96_22_Y_u6_div_90_17_n_973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9730;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9731;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9732;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9733;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9734;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9735;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9736;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9737;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9739;
 wire u6_rem_96_22_Y_u6_div_90_17_n_974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9740;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9741;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9742;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9743;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9744;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9745;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9746;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9747;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9748;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9749;
 wire u6_rem_96_22_Y_u6_div_90_17_n_975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9750;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9751;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9752;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9753;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9754;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9755;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9756;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9757;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9758;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9759;
 wire u6_rem_96_22_Y_u6_div_90_17_n_976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9760;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9761;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9762;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9763;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9764;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9765;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9766;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9768;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9769;
 wire u6_rem_96_22_Y_u6_div_90_17_n_977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9770;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9771;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9772;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9773;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9774;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9775;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9776;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9777;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9778;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9779;
 wire u6_rem_96_22_Y_u6_div_90_17_n_978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9780;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9781;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9782;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9783;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9784;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9785;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9786;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9787;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9788;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9789;
 wire u6_rem_96_22_Y_u6_div_90_17_n_979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9790;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9791;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9792;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9793;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9794;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9795;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9796;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9797;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9798;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9799;
 wire u6_rem_96_22_Y_u6_div_90_17_n_98;
 wire u6_rem_96_22_Y_u6_div_90_17_n_980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9801;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9802;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9803;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9804;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9805;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9806;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9807;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9808;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9809;
 wire u6_rem_96_22_Y_u6_div_90_17_n_981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9810;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9811;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9812;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9813;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9814;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9815;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9816;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9817;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9818;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9819;
 wire u6_rem_96_22_Y_u6_div_90_17_n_982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9820;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9821;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9822;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9823;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9824;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9825;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9826;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9827;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9828;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9829;
 wire u6_rem_96_22_Y_u6_div_90_17_n_983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9830;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9831;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9832;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9833;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9834;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9835;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9836;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9837;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9838;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9839;
 wire u6_rem_96_22_Y_u6_div_90_17_n_984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9840;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9841;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9842;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9843;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9844;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9845;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9846;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9847;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9848;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9849;
 wire u6_rem_96_22_Y_u6_div_90_17_n_985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9850;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9851;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9852;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9853;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9854;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9855;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9856;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9857;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9858;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9859;
 wire u6_rem_96_22_Y_u6_div_90_17_n_986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9860;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9861;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9862;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9863;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9864;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9865;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9866;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9867;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9868;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9869;
 wire u6_rem_96_22_Y_u6_div_90_17_n_987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9870;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9871;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9872;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9873;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9874;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9875;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9876;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9877;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9878;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9879;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9880;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9881;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9882;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9883;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9884;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9885;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9886;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9887;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9888;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9889;
 wire u6_rem_96_22_Y_u6_div_90_17_n_989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9890;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9891;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9892;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9893;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9894;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9895;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9896;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9897;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9898;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9899;
 wire u6_rem_96_22_Y_u6_div_90_17_n_99;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9900;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9901;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9902;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9903;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9904;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9905;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9906;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9908;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9909;
 wire u6_rem_96_22_Y_u6_div_90_17_n_991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9910;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9911;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9912;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9913;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9914;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9915;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9916;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9917;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9918;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9919;
 wire u6_rem_96_22_Y_u6_div_90_17_n_992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9920;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9921;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9923;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9924;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9925;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9926;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9927;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9928;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9929;
 wire u6_rem_96_22_Y_u6_div_90_17_n_993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9930;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9931;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9932;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9933;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9934;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9935;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9936;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9937;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9938;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9939;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9940;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9941;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9942;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9943;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9944;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9945;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9946;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9947;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9948;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9949;
 wire u6_rem_96_22_Y_u6_div_90_17_n_995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9950;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9951;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9952;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9953;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9954;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9955;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9956;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9957;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9958;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9959;
 wire u6_rem_96_22_Y_u6_div_90_17_n_996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9960;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9961;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9962;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9963;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9964;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9965;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9966;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9967;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9968;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9969;
 wire u6_rem_96_22_Y_u6_div_90_17_n_997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9970;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9971;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9972;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9973;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9974;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9975;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9976;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9977;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9978;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9979;
 wire u6_rem_96_22_Y_u6_div_90_17_n_998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9980;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9981;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9982;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9983;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9984;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9985;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9986;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9987;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9988;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9989;
 wire u6_rem_96_22_Y_u6_div_90_17_n_999;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9990;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9991;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9992;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9993;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9994;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9995;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9996;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9997;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9998;
 wire u6_rem_96_22_Y_u6_div_90_17_n_9999;
 wire [4:0] div_opa_ldz_r1;
 wire [4:0] div_opa_ldz_r2;
 wire [7:0] exp_fasu;
 wire [7:0] exp_mul;
 wire [1:0] exp_ovf;
 wire [1:0] exp_ovf_r;
 wire [7:0] exp_r;
 wire [2:0] fpu_op_r1;
 wire [2:0] fpu_op_r2;
 wire [2:0] fpu_op_r3;
 wire [47:0] fract_denorm;
 wire [47:0] fract_i2f;
 wire [27:0] fract_out_q;
 wire [26:0] fracta;
 wire [23:0] fracta_mul;
 wire [26:0] fractb;
 wire [23:0] fractb_mul;
 wire [31:0] opa_r;
 wire [30:0] opa_r1;
 wire [31:0] opb_r;
 wire [47:0] prod;
 wire [49:0] quo;
 wire [23:0] remainder;
 wire [1:0] rmode_r1;
 wire [1:0] rmode_r2;
 wire [1:0] rmode_r3;
 wire [7:0] u1_exp_large;
 wire [26:0] u1_fracta_s;
 wire [26:0] u1_fractb_s;
 wire [1:0] u2_exp_ovf_d;
 wire [7:0] u2_exp_tmp1;
 wire [7:0] u4_exp_div;
 wire [7:0] u4_exp_out;
 wire [22:0] u4_fract_out;
 wire [23:0] u4_fract_out_pl1;
 wire [24:0] u4_fract_trunc;
 wire [47:0] u5_prod1;
 wire [49:0] u6_quo1;
 wire [23:0] u6_remainder;
 wire [2:0] underflow_fmul_d;
 wire [2:0] underflow_fmul_r;

 DFFHQNx1_ASAP7_75t_R div_by_zero_reg (.CLK(clk),
    .D(n_259),
    .QN(div_by_zero));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r1_reg[0]  (.CLK(clk),
    .D(n_1071),
    .QN(div_opa_ldz_r1[0]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r1_reg[1]  (.CLK(clk),
    .D(n_1072),
    .QN(div_opa_ldz_r1[1]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r1_reg[2]  (.CLK(clk),
    .D(n_1079),
    .QN(div_opa_ldz_r1[2]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r1_reg[3]  (.CLK(clk),
    .D(n_1075),
    .QN(div_opa_ldz_r1[3]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r1_reg[4]  (.CLK(clk),
    .D(n_1058),
    .QN(div_opa_ldz_r1[4]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r2_reg[0]  (.CLK(clk),
    .D(n_1087),
    .QN(div_opa_ldz_r2[0]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r2_reg[1]  (.CLK(clk),
    .D(n_1086),
    .QN(div_opa_ldz_r2[1]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r2_reg[2]  (.CLK(clk),
    .D(n_1120),
    .QN(div_opa_ldz_r2[2]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r2_reg[3]  (.CLK(clk),
    .D(n_1121),
    .QN(div_opa_ldz_r2[3]));
 DFFHQNx1_ASAP7_75t_R \div_opa_ldz_r2_reg[4]  (.CLK(clk),
    .D(n_1074),
    .QN(div_opa_ldz_r2[4]));
 HB1xp67_ASAP7_75t_R drc_buf_sp234637 (.A(fracta_mul[23]),
    .Y(n_13883));
 HB1xp67_ASAP7_75t_R drc_buf_sp234638 (.A(fracta_mul[23]),
    .Y(n_13884));
 HB1xp67_ASAP7_75t_R drc_buf_sp234673 (.A(n_13919),
    .Y(n_13920));
 HB1xp67_ASAP7_75t_R drc_buf_sp234674 (.A(u4_n_1362),
    .Y(n_13919));
 HB1xp67_ASAP7_75t_R drc_buf_sp234698 (.A(exp_r[5]),
    .Y(n_13946));
 HB1xp67_ASAP7_75t_R drc_buf_sp234723 (.A(exp_r[0]),
    .Y(n_13972));
 HB1xp67_ASAP7_75t_R drc_buf_sp234731 (.A(u2_n_606),
    .Y(n_13981));
 INVx2_ASAP7_75t_SL drc_bufs36417 (.A(n_2944),
    .Y(n_2940));
 INVx2_ASAP7_75t_L drc_bufs36418 (.A(n_2943),
    .Y(n_2944));
 INVxp33_ASAP7_75t_R drc_bufs37394 (.A(n_9),
    .Y(n_12));
 INVxp33_ASAP7_75t_R drc_bufs37395 (.A(n_9),
    .Y(n_11));
 INVxp33_ASAP7_75t_R drc_bufs37396 (.A(n_9),
    .Y(n_10));
 INVxp33_ASAP7_75t_R drc_bufs37407 (.A(n_13),
    .Y(n_8));
 INVxp33_ASAP7_75t_R drc_bufs37415 (.A(u1_n_1066),
    .Y(n_7));
 INVxp33_ASAP7_75t_R drc_bufs37423 (.A(n_4),
    .Y(n_5));
 INVxp33_ASAP7_75t_R drc_bufs37424 (.A(n_541),
    .Y(n_4));
 INVxp33_ASAP7_75t_R drc_bufs37431 (.A(n_15),
    .Y(n_3));
 INVxp33_ASAP7_75t_R drc_bufs37432 (.A(n_539),
    .Y(n_15));
 INVxp33_ASAP7_75t_R drc_bufs37439 (.A(n_14),
    .Y(n_2));
 INVxp33_ASAP7_75t_R drc_bufs37440 (.A(n_538),
    .Y(n_14));
 INVxp33_ASAP7_75t_R drc_bufs37447 (.A(u1_n_1066),
    .Y(n_1));
 INVxp33_ASAP7_75t_R drc_bufs44686 (.A(n_3497),
    .Y(n_681));
 INVxp33_ASAP7_75t_R drc_bufs44687 (.A(n_3497),
    .Y(n_680));
 INVxp33_ASAP7_75t_R drc_bufs44688 (.A(n_3497),
    .Y(n_679));
 INVxp33_ASAP7_75t_R drc_bufs44689 (.A(n_682),
    .Y(n_3497));
 INVxp33_ASAP7_75t_R drc_bufs44699 (.A(n_675),
    .Y(n_678));
 INVxp33_ASAP7_75t_R drc_bufs44700 (.A(n_675),
    .Y(n_677));
 INVxp33_ASAP7_75t_R drc_bufs44701 (.A(n_675),
    .Y(n_676));
 INVxp33_ASAP7_75t_R drc_bufs44702 (.A(n_1059),
    .Y(n_675));
 INVxp33_ASAP7_75t_R drc_bufs44711 (.A(n_3850),
    .Y(n_674));
 INVxp33_ASAP7_75t_R drc_bufs44712 (.A(n_3850),
    .Y(n_23));
 INVxp33_ASAP7_75t_R drc_bufs44713 (.A(n_3850),
    .Y(n_672));
 INVxp33_ASAP7_75t_R drc_bufs44714 (.A(n_3850),
    .Y(n_671));
 INVxp33_ASAP7_75t_R drc_bufs44721 (.A(n_691),
    .Y(n_670));
 INVxp67_ASAP7_75t_R drc_bufs44722 (.A(n_690),
    .Y(n_691));
 INVxp33_ASAP7_75t_R drc_bufs44728 (.A(n_668),
    .Y(n_669));
 INVxp33_ASAP7_75t_R drc_bufs44729 (.A(n_1432),
    .Y(n_668));
 INVxp33_ASAP7_75t_R drc_bufs44735 (.A(n_666),
    .Y(n_667));
 INVxp33_ASAP7_75t_R drc_bufs44736 (.A(n_1433),
    .Y(n_666));
 INVxp33_ASAP7_75t_R drc_bufs44743 (.A(n_1150),
    .Y(n_689));
 INVxp33_ASAP7_75t_R drc_bufs44750 (.A(n_1218),
    .Y(n_693));
 INVxp33_ASAP7_75t_R drc_bufs44755 (.A(n_3498),
    .Y(n_653));
 INVxp33_ASAP7_75t_R drc_bufs44756 (.A(n_3498),
    .Y(n_652));
 INVxp33_ASAP7_75t_R drc_bufs44763 (.A(n_664),
    .Y(n_665));
 INVxp33_ASAP7_75t_R drc_bufs44764 (.A(n_1060),
    .Y(n_664));
 INVxp33_ASAP7_75t_R drc_bufs44769 (.A(n_688),
    .Y(n_663));
 INVxp33_ASAP7_75t_R drc_bufs44770 (.A(n_688),
    .Y(n_686));
 INVxp33_ASAP7_75t_R drc_bufs44771 (.A(n_1150),
    .Y(n_688));
 INVxp33_ASAP7_75t_R drc_bufs44777 (.A(n_661),
    .Y(n_662));
 INVxp33_ASAP7_75t_R drc_bufs44778 (.A(n_1443),
    .Y(n_661));
 INVxp33_ASAP7_75t_R drc_bufs44784 (.A(n_687),
    .Y(n_660));
 INVxp67_ASAP7_75t_R drc_bufs44785 (.A(n_686),
    .Y(n_687));
 INVxp33_ASAP7_75t_R drc_bufs44791 (.A(n_699),
    .Y(n_659));
 INVxp33_ASAP7_75t_R drc_bufs44792 (.A(n_1436),
    .Y(n_699));
 INVxp33_ASAP7_75t_R drc_bufs44798 (.A(n_697),
    .Y(n_658));
 INVxp33_ASAP7_75t_R drc_bufs44799 (.A(n_1290),
    .Y(n_697));
 INVxp33_ASAP7_75t_R drc_bufs44805 (.A(n_1153),
    .Y(n_690));
 INVxp33_ASAP7_75t_R drc_bufs44811 (.A(u1_n_853),
    .Y(n_657));
 INVxp33_ASAP7_75t_R drc_bufs44813 (.A(n_693),
    .Y(u1_n_853));
 HB1xp67_ASAP7_75t_R drc_bufs44829 (.A(n_1435),
    .Y(n_655));
 HB1xp67_ASAP7_75t_R drc_bufs44835 (.A(n_1291),
    .Y(n_654));
 INVxp33_ASAP7_75t_R drc_bufs53377 (.A(n_1843),
    .Y(n_1823));
 INVxp33_ASAP7_75t_R drc_bufs53378 (.A(n_2595),
    .Y(n_1843));
 INVxp33_ASAP7_75t_R drc_bufs53383 (.A(n_2592),
    .Y(n_1822));
 INVxp33_ASAP7_75t_R drc_bufs53384 (.A(n_2592),
    .Y(n_1821));
 INVxp33_ASAP7_75t_R drc_bufs53391 (.A(n_1824),
    .Y(n_1820));
 INVxp33_ASAP7_75t_R drc_bufs53392 (.A(n_2233),
    .Y(n_1824));
 INVxp33_ASAP7_75t_R drc_bufs53398 (.A(n_1818),
    .Y(n_1819));
 INVxp33_ASAP7_75t_R drc_bufs53399 (.A(n_2235),
    .Y(n_1818));
 INVxp33_ASAP7_75t_R drc_bufs53405 (.A(n_2233),
    .Y(n_1817));
 HB1xp67_ASAP7_75t_R drc_bufs53418 (.A(n_1832),
    .Y(n_1830));
 HB1xp67_ASAP7_75t_R drc_bufs53470 (.A(n_2525),
    .Y(n_1816));
 DFFHQNx1_ASAP7_75t_R \exp_ovf_r_reg[0]  (.CLK(clk),
    .D(n_1289),
    .QN(exp_ovf_r[0]));
 DFFHQNx1_ASAP7_75t_R \exp_ovf_r_reg[1]  (.CLK(clk),
    .D(n_1274),
    .QN(exp_ovf_r[1]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[0]  (.CLK(clk),
    .D(n_635),
    .QN(exp_r[0]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[1]  (.CLK(clk),
    .D(n_633),
    .QN(exp_r[1]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[2]  (.CLK(clk),
    .D(n_632),
    .QN(exp_r[2]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[3]  (.CLK(clk),
    .D(n_637),
    .QN(exp_r[3]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[4]  (.CLK(clk),
    .D(n_638),
    .QN(exp_r[4]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[5]  (.CLK(clk),
    .D(n_639),
    .QN(exp_r[5]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[6]  (.CLK(clk),
    .D(n_636),
    .QN(exp_r[6]));
 DFFHQNx1_ASAP7_75t_R \exp_r_reg[7]  (.CLK(clk),
    .D(n_634),
    .QN(exp_r[7]));
 DFFHQNx1_ASAP7_75t_R fasu_op_r1_reg (.CLK(clk),
    .D(u3_sub_52_45_Y_add_52_31_n_841),
    .QN(fasu_op_r1));
 DFFHQNx1_ASAP7_75t_R fasu_op_r2_reg (.CLK(clk),
    .D(n_2043),
    .QN(fasu_op_r2));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r1_reg[0]  (.CLK(clk),
    .D(n_3287),
    .QN(fpu_op_r1[0]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r1_reg[1]  (.CLK(clk),
    .D(n_834),
    .QN(fpu_op_r1[1]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r1_reg[2]  (.CLK(clk),
    .D(n_822),
    .QN(fpu_op_r1[2]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r2_reg[0]  (.CLK(clk),
    .D(n_726),
    .QN(fpu_op_r2[0]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r2_reg[1]  (.CLK(clk),
    .D(n_64),
    .QN(fpu_op_r2[1]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r2_reg[2]  (.CLK(clk),
    .D(n_56),
    .QN(fpu_op_r2[2]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r3_reg[0]  (.CLK(clk),
    .D(n_875),
    .QN(fpu_op_r3[0]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r3_reg[1]  (.CLK(clk),
    .D(n_801),
    .QN(fpu_op_r3[1]));
 DFFHQNx1_ASAP7_75t_R \fpu_op_r3_reg[2]  (.CLK(clk),
    .D(n_727),
    .QN(fpu_op_r3[2]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[0]  (.CLK(n_1602),
    .D(n_1098),
    .Q(fract_denorm[0]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[10]  (.CLK(n_1602),
    .D(n_1534),
    .Q(fract_denorm[10]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[11]  (.CLK(n_1602),
    .D(n_1533),
    .Q(fract_denorm[11]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[12]  (.CLK(n_1602),
    .D(n_1532),
    .Q(fract_denorm[12]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[13]  (.CLK(n_1602),
    .D(n_1531),
    .Q(fract_denorm[13]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[14]  (.CLK(n_1602),
    .D(n_1530),
    .Q(fract_denorm[14]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[15]  (.CLK(n_1602),
    .D(n_1529),
    .Q(fract_denorm[15]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[16]  (.CLK(n_1602),
    .D(n_1528),
    .Q(fract_denorm[16]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[17]  (.CLK(n_1602),
    .D(n_651),
    .Q(fract_denorm[17]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[18]  (.CLK(n_1602),
    .D(n_650),
    .Q(fract_denorm[18]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[19]  (.CLK(n_1602),
    .D(n_649),
    .Q(fract_denorm[19]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[1]  (.CLK(n_1602),
    .D(n_1527),
    .Q(fract_denorm[1]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[20]  (.CLK(n_1602),
    .D(n_1560),
    .Q(fract_denorm[20]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[21]  (.CLK(n_1602),
    .D(n_1561),
    .Q(fract_denorm[21]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[22]  (.CLK(n_1602),
    .D(n_1562),
    .Q(fract_denorm[22]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[23]  (.CLK(n_1602),
    .D(n_1563),
    .Q(fract_denorm[23]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[24]  (.CLK(n_1602),
    .D(n_1564),
    .Q(fract_denorm[24]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[25]  (.CLK(n_1602),
    .D(n_1565),
    .Q(fract_denorm[25]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[26]  (.CLK(n_1602),
    .D(n_1566),
    .Q(fract_denorm[26]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[27]  (.CLK(n_1602),
    .D(n_1559),
    .Q(fract_denorm[27]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[28]  (.CLK(n_1602),
    .D(n_1558),
    .Q(fract_denorm[28]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[29]  (.CLK(n_1602),
    .D(n_1557),
    .Q(fract_denorm[29]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[2]  (.CLK(n_1602),
    .D(n_1526),
    .Q(fract_denorm[2]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[30]  (.CLK(n_1602),
    .D(n_1556),
    .Q(fract_denorm[30]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[31]  (.CLK(n_1602),
    .D(n_1555),
    .Q(fract_denorm[31]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[32]  (.CLK(n_1602),
    .D(n_1554),
    .Q(fract_denorm[32]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[33]  (.CLK(n_1602),
    .D(n_1553),
    .Q(fract_denorm[33]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[34]  (.CLK(n_1602),
    .D(n_1552),
    .Q(fract_denorm[34]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[35]  (.CLK(n_1602),
    .D(n_1551),
    .Q(fract_denorm[35]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[36]  (.CLK(n_1602),
    .D(n_1550),
    .Q(fract_denorm[36]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[37]  (.CLK(n_1602),
    .D(n_1549),
    .Q(fract_denorm[37]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[38]  (.CLK(n_1602),
    .D(n_1548),
    .Q(fract_denorm[38]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[39]  (.CLK(n_1602),
    .D(n_1547),
    .Q(fract_denorm[39]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[3]  (.CLK(n_1602),
    .D(n_1525),
    .Q(fract_denorm[3]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[40]  (.CLK(n_1602),
    .D(n_1546),
    .Q(fract_denorm[40]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[41]  (.CLK(n_1602),
    .D(n_1545),
    .Q(fract_denorm[41]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[42]  (.CLK(n_1602),
    .D(n_1544),
    .Q(fract_denorm[42]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[43]  (.CLK(n_1602),
    .D(n_1574),
    .Q(fract_denorm[43]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[44]  (.CLK(n_1602),
    .D(n_1543),
    .Q(fract_denorm[44]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[45]  (.CLK(n_1602),
    .D(n_1573),
    .Q(fract_denorm[45]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[46]  (.CLK(n_1602),
    .D(n_1542),
    .Q(fract_denorm[46]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[47]  (.CLK(n_1602),
    .D(n_1541),
    .Q(fract_denorm[47]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[4]  (.CLK(n_1602),
    .D(n_1524),
    .Q(fract_denorm[4]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[5]  (.CLK(n_1602),
    .D(n_1523),
    .Q(fract_denorm[5]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[6]  (.CLK(n_1602),
    .D(n_1518),
    .Q(fract_denorm[6]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[7]  (.CLK(n_1602),
    .D(n_1537),
    .Q(fract_denorm[7]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[8]  (.CLK(n_1602),
    .D(n_1536),
    .Q(fract_denorm[8]));
 DHLx1_ASAP7_75t_R \fract_denorm_reg[9]  (.CLK(n_1602),
    .D(n_1535),
    .Q(fract_denorm[9]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[0]  (.CLK(clk),
    .D(n_1033),
    .QN(fract_i2f[0]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[10]  (.CLK(clk),
    .D(n_1460),
    .QN(fract_i2f[10]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[11]  (.CLK(clk),
    .D(n_1449),
    .QN(fract_i2f[11]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[12]  (.CLK(clk),
    .D(n_1454),
    .QN(fract_i2f[12]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[13]  (.CLK(clk),
    .D(n_1453),
    .QN(fract_i2f[13]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[14]  (.CLK(clk),
    .D(n_1452),
    .QN(fract_i2f[14]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[15]  (.CLK(clk),
    .D(n_1451),
    .QN(fract_i2f[15]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[16]  (.CLK(clk),
    .D(n_1450),
    .QN(fract_i2f[16]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[17]  (.CLK(clk),
    .D(n_1466),
    .QN(fract_i2f[17]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[18]  (.CLK(clk),
    .D(n_1472),
    .QN(fract_i2f[18]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[19]  (.CLK(clk),
    .D(n_1470),
    .QN(fract_i2f[19]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[1]  (.CLK(clk),
    .D(n_1444),
    .QN(fract_i2f[1]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[20]  (.CLK(clk),
    .D(n_1469),
    .QN(fract_i2f[20]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[21]  (.CLK(clk),
    .D(n_1471),
    .QN(fract_i2f[21]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[22]  (.CLK(clk),
    .D(n_1468),
    .QN(fract_i2f[22]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[23]  (.CLK(clk),
    .D(n_1467),
    .QN(fract_i2f[23]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[24]  (.CLK(clk),
    .D(n_1496),
    .QN(fract_i2f[24]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[25]  (.CLK(clk),
    .D(n_1495),
    .QN(fract_i2f[25]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[26]  (.CLK(clk),
    .D(n_1494),
    .QN(fract_i2f[26]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[27]  (.CLK(clk),
    .D(n_1493),
    .QN(fract_i2f[27]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[28]  (.CLK(clk),
    .D(n_1492),
    .QN(fract_i2f[28]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[29]  (.CLK(clk),
    .D(n_1491),
    .QN(fract_i2f[29]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[2]  (.CLK(clk),
    .D(n_1464),
    .QN(fract_i2f[2]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[30]  (.CLK(clk),
    .D(n_1490),
    .QN(fract_i2f[30]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[31]  (.CLK(clk),
    .D(n_1489),
    .QN(fract_i2f[31]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[32]  (.CLK(clk),
    .D(n_1488),
    .QN(fract_i2f[32]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[33]  (.CLK(clk),
    .D(n_1487),
    .QN(fract_i2f[33]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[34]  (.CLK(clk),
    .D(n_1486),
    .QN(fract_i2f[34]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[35]  (.CLK(clk),
    .D(n_1485),
    .QN(fract_i2f[35]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[36]  (.CLK(clk),
    .D(n_1484),
    .QN(fract_i2f[36]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[37]  (.CLK(clk),
    .D(n_1483),
    .QN(fract_i2f[37]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[38]  (.CLK(clk),
    .D(n_1482),
    .QN(fract_i2f[38]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[39]  (.CLK(clk),
    .D(n_1481),
    .QN(fract_i2f[39]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[3]  (.CLK(clk),
    .D(n_1463),
    .QN(fract_i2f[3]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[40]  (.CLK(clk),
    .D(n_1480),
    .QN(fract_i2f[40]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[41]  (.CLK(clk),
    .D(n_1479),
    .QN(fract_i2f[41]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[42]  (.CLK(clk),
    .D(n_1478),
    .QN(fract_i2f[42]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[43]  (.CLK(clk),
    .D(n_1477),
    .QN(fract_i2f[43]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[44]  (.CLK(clk),
    .D(n_1476),
    .QN(fract_i2f[44]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[45]  (.CLK(clk),
    .D(n_1475),
    .QN(fract_i2f[45]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[46]  (.CLK(clk),
    .D(n_1474),
    .QN(fract_i2f[46]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[47]  (.CLK(clk),
    .D(n_1473),
    .QN(fract_i2f[47]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[4]  (.CLK(clk),
    .D(n_1462),
    .QN(fract_i2f[4]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[5]  (.CLK(clk),
    .D(n_1465),
    .QN(fract_i2f[5]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[6]  (.CLK(clk),
    .D(n_1459),
    .QN(fract_i2f[6]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[7]  (.CLK(clk),
    .D(n_1458),
    .QN(fract_i2f[7]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[8]  (.CLK(clk),
    .D(n_1457),
    .QN(fract_i2f[8]));
 DFFHQNx1_ASAP7_75t_R \fract_i2f_reg[9]  (.CLK(clk),
    .D(n_1456),
    .QN(fract_i2f[9]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[0]  (.CLK(clk),
    .D(n_751),
    .QN(fract_out_q[0]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[10]  (.CLK(clk),
    .D(n_14497),
    .QN(fract_out_q[10]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[11]  (.CLK(clk),
    .D(n_14515),
    .QN(fract_out_q[11]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[12]  (.CLK(clk),
    .D(n_14499),
    .QN(fract_out_q[12]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[13]  (.CLK(clk),
    .D(n_14498),
    .QN(fract_out_q[13]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[14]  (.CLK(clk),
    .D(n_14508),
    .QN(fract_out_q[14]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[15]  (.CLK(clk),
    .D(n_14504),
    .QN(fract_out_q[15]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[16]  (.CLK(clk),
    .D(n_14505),
    .QN(fract_out_q[16]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[17]  (.CLK(clk),
    .D(n_14514),
    .QN(fract_out_q[17]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[18]  (.CLK(clk),
    .D(n_14506),
    .QN(fract_out_q[18]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[19]  (.CLK(clk),
    .D(n_14507),
    .QN(fract_out_q[19]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[1]  (.CLK(clk),
    .D(n_14258),
    .QN(fract_out_q[1]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[20]  (.CLK(clk),
    .D(n_14503),
    .QN(fract_out_q[20]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[21]  (.CLK(clk),
    .D(n_14512),
    .QN(fract_out_q[21]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[22]  (.CLK(clk),
    .D(n_14502),
    .QN(fract_out_q[22]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[23]  (.CLK(clk),
    .D(n_14501),
    .QN(fract_out_q[23]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[24]  (.CLK(clk),
    .D(n_14495),
    .QN(fract_out_q[24]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[25]  (.CLK(clk),
    .D(n_14513),
    .QN(fract_out_q[25]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[26]  (.CLK(clk),
    .D(n_14509),
    .QN(fract_out_q[26]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[27]  (.CLK(clk),
    .D(n_14246),
    .QN(fract_out_q[27]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[2]  (.CLK(clk),
    .D(n_14185),
    .QN(fract_out_q[2]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[3]  (.CLK(clk),
    .D(n_14494),
    .QN(fract_out_q[3]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[4]  (.CLK(clk),
    .D(n_14259),
    .QN(fract_out_q[4]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[5]  (.CLK(clk),
    .D(n_14516),
    .QN(fract_out_q[5]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[6]  (.CLK(clk),
    .D(n_14496),
    .QN(fract_out_q[6]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[7]  (.CLK(clk),
    .D(n_14500),
    .QN(fract_out_q[7]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[8]  (.CLK(clk),
    .D(n_14511),
    .QN(fract_out_q[8]));
 DFFHQNx1_ASAP7_75t_R \fract_out_q_reg[9]  (.CLK(clk),
    .D(n_14510),
    .QN(fract_out_q[9]));
 INVxp33_ASAP7_75t_R g100 (.A(u6_remainder[15]),
    .Y(n_14071));
 INVxp33_ASAP7_75t_R g106 (.A(u6_remainder[16]),
    .Y(n_14072));
 INVxp33_ASAP7_75t_R g110 (.A(u6_remainder[8]),
    .Y(n_14064));
 INVxp33_ASAP7_75t_R g112 (.A(u6_remainder[17]),
    .Y(n_14073));
 INVxp33_ASAP7_75t_R g116 (.A(u6_remainder[18]),
    .Y(n_14074));
 INVxp33_ASAP7_75t_R g120 (.A(u6_remainder[4]),
    .Y(n_14060));
 INVxp33_ASAP7_75t_R g122 (.A(u6_remainder[9]),
    .Y(n_14065));
 INVxp33_ASAP7_75t_R g124 (.A(u6_remainder[19]),
    .Y(n_14075));
 INVxp33_ASAP7_75t_R g128 (.A(u6_remainder[20]),
    .Y(n_14076));
 INVxp33_ASAP7_75t_R g132 (.A(u6_remainder[10]),
    .Y(n_14066));
 INVxp33_ASAP7_75t_R g134 (.A(u6_remainder[21]),
    .Y(n_14077));
 INVxp33_ASAP7_75t_R g138 (.A(u6_remainder[22]),
    .Y(n_14078));
 INVxp33_ASAP7_75t_R g142 (.A(u6_remainder[2]),
    .Y(n_14058));
 INVxp33_ASAP7_75t_R g144 (.A(u6_remainder[5]),
    .Y(n_14061));
 INVxp33_ASAP7_75t_R g146 (.A(u6_remainder[11]),
    .Y(n_14067));
 INVxp33_ASAP7_75t_R g148 (.A(u6_remainder[23]),
    .Y(n_14079));
 INVxp33_ASAP7_75t_R g15 (.A(opa[16]),
    .Y(n_14167));
 INVxp33_ASAP7_75t_R g152 (.A(n_14081),
    .Y(n_14082));
 INVxp33_ASAP7_75t_R g156 (.A(u6_remainder[12]),
    .Y(n_14068));
 INVxp33_ASAP7_75t_R g158 (.A(n_14085),
    .Y(n_14086));
 INVxp33_ASAP7_75t_R g16 (.A(opa[15]),
    .Y(n_14165));
 INVxp33_ASAP7_75t_R g165 (.A(u6_remainder[6]),
    .Y(n_14062));
 INVxp33_ASAP7_75t_R g167 (.A(u6_remainder[13]),
    .Y(n_14069));
 INVxp33_ASAP7_75t_R g17 (.A(opa[18]),
    .Y(n_14171));
 INVxp33_ASAP7_75t_R g175 (.A(u6_remainder[14]),
    .Y(n_14070));
 INVxp33_ASAP7_75t_R g18 (.A(opa[19]),
    .Y(n_14173));
 INVxp67_ASAP7_75t_R g183 (.A(u6_n_126),
    .Y(n_14054));
 INVxp33_ASAP7_75t_R g184 (.A(opb[22]),
    .Y(n_14163));
 INVxp33_ASAP7_75t_R g185 (.A(u6_n_76),
    .Y(n_14080));
 INVxp33_ASAP7_75t_R g187 (.A(opa[2]),
    .Y(n_14091));
 INVxp33_ASAP7_75t_R g188 (.A(opa[3]),
    .Y(n_14093));
 INVxp33_ASAP7_75t_R g189 (.A(opa[5]),
    .Y(n_14097));
 INVxp33_ASAP7_75t_R g19 (.A(opb[2]),
    .Y(n_14177));
 INVxp33_ASAP7_75t_R g190 (.A(opa[6]),
    .Y(n_14099));
 INVxp33_ASAP7_75t_R g191 (.A(opa[11]),
    .Y(n_14109));
 INVxp33_ASAP7_75t_R g192 (.A(opa[12]),
    .Y(n_14111));
 INVxp33_ASAP7_75t_R g193 (.A(opa[14]),
    .Y(n_14115));
 INVxp33_ASAP7_75t_R g194 (.A(opa[20]),
    .Y(n_14117));
 INVxp33_ASAP7_75t_R g195 (.A(opb[1]),
    .Y(n_14123));
 INVxp33_ASAP7_75t_R g196 (.A(opb[3]),
    .Y(n_14125));
 INVxp33_ASAP7_75t_R g197 (.A(opb[5]),
    .Y(n_14129));
 INVxp33_ASAP7_75t_R g198 (.A(opb[6]),
    .Y(n_14131));
 INVxp33_ASAP7_75t_R g199 (.A(opb[10]),
    .Y(n_14139));
 O2A1O1Ixp33_ASAP7_75t_SL g2 (.A1(n_3146),
    .A2(n_3137),
    .B(n_2940),
    .C(n_3200),
    .Y(n_13834));
 INVxp33_ASAP7_75t_R g20 (.A(opa[17]),
    .Y(n_14169));
 INVxp33_ASAP7_75t_R g200 (.A(opb[11]),
    .Y(n_14141));
 INVxp33_ASAP7_75t_R g201 (.A(opb[13]),
    .Y(n_14145));
 INVxp33_ASAP7_75t_R g202 (.A(opb[14]),
    .Y(n_14147));
 INVxp33_ASAP7_75t_R g203 (.A(opb[17]),
    .Y(n_14153));
 INVxp33_ASAP7_75t_R g204 (.A(opb[18]),
    .Y(n_14155));
 INVxp33_ASAP7_75t_R g205 (.A(opb[20]),
    .Y(n_14159));
 INVxp33_ASAP7_75t_R g206 (.A(opb[21]),
    .Y(n_14161));
 INVxp33_ASAP7_75t_R g207 (.A(opa[1]),
    .Y(n_14089));
 INVxp33_ASAP7_75t_R g208 (.A(opa[4]),
    .Y(n_14095));
 INVxp33_ASAP7_75t_R g209 (.A(opa[10]),
    .Y(n_14107));
 INVxp33_ASAP7_75t_R g21 (.A(opa[22]),
    .Y(n_14175));
 INVxp33_ASAP7_75t_R g210 (.A(opa[13]),
    .Y(n_14113));
 INVxp33_ASAP7_75t_R g211 (.A(opb[0]),
    .Y(n_14121));
 INVxp33_ASAP7_75t_R g212 (.A(opb[4]),
    .Y(n_14127));
 INVxp33_ASAP7_75t_R g213 (.A(opb[9]),
    .Y(n_14137));
 INVxp33_ASAP7_75t_R g214 (.A(opb[12]),
    .Y(n_14143));
 INVxp33_ASAP7_75t_R g215 (.A(opb[16]),
    .Y(n_14151));
 INVxp33_ASAP7_75t_R g216 (.A(opb[19]),
    .Y(n_14157));
 INVxp33_ASAP7_75t_R g217 (.A(opa[0]),
    .Y(n_14087));
 INVxp33_ASAP7_75t_R g218 (.A(opa[9]),
    .Y(n_14105));
 INVxp33_ASAP7_75t_R g219 (.A(opa[21]),
    .Y(n_14119));
 INVxp33_ASAP7_75t_R g220 (.A(opb[8]),
    .Y(n_14135));
 INVxp33_ASAP7_75t_R g221 (.A(opb[15]),
    .Y(n_14149));
 INVxp33_ASAP7_75t_R g222 (.A(opa[8]),
    .Y(n_14103));
 INVxp33_ASAP7_75t_R g223 (.A(opb[7]),
    .Y(n_14133));
 INVxp33_ASAP7_75t_R g224 (.A(opa[7]),
    .Y(n_14101));
 INVxp33_ASAP7_75t_R g234590 (.A(n_3302),
    .Y(u5_mul_69_18_n_115));
 A2O1A1Ixp33_ASAP7_75t_L g234591 (.A1(n_2953),
    .A2(n_2888),
    .B(n_3163),
    .C(n_2940),
    .Y(n_13835));
 OAI21xp33_ASAP7_75t_SL g234592 (.A1(n_3151),
    .A2(n_3136),
    .B(n_2940),
    .Y(n_13836));
 OAI21xp33_ASAP7_75t_L g234593 (.A1(n_3154),
    .A2(n_3144),
    .B(n_2940),
    .Y(n_13837));
 NOR2xp33_ASAP7_75t_R g234594 (.A(n_2882),
    .B(n_2943),
    .Y(n_13838));
 NAND2xp33_ASAP7_75t_R g234595 (.A(n_76),
    .B(n_14118),
    .Y(n_13839));
 NAND3xp33_ASAP7_75t_R g234596 (.A(exp_r[5]),
    .B(n_2278),
    .C(exp_r[7]),
    .Y(n_13840));
 NOR2xp33_ASAP7_75t_R g234597 (.A(n_13841),
    .B(n_2149),
    .Y(n_13842));
 AOI21xp33_ASAP7_75t_R g234598 (.A1(n_1412),
    .A2(n_1411),
    .B(n_1413),
    .Y(n_13843));
 OAI21xp33_ASAP7_75t_R g234599 (.A1(u2_exp_ovf_d[1]),
    .A2(n_1040),
    .B(opa_r[30]),
    .Y(n_13844));
 AND2x2_ASAP7_75t_R g234600 (.A(n_13846),
    .B(n_425),
    .Y(n_13845));
 NAND3xp33_ASAP7_75t_R g234601 (.A(n_383),
    .B(n_478),
    .C(n_3503),
    .Y(n_13846));
 OA21x2_ASAP7_75t_R g234602 (.A1(n_270),
    .A2(n_3514),
    .B(n_3766),
    .Y(n_13847));
 NAND4xp25_ASAP7_75t_L g234603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_432),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12392),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12383),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .Y(n_13848));
 AOI21xp33_ASAP7_75t_L g234604 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10834),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10769),
    .Y(n_13849));
 MAJx2_ASAP7_75t_SL g234605 (.A(n_13850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .Y(n_13851));
 AO21x1_ASAP7_75t_SL g234606 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7180),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1593),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6931),
    .Y(n_13850));
 MAJx2_ASAP7_75t_SL g234607 (.A(n_13852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6098));
 AOI21xp5_ASAP7_75t_R g234608 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1360),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5865),
    .Y(n_13852));
 MAJx2_ASAP7_75t_R g234611 (.A(n_13856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(n_13857));
 OR2x2_ASAP7_75t_R g234612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .Y(n_13856));
 MAJx2_ASAP7_75t_L g234613 (.A(n_13858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(n_13859));
 NAND2xp5_ASAP7_75t_L g234614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_44),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3642),
    .Y(n_13858));
 MAJx2_ASAP7_75t_L g234615 (.A(n_13860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3372),
    .Y(n_13861));
 OR2x2_ASAP7_75t_SL g234616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3371),
    .Y(n_13860));
 AOI21xp33_ASAP7_75t_R g234617 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_234),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2687),
    .Y(n_13862));
 NOR2xp33_ASAP7_75t_R g234618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .Y(n_13863));
 AND2x2_ASAP7_75t_R g234619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .Y(n_13864));
 NAND2xp33_ASAP7_75t_R g234620 (.A(n_14178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_789),
    .Y(n_13865));
 NOR2xp33_ASAP7_75t_R g234621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .Y(n_13866));
 OAI21xp33_ASAP7_75t_R g234622 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(n_14134),
    .Y(n_13867));
 MAJIxp5_ASAP7_75t_R g234623 (.A(n_13868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(n_13869));
 AOI21xp5_ASAP7_75t_R g234624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5290),
    .Y(n_13868));
 NOR2xp33_ASAP7_75t_R g234780 (.A(opa_r1[0]),
    .B(opa_r1[1]),
    .Y(n_14033));
 AND2x2_ASAP7_75t_R g234882 (.A(exp_ovf_r[0]),
    .B(u4_op_dn),
    .Y(n_14180));
 OA21x2_ASAP7_75t_R g234883 (.A1(n_1681),
    .A2(n_3588),
    .B(n_3587),
    .Y(n_14181));
 AO21x1_ASAP7_75t_R g234884 (.A1(n_1022),
    .A2(n_790),
    .B(n_1036),
    .Y(n_14182));
 XNOR2xp5_ASAP7_75t_R g234885 (.A(u5_mul_69_18_n_2026),
    .B(u5_mul_69_18_n_1803),
    .Y(n_14183));
 AND2x2_ASAP7_75t_R g234886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .Y(n_14184));
 XNOR2xp5_ASAP7_75t_R g234887 (.A(u3_sub_52_45_Y_add_52_31_n_767),
    .B(u3_sub_52_45_Y_add_52_31_n_784),
    .Y(n_14185));
 XNOR2xp5_ASAP7_75t_R g234888 (.A(u5_mul_69_18_n_1978),
    .B(u5_mul_69_18_n_1881),
    .Y(n_14186));
 AND2x2_ASAP7_75t_R g234892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(n_14190));
 XNOR2xp5_ASAP7_75t_R g234893 (.A(u5_mul_69_18_n_1988),
    .B(u5_mul_69_18_n_1920),
    .Y(n_14191));
 AND2x2_ASAP7_75t_R g234894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .Y(n_14192));
 XNOR2xp5_ASAP7_75t_R g234895 (.A(u5_mul_69_18_n_2004),
    .B(u5_mul_69_18_n_1946),
    .Y(n_14193));
 XNOR2xp5_ASAP7_75t_R g234896 (.A(u5_mul_69_18_n_2024),
    .B(u5_mul_69_18_n_1831),
    .Y(n_14194));
 XNOR2xp5_ASAP7_75t_R g234898 (.A(u5_mul_69_18_n_1949),
    .B(u5_mul_69_18_n_1800),
    .Y(n_14196));
 OR2x2_ASAP7_75t_R g234899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1073),
    .Y(n_14197));
 AND2x2_ASAP7_75t_R g234901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .Y(n_14199));
 XNOR2xp5_ASAP7_75t_R g234902 (.A(u5_mul_69_18_n_2014),
    .B(u5_mul_69_18_n_1910),
    .Y(n_14200));
 XNOR2xp5_ASAP7_75t_R g234903 (.A(u5_mul_69_18_n_1974),
    .B(u5_mul_69_18_n_1858),
    .Y(n_14201));
 XNOR2xp5_ASAP7_75t_R g234905 (.A(u5_mul_69_18_n_2002),
    .B(u5_mul_69_18_n_1953),
    .Y(n_14203));
 AND2x2_ASAP7_75t_R g234906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_469),
    .Y(n_14204));
 XNOR2xp5_ASAP7_75t_R g234907 (.A(u5_mul_69_18_n_2036),
    .B(n_14374),
    .Y(n_14205));
 XNOR2xp5_ASAP7_75t_R g234911 (.A(u5_mul_69_18_n_2032),
    .B(u5_mul_69_18_n_1680),
    .Y(n_14209));
 XNOR2xp5_ASAP7_75t_R g234912 (.A(u5_mul_69_18_n_1641),
    .B(u5_mul_69_18_n_1511),
    .Y(n_14210));
 XNOR2xp5_ASAP7_75t_R g234914 (.A(u5_mul_69_18_n_2034),
    .B(u5_mul_69_18_n_1634),
    .Y(n_14212));
 OR2x2_ASAP7_75t_R g234916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2675),
    .Y(n_14214));
 XNOR2xp5_ASAP7_75t_R g234917 (.A(u5_mul_69_18_n_2028),
    .B(u5_mul_69_18_n_1758),
    .Y(n_14215));
 XNOR2xp5_ASAP7_75t_R g234920 (.A(u5_mul_69_18_n_1807),
    .B(u5_mul_69_18_n_1633),
    .Y(n_14218));
 AND2x2_ASAP7_75t_R g234921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .Y(n_14219));
 XNOR2xp5_ASAP7_75t_R g234922 (.A(u5_mul_69_18_n_2030),
    .B(u5_mul_69_18_n_1721),
    .Y(n_14220));
 XNOR2xp5_ASAP7_75t_R g234923 (.A(u5_mul_69_18_n_1893),
    .B(u5_mul_69_18_n_1722),
    .Y(n_14221));
 XNOR2xp5_ASAP7_75t_R g234924 (.A(u5_mul_69_18_n_1982),
    .B(u5_mul_69_18_n_1909),
    .Y(n_14222));
 AND2x2_ASAP7_75t_R g234926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .Y(n_14224));
 XNOR2xp5_ASAP7_75t_R g234927 (.A(u5_mul_69_18_n_2000),
    .B(u5_mul_69_18_n_1960),
    .Y(n_14225));
 XNOR2xp5_ASAP7_75t_R g234928 (.A(u5_mul_69_18_n_1976),
    .B(u5_mul_69_18_n_1882),
    .Y(n_14226));
 XNOR2xp5_ASAP7_75t_R g234930 (.A(u5_mul_69_18_n_1732),
    .B(u5_mul_69_18_n_1579),
    .Y(n_14228));
 XNOR2xp5_ASAP7_75t_R g234931 (.A(u5_mul_69_18_n_1996),
    .B(u5_mul_69_18_n_1966),
    .Y(n_14229));
 XNOR2xp5_ASAP7_75t_R g234932 (.A(u5_mul_69_18_n_1990),
    .B(u5_mul_69_18_n_1954),
    .Y(n_14230));
 XNOR2xp5_ASAP7_75t_R g234933 (.A(u5_mul_69_18_n_1970),
    .B(u5_mul_69_18_n_1829),
    .Y(n_14231));
 XNOR2xp5_ASAP7_75t_R g234935 (.A(u5_mul_69_18_n_1994),
    .B(u5_mul_69_18_n_1963),
    .Y(n_14233));
 XNOR2xp5_ASAP7_75t_R g234936 (.A(u5_mul_69_18_n_1965),
    .B(u5_mul_69_18_n_1802),
    .Y(n_14234));
 XNOR2xp5_ASAP7_75t_R g234937 (.A(u5_mul_69_18_n_1439),
    .B(u5_mul_69_18_n_1335),
    .Y(n_14235));
 XNOR2xp5_ASAP7_75t_R g234938 (.A(u5_mul_69_18_n_2008),
    .B(u5_mul_69_18_n_1955),
    .Y(n_14236));
 XNOR2xp5_ASAP7_75t_R g234939 (.A(u5_mul_69_18_n_2018),
    .B(u5_mul_69_18_n_1856),
    .Y(n_14237));
 XNOR2xp5_ASAP7_75t_R g234943 (.A(u5_mul_69_18_n_1986),
    .B(u5_mul_69_18_n_1923),
    .Y(n_14241));
 XNOR2xp5_ASAP7_75t_R g234945 (.A(u5_mul_69_18_n_1972),
    .B(u5_mul_69_18_n_1830),
    .Y(n_14243));
 XNOR2xp5_ASAP7_75t_R g234946 (.A(u5_mul_69_18_n_2016),
    .B(u5_mul_69_18_n_1883),
    .Y(n_14244));
 XNOR2xp5_ASAP7_75t_R g234947 (.A(u5_mul_69_18_n_2020),
    .B(u5_mul_69_18_n_1859),
    .Y(n_14245));
 XOR2xp5_ASAP7_75t_R g234948 (.A(u3_sub_52_45_Y_add_52_31_n_630),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(n_14246));
 XNOR2xp5_ASAP7_75t_R g234949 (.A(u5_mul_69_18_n_1864),
    .B(u5_mul_69_18_n_1678),
    .Y(n_14247));
 AND2x2_ASAP7_75t_R g234950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .Y(n_14248));
 XNOR2xp5_ASAP7_75t_R g234951 (.A(u5_mul_69_18_n_2022),
    .B(u5_mul_69_18_n_1828),
    .Y(n_14249));
 XNOR2xp5_ASAP7_75t_R g234952 (.A(u5_mul_69_18_n_2012),
    .B(u5_mul_69_18_n_1935),
    .Y(n_14250));
 XOR2xp5_ASAP7_75t_R g234953 (.A(u5_mul_69_18_n_1453),
    .B(u5_mul_69_18_n_1535),
    .Y(n_14251));
 XNOR2xp5_ASAP7_75t_R g234954 (.A(u5_mul_69_18_n_1998),
    .B(u5_mul_69_18_n_1959),
    .Y(n_14252));
 XNOR2xp5_ASAP7_75t_R g234956 (.A(u5_mul_69_18_n_1181),
    .B(u5_mul_69_18_n_1121),
    .Y(n_14254));
 XNOR2xp5_ASAP7_75t_R g234957 (.A(u5_mul_69_18_n_1992),
    .B(u5_mul_69_18_n_1952),
    .Y(n_14255));
 XNOR2xp5_ASAP7_75t_R g234958 (.A(u5_mul_69_18_n_2010),
    .B(u5_mul_69_18_n_1933),
    .Y(n_14256));
 XNOR2xp5_ASAP7_75t_R g234959 (.A(u5_mul_69_18_n_1968),
    .B(u5_mul_69_18_n_1801),
    .Y(n_14257));
 XNOR2xp5_ASAP7_75t_R g234960 (.A(u3_sub_52_45_Y_add_52_31_n_785),
    .B(u3_sub_52_45_Y_add_52_31_n_797),
    .Y(n_14258));
 XNOR2xp5_ASAP7_75t_R g234961 (.A(u3_sub_52_45_Y_add_52_31_n_699),
    .B(u3_sub_52_45_Y_add_52_31_n_762),
    .Y(n_14259));
 XNOR2xp5_ASAP7_75t_R g234963 (.A(u5_mul_69_18_n_2006),
    .B(u5_mul_69_18_n_1947),
    .Y(n_14261));
 XNOR2xp5_ASAP7_75t_R g234964 (.A(u5_mul_69_18_n_996),
    .B(u5_mul_69_18_n_891),
    .Y(n_14262));
 XNOR2xp5_ASAP7_75t_R g234965 (.A(u5_mul_69_18_n_1984),
    .B(u5_mul_69_18_n_1937),
    .Y(n_14263));
 AND2x2_ASAP7_75t_R g234966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(n_14264));
 AO21x1_ASAP7_75t_R g234968 (.A1(u5_mul_69_18_n_690),
    .A2(u5_mul_69_18_n_584),
    .B(u5_mul_69_18_n_891),
    .Y(n_14266));
 XNOR2xp5_ASAP7_75t_R g234969 (.A(u5_mul_69_18_n_1980),
    .B(u5_mul_69_18_n_1908),
    .Y(n_14267));
 AND2x2_ASAP7_75t_R g234970 (.A(u1_n_852),
    .B(n_1293),
    .Y(n_14268));
 AND2x2_ASAP7_75t_L g234971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_738),
    .Y(n_14269));
 AND3x1_ASAP7_75t_SL g234972 (.A(n_3198),
    .B(n_3213),
    .C(n_13837),
    .Y(n_14270));
 NAND2x1_ASAP7_75t_SL g234973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13674),
    .Y(n_14271));
 AND2x2_ASAP7_75t_R g234979 (.A(n_1186),
    .B(n_1177),
    .Y(n_14277));
 AND2x2_ASAP7_75t_R g234980 (.A(n_1184),
    .B(n_1183),
    .Y(n_14278));
 AND3x1_ASAP7_75t_R g234981 (.A(n_310),
    .B(n_1179),
    .C(n_1178),
    .Y(n_14279));
 XOR2x2_ASAP7_75t_L g234982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13355),
    .Y(n_14280));
 XOR2xp5_ASAP7_75t_L g234984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5932),
    .Y(n_14282));
 XNOR2xp5_ASAP7_75t_R g234985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5447),
    .Y(n_14283));
 XNOR2xp5_ASAP7_75t_R g234986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4932),
    .Y(n_14284));
 XOR2xp5_ASAP7_75t_R g234987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5103),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4942),
    .Y(n_14285));
 XNOR2xp5_ASAP7_75t_R g234988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4937),
    .Y(n_14286));
 XOR2xp5_ASAP7_75t_L g234989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4517),
    .Y(n_14287));
 XOR2xp5_ASAP7_75t_SL g234990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4487),
    .Y(n_14288));
 XOR2xp5_ASAP7_75t_R g234991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(n_14289));
 AO21x1_ASAP7_75t_SL g234992 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2851),
    .A2(n_3646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .Y(n_14290));
 XNOR2xp5_ASAP7_75t_L g234993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2772),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2670),
    .Y(n_14291));
 XNOR2xp5_ASAP7_75t_R g234994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3230),
    .B(n_14536),
    .Y(n_14292));
 NAND4xp75_ASAP7_75t_R g234995 (.A(n_2997),
    .B(n_2999),
    .C(n_14108),
    .D(n_3037),
    .Y(n_14293));
 NAND3xp33_ASAP7_75t_SL g234996 (.A(n_14114),
    .B(n_72),
    .C(n_3037),
    .Y(n_14294));
 FAx1_ASAP7_75t_R g234997 (.SN(n_14295),
    .A(n_1141),
    .B(n_1052),
    .CI(n_41),
    .CON(UNCONNECTED0));
 OAI221xp5_ASAP7_75t_R g234998 (.A1(n_13981),
    .A2(n_1228),
    .B1(u2_n_1831),
    .B2(n_134),
    .C(n_152),
    .Y(n_14296));
 NAND3xp33_ASAP7_75t_R g234999 (.A(n_14277),
    .B(n_1187),
    .C(n_1188),
    .Y(n_14297));
 FAx1_ASAP7_75t_R g235000 (.SN(n_14298),
    .A(u5_mul_69_18_n_1817),
    .B(u5_mul_69_18_n_1694),
    .CI(u5_mul_69_18_n_1788),
    .CON(UNCONNECTED1));
 FAx1_ASAP7_75t_R g235001 (.SN(n_14299),
    .A(u5_mul_69_18_n_1818),
    .B(n_14325),
    .CI(u5_mul_69_18_n_1821),
    .CON(UNCONNECTED2));
 FAx1_ASAP7_75t_R g235002 (.SN(n_14300),
    .A(u5_mul_69_18_n_1806),
    .B(n_14340),
    .CI(u5_mul_69_18_n_1790),
    .CON(UNCONNECTED3));
 FAx1_ASAP7_75t_R g235003 (.SN(n_14301),
    .A(u5_mul_69_18_n_1833),
    .B(u5_mul_69_18_n_1748),
    .CI(n_14341),
    .CON(UNCONNECTED4));
 FAx1_ASAP7_75t_R g235004 (.SN(n_14302),
    .A(n_14330),
    .B(n_14334),
    .CI(u5_mul_69_18_n_1749),
    .CON(UNCONNECTED5));
 FAx1_ASAP7_75t_R g235005 (.SN(n_14303),
    .A(n_14320),
    .B(u5_mul_69_18_n_1688),
    .CI(u5_mul_69_18_n_1789),
    .CON(UNCONNECTED6));
 FAx1_ASAP7_75t_R g235006 (.SN(n_14304),
    .A(n_14319),
    .B(u5_mul_69_18_n_1639),
    .CI(u5_mul_69_18_n_1750),
    .CON(UNCONNECTED7));
 FAx1_ASAP7_75t_R g235007 (.SN(n_14305),
    .A(u5_mul_69_18_n_1745),
    .B(n_14338),
    .CI(u5_mul_69_18_n_1783),
    .CON(UNCONNECTED8));
 FAx1_ASAP7_75t_R g235008 (.SN(n_14306),
    .A(n_14336),
    .B(n_14358),
    .CI(u5_mul_69_18_n_1707),
    .CON(UNCONNECTED9));
 FAx1_ASAP7_75t_R g235009 (.SN(n_14307),
    .A(u5_mul_69_18_n_1697),
    .B(u5_mul_69_18_n_1581),
    .CI(n_14335),
    .CON(UNCONNECTED10));
 FAx1_ASAP7_75t_R g235010 (.SN(n_14308),
    .A(u5_mul_69_18_n_1731),
    .B(u5_mul_69_18_n_1660),
    .CI(u5_mul_69_18_n_1692),
    .CON(UNCONNECTED11));
 FAx1_ASAP7_75t_R g235011 (.SN(n_14309),
    .A(u5_mul_69_18_n_1703),
    .B(n_14345),
    .CI(n_14329),
    .CON(UNCONNECTED12));
 FAx1_ASAP7_75t_R g235012 (.SN(n_14310),
    .A(u5_mul_69_18_n_1689),
    .B(u5_mul_69_18_n_1652),
    .CI(u5_mul_69_18_n_1696),
    .CON(UNCONNECTED13));
 FAx1_ASAP7_75t_R g235013 (.SN(n_14311),
    .A(u5_mul_69_18_n_1659),
    .B(n_14366),
    .CI(n_14337),
    .CON(UNCONNECTED14));
 FAx1_ASAP7_75t_R g235014 (.SN(n_14312),
    .A(u5_mul_69_18_n_1746),
    .B(u5_mul_69_18_n_1657),
    .CI(n_14365),
    .CON(UNCONNECTED15));
 FAx1_ASAP7_75t_R g235015 (.SN(n_14313),
    .A(n_14343),
    .B(n_14353),
    .CI(u5_mul_69_18_n_1658),
    .CON(UNCONNECTED16));
 FAx1_ASAP7_75t_R g235016 (.SN(n_14314),
    .A(u5_mul_69_18_n_1638),
    .B(u5_mul_69_18_n_1473),
    .CI(u5_mul_69_18_n_1618),
    .CON(UNCONNECTED17));
 FAx1_ASAP7_75t_R g235017 (.SN(n_14315),
    .A(u5_mul_69_18_n_1695),
    .B(u5_mul_69_18_n_1566),
    .CI(u5_mul_69_18_n_1554),
    .CON(UNCONNECTED18));
 FAx1_ASAP7_75t_R g235018 (.SN(n_14316),
    .A(n_14344),
    .B(n_14378),
    .CI(u5_mul_69_18_n_1621),
    .CON(UNCONNECTED19));
 FAx1_ASAP7_75t_R g235019 (.SN(n_14317),
    .A(u5_mul_69_18_n_1620),
    .B(u5_mul_69_18_n_1594),
    .CI(u5_mul_69_18_n_1654),
    .CON(UNCONNECTED20));
 FAx1_ASAP7_75t_R g235020 (.SN(n_14318),
    .A(u5_mul_69_18_n_1587),
    .B(u5_mul_69_18_n_1467),
    .CI(u5_mul_69_18_n_1619),
    .CON(UNCONNECTED21));
 FAx1_ASAP7_75t_R g235021 (.SN(n_14319),
    .A(n_14371),
    .B(u5_mul_69_18_n_1462),
    .CI(u5_mul_69_18_n_1568),
    .CON(UNCONNECTED22));
 FAx1_ASAP7_75t_R g235022 (.SN(n_14320),
    .A(n_14354),
    .B(u5_mul_69_18_n_1494),
    .CI(n_14350),
    .CON(UNCONNECTED23));
 FAx1_ASAP7_75t_R g235023 (.SN(n_14321),
    .A(n_14372),
    .B(u5_mul_69_18_n_1497),
    .CI(n_14369),
    .CON(UNCONNECTED24));
 FAx1_ASAP7_75t_R g235024 (.SN(n_14322),
    .A(n_14363),
    .B(n_14464),
    .CI(u5_mul_69_18_n_1463),
    .CON(UNCONNECTED25));
 FAx1_ASAP7_75t_R g235025 (.SN(n_14323),
    .A(u5_mul_69_18_n_1583),
    .B(u5_mul_69_18_n_1461),
    .CI(u5_mul_69_18_n_1564),
    .CON(UNCONNECTED26));
 FAx1_ASAP7_75t_R g235026 (.SN(n_14324),
    .A(n_14361),
    .B(u5_mul_69_18_n_1474),
    .CI(u5_mul_69_18_n_1598),
    .CON(UNCONNECTED27));
 FAx1_ASAP7_75t_R g235027 (.SN(n_14325),
    .A(u5_mul_69_18_n_1548),
    .B(n_14351),
    .CI(u5_mul_69_18_n_1565),
    .CON(UNCONNECTED28));
 FAx1_ASAP7_75t_R g235028 (.SN(n_14326),
    .A(n_14352),
    .B(u5_mul_69_18_n_1359),
    .CI(u5_mul_69_18_n_1563),
    .CON(UNCONNECTED29));
 FAx1_ASAP7_75t_R g235029 (.SN(n_14327),
    .A(u5_mul_69_18_n_1567),
    .B(n_14367),
    .CI(n_14346),
    .CON(UNCONNECTED30));
 FAx1_ASAP7_75t_R g235030 (.SN(n_14328),
    .A(u5_mul_69_18_n_1560),
    .B(u5_mul_69_18_n_1485),
    .CI(u5_mul_69_18_n_1684),
    .CON(UNCONNECTED31));
 FAx1_ASAP7_75t_R g235031 (.SN(n_14329),
    .A(u5_mul_69_18_n_1558),
    .B(n_14384),
    .CI(u5_mul_69_18_n_1491),
    .CON(UNCONNECTED32));
 FAx1_ASAP7_75t_R g235032 (.SN(n_14330),
    .A(u5_mul_69_18_n_1656),
    .B(n_14364),
    .CI(n_14370),
    .CON(UNCONNECTED33));
 FAx1_ASAP7_75t_R g235033 (.SN(n_14331),
    .A(u5_mul_69_18_n_1591),
    .B(u5_mul_69_18_n_1490),
    .CI(u5_mul_69_18_n_1470),
    .CON(UNCONNECTED34));
 FAx1_ASAP7_75t_R g235034 (.SN(n_14332),
    .A(n_14377),
    .B(u5_mul_69_18_n_1305),
    .CI(u5_mul_69_18_n_1534),
    .CON(UNCONNECTED35));
 FAx1_ASAP7_75t_R g235035 (.SN(n_14333),
    .A(n_14380),
    .B(u5_mul_69_18_n_1316),
    .CI(u5_mul_69_18_n_1499),
    .CON(UNCONNECTED36));
 FAx1_ASAP7_75t_R g235036 (.SN(n_14334),
    .A(u5_mul_69_18_n_1524),
    .B(u5_mul_69_18_n_1488),
    .CI(u5_mul_69_18_n_1464),
    .CON(UNCONNECTED37));
 FAx1_ASAP7_75t_R g235037 (.SN(n_14335),
    .A(n_14385),
    .B(u5_mul_69_18_n_1365),
    .CI(u5_mul_69_18_n_1475),
    .CON(UNCONNECTED38));
 FAx1_ASAP7_75t_R g235038 (.SN(n_14336),
    .A(u5_mul_69_18_n_1476),
    .B(n_14383),
    .CI(u5_mul_69_18_n_1466),
    .CON(UNCONNECTED39));
 FAx1_ASAP7_75t_R g235039 (.SN(n_14337),
    .A(u5_mul_69_18_n_1531),
    .B(u5_mul_69_18_n_1423),
    .CI(u5_mul_69_18_n_1465),
    .CON(UNCONNECTED40));
 FAx1_ASAP7_75t_R g235040 (.SN(n_14338),
    .A(u5_mul_69_18_n_1528),
    .B(n_14390),
    .CI(u5_mul_69_18_n_1484),
    .CON(UNCONNECTED41));
 FAx1_ASAP7_75t_R g235041 (.SN(n_14339),
    .A(u5_mul_69_18_n_1486),
    .B(u5_mul_69_18_n_1360),
    .CI(u5_mul_69_18_n_1546),
    .CON(UNCONNECTED42));
 FAx1_ASAP7_75t_R g235042 (.SN(n_14340),
    .A(u5_mul_69_18_n_1477),
    .B(n_14414),
    .CI(n_14373),
    .CON(UNCONNECTED43));
 FAx1_ASAP7_75t_R g235043 (.SN(n_14341),
    .A(u5_mul_69_18_n_1482),
    .B(n_14379),
    .CI(u5_mul_69_18_n_1551),
    .CON(UNCONNECTED44));
 FAx1_ASAP7_75t_R g235044 (.SN(n_14342),
    .A(u5_mul_69_18_n_1455),
    .B(u5_mul_69_18_n_1197),
    .CI(u5_mul_69_18_n_1418),
    .CON(UNCONNECTED45));
 FAx1_ASAP7_75t_R g235045 (.SN(n_14343),
    .A(u5_mul_69_18_n_1411),
    .B(u5_mul_69_18_n_1384),
    .CI(u5_mul_69_18_n_1498),
    .CON(UNCONNECTED46));
 FAx1_ASAP7_75t_R g235046 (.SN(n_14344),
    .A(u5_mul_69_18_n_1537),
    .B(u5_mul_69_18_n_1354),
    .CI(n_14408),
    .CON(UNCONNECTED47));
 FAx1_ASAP7_75t_R g235047 (.SN(n_14345),
    .A(u5_mul_69_18_n_1483),
    .B(u5_mul_69_18_n_1357),
    .CI(n_14442),
    .CON(UNCONNECTED48));
 FAx1_ASAP7_75t_R g235048 (.SN(n_14346),
    .A(n_14393),
    .B(u5_mul_69_18_n_1200),
    .CI(u5_mul_69_18_n_1421),
    .CON(UNCONNECTED49));
 FAx1_ASAP7_75t_R g235049 (.SN(n_14347),
    .A(u5_mul_69_18_n_1481),
    .B(n_14402),
    .CI(u5_mul_69_18_n_1188),
    .CON(UNCONNECTED50));
 FAx1_ASAP7_75t_R g235050 (.SN(n_14348),
    .A(u5_mul_69_18_n_1362),
    .B(n_14415),
    .CI(n_14381),
    .CON(UNCONNECTED51));
 FAx1_ASAP7_75t_R g235051 (.SN(n_14349),
    .A(n_14395),
    .B(n_14410),
    .CI(u5_mul_69_18_n_1419),
    .CON(UNCONNECTED52));
 FAx1_ASAP7_75t_R g235052 (.SN(n_14350),
    .A(u5_mul_69_18_n_1358),
    .B(n_14451),
    .CI(u5_mul_69_18_n_1417),
    .CON(UNCONNECTED53));
 FAx1_ASAP7_75t_R g235053 (.SN(n_14351),
    .A(u5_mul_69_18_n_1291),
    .B(u5_mul_69_18_n_1202),
    .CI(n_14425),
    .CON(UNCONNECTED54));
 FAx1_ASAP7_75t_R g235054 (.SN(n_14352),
    .A(u5_mul_69_18_n_1312),
    .B(u5_mul_69_18_n_1221),
    .CI(n_14421),
    .CON(UNCONNECTED55));
 FAx1_ASAP7_75t_R g235055 (.SN(n_14353),
    .A(u5_mul_69_18_n_1267),
    .B(u5_mul_69_18_n_1225),
    .CI(u5_mul_69_18_n_1310),
    .CON(UNCONNECTED56));
 FAx1_ASAP7_75t_R g235056 (.SN(n_14354),
    .A(n_14406),
    .B(u5_mul_69_18_n_1131),
    .CI(u5_mul_69_18_n_1213),
    .CON(UNCONNECTED57));
 FAx1_ASAP7_75t_R g235057 (.SN(n_14355),
    .A(n_14450),
    .B(u5_mul_69_18_n_1224),
    .CI(u5_mul_69_18_n_1327),
    .CON(UNCONNECTED58));
 FAx1_ASAP7_75t_R g235058 (.SN(n_14356),
    .A(n_14432),
    .B(u5_mul_69_18_n_1258),
    .CI(u5_mul_69_18_n_1205),
    .CON(UNCONNECTED59));
 FAx1_ASAP7_75t_R g235059 (.SN(n_14357),
    .A(n_14444),
    .B(u5_mul_69_18_n_1211),
    .CI(n_14429),
    .CON(UNCONNECTED60));
 FAx1_ASAP7_75t_R g235060 (.SN(n_14358),
    .A(u5_mul_69_18_n_1246),
    .B(u5_mul_69_18_n_1219),
    .CI(u5_mul_69_18_n_1331),
    .CON(UNCONNECTED61));
 FAx1_ASAP7_75t_R g235061 (.SN(n_14359),
    .A(u5_mul_69_18_n_1415),
    .B(u5_mul_69_18_n_1239),
    .CI(n_14407),
    .CON(UNCONNECTED62));
 FAx1_ASAP7_75t_R g235062 (.SN(n_14360),
    .A(n_14453),
    .B(n_14452),
    .CI(u5_mul_69_18_n_1364),
    .CON(UNCONNECTED63));
 FAx1_ASAP7_75t_R g235063 (.SN(n_14361),
    .A(u5_mul_69_18_n_1257),
    .B(u5_mul_69_18_n_1137),
    .CI(u5_mul_69_18_n_1203),
    .CON(UNCONNECTED64));
 FAx1_ASAP7_75t_R g235064 (.SN(n_14362),
    .A(u5_mul_69_18_n_1303),
    .B(u5_mul_69_18_n_845),
    .CI(u5_mul_69_18_n_1210),
    .CON(UNCONNECTED65));
 FAx1_ASAP7_75t_R g235065 (.SN(n_14363),
    .A(n_14399),
    .B(u5_mul_69_18_n_1241),
    .CI(u5_mul_69_18_n_1128),
    .CON(UNCONNECTED66));
 FAx1_ASAP7_75t_R g235066 (.SN(n_14364),
    .A(u5_mul_69_18_n_1260),
    .B(n_14456),
    .CI(u5_mul_69_18_n_1363),
    .CON(UNCONNECTED67));
 FAx1_ASAP7_75t_R g235067 (.SN(n_14365),
    .A(u5_mul_69_18_n_1232),
    .B(n_14420),
    .CI(n_14392),
    .CON(UNCONNECTED68));
 FAx1_ASAP7_75t_R g235068 (.SN(n_14366),
    .A(n_14446),
    .B(u5_mul_69_18_n_1339),
    .CI(u5_mul_69_18_n_1324),
    .CON(UNCONNECTED69));
 FAx1_ASAP7_75t_R g235069 (.SN(n_14367),
    .A(n_14448),
    .B(u5_mul_69_18_n_1171),
    .CI(n_14449),
    .CON(UNCONNECTED70));
 FAx1_ASAP7_75t_R g235070 (.SN(n_14368),
    .A(n_14447),
    .B(u5_mul_69_18_n_1130),
    .CI(u5_mul_69_18_n_1278),
    .CON(UNCONNECTED71));
 FAx1_ASAP7_75t_R g235071 (.SN(n_14369),
    .A(n_14436),
    .B(u5_mul_69_18_n_1144),
    .CI(u5_mul_69_18_n_1222),
    .CON(UNCONNECTED72));
 FAx1_ASAP7_75t_R g235072 (.SN(n_14370),
    .A(n_14437),
    .B(u5_mul_69_18_n_1147),
    .CI(u5_mul_69_18_n_1298),
    .CON(UNCONNECTED73));
 FAx1_ASAP7_75t_R g235073 (.SN(n_14371),
    .A(u5_mul_69_18_n_1306),
    .B(u5_mul_69_18_n_1164),
    .CI(n_14445),
    .CON(UNCONNECTED74));
 FAx1_ASAP7_75t_R g235074 (.SN(n_14372),
    .A(n_14439),
    .B(u5_mul_69_18_n_1148),
    .CI(n_14411),
    .CON(UNCONNECTED75));
 FAx1_ASAP7_75t_R g235075 (.SN(n_14373),
    .A(n_14400),
    .B(u5_mul_69_18_n_703),
    .CI(u5_mul_69_18_n_1126),
    .CON(UNCONNECTED76));
 FAx1_ASAP7_75t_R g235076 (.SN(n_14374),
    .A(u5_mul_69_18_n_1352),
    .B(u5_mul_69_18_n_1104),
    .CI(u5_mul_69_18_n_166),
    .CON(UNCONNECTED77));
 FAx1_ASAP7_75t_R g235077 (.SN(n_14375),
    .A(u5_mul_69_18_n_1158),
    .B(n_14460),
    .CI(u5_mul_69_18_n_1329),
    .CON(UNCONNECTED78));
 FAx1_ASAP7_75t_R g235078 (.SN(n_14376),
    .A(u5_mul_69_18_n_1229),
    .B(u5_mul_69_18_n_695),
    .CI(n_14413),
    .CON(UNCONNECTED79));
 FAx1_ASAP7_75t_R g235079 (.SN(n_14377),
    .A(u5_mul_69_18_n_1133),
    .B(u5_mul_69_18_n_1216),
    .CI(n_14416),
    .CON(UNCONNECTED80));
 FAx1_ASAP7_75t_R g235080 (.SN(n_14378),
    .A(u5_mul_69_18_n_1125),
    .B(u5_mul_69_18_n_1161),
    .CI(n_14433),
    .CON(UNCONNECTED81));
 FAx1_ASAP7_75t_R g235081 (.SN(n_14379),
    .A(u5_mul_69_18_n_1138),
    .B(u5_mul_69_18_n_1204),
    .CI(u5_mul_69_18_n_1132),
    .CON(UNCONNECTED82));
 FAx1_ASAP7_75t_R g235082 (.SN(n_14380),
    .A(u5_mul_69_18_n_1123),
    .B(u5_mul_69_18_n_699),
    .CI(u5_mul_69_18_n_1214),
    .CON(UNCONNECTED83));
 FAx1_ASAP7_75t_R g235083 (.SN(n_14381),
    .A(u5_mul_69_18_n_1215),
    .B(u5_mul_69_18_n_1000),
    .CI(n_14455),
    .CON(UNCONNECTED84));
 FAx1_ASAP7_75t_R g235084 (.SN(n_14382),
    .A(u5_mul_69_18_n_1206),
    .B(u5_mul_69_18_n_207),
    .CI(u5_mul_69_18_n_1266),
    .CON(UNCONNECTED85));
 FAx1_ASAP7_75t_R g235085 (.SN(n_14383),
    .A(u5_mul_69_18_n_1175),
    .B(u5_mul_69_18_n_173),
    .CI(u5_mul_69_18_n_1141),
    .CON(UNCONNECTED86));
 FAx1_ASAP7_75t_R g235086 (.SN(n_14384),
    .A(u5_mul_69_18_n_1163),
    .B(u5_mul_69_18_n_1116),
    .CI(u5_mul_69_18_n_1198),
    .CON(UNCONNECTED87));
 FAx1_ASAP7_75t_R g235087 (.SN(n_14385),
    .A(u5_mul_69_18_n_1191),
    .B(u5_mul_69_18_n_1159),
    .CI(u5_mul_69_18_n_1201),
    .CON(UNCONNECTED88));
 FAx1_ASAP7_75t_R g235088 (.SN(n_14386),
    .A(u5_mul_69_18_n_1189),
    .B(u5_mul_69_18_n_1217),
    .CI(n_14431),
    .CON(UNCONNECTED89));
 FAx1_ASAP7_75t_R g235089 (.SN(n_14387),
    .A(u5_mul_69_18_n_1145),
    .B(u5_mul_69_18_n_872),
    .CI(u5_mul_69_18_n_1167),
    .CON(UNCONNECTED90));
 FAx1_ASAP7_75t_R g235090 (.SN(n_14388),
    .A(u5_mul_69_18_n_1060),
    .B(u5_mul_69_18_n_992),
    .CI(n_14427),
    .CON(UNCONNECTED91));
 FAx1_ASAP7_75t_R g235091 (.SN(n_14389),
    .A(u5_mul_69_18_n_1119),
    .B(u5_mul_69_18_n_897),
    .CI(u5_mul_69_18_n_867),
    .CON(UNCONNECTED92));
 FAx1_ASAP7_75t_R g235092 (.SN(n_14390),
    .A(u5_mul_69_18_n_1117),
    .B(u5_mul_69_18_n_851),
    .CI(u5_mul_69_18_n_1146),
    .CON(UNCONNECTED93));
 FAx1_ASAP7_75t_R g235093 (.SN(n_14391),
    .A(n_14457),
    .B(u5_mul_69_18_n_855),
    .CI(u5_mul_69_18_n_905),
    .CON(UNCONNECTED94));
 FAx1_ASAP7_75t_R g235094 (.SN(n_14392),
    .A(u5_mul_69_18_n_1155),
    .B(u5_mul_69_18_n_998),
    .CI(u5_mul_69_18_n_773),
    .CON(UNCONNECTED95));
 FAx1_ASAP7_75t_R g235095 (.SN(n_14393),
    .A(u5_mul_69_18_n_994),
    .B(u5_mul_69_18_n_731),
    .CI(u5_mul_69_18_n_1062),
    .CON(UNCONNECTED96));
 FAx1_ASAP7_75t_R g235096 (.SN(n_14394),
    .A(u5_mul_69_18_n_1002),
    .B(u5_mul_69_18_n_784),
    .CI(u5_mul_69_18_n_1220),
    .CON(UNCONNECTED97));
 FAx1_ASAP7_75t_R g235097 (.SN(n_14395),
    .A(u5_mul_69_18_n_1154),
    .B(u5_mul_69_18_n_1001),
    .CI(u5_mul_69_18_n_874),
    .CON(UNCONNECTED98));
 FAx1_ASAP7_75t_R g235098 (.SN(n_14396),
    .A(u5_mul_69_18_n_1176),
    .B(u5_mul_69_18_n_706),
    .CI(u5_mul_69_18_n_210),
    .CON(UNCONNECTED99));
 FAx1_ASAP7_75t_R g235099 (.SN(n_14397),
    .A(u5_mul_69_18_n_952),
    .B(u5_mul_69_18_n_653),
    .CI(u5_mul_69_18_n_660),
    .CON(UNCONNECTED100));
 FAx1_ASAP7_75t_R g235100 (.SN(n_14398),
    .A(u5_mul_69_18_n_785),
    .B(u5_mul_69_18_n_961),
    .CI(u5_mul_69_18_n_993),
    .CON(UNCONNECTED101));
 FAx1_ASAP7_75t_R g235101 (.SN(n_14399),
    .A(u5_mul_69_18_n_930),
    .B(u5_mul_69_18_n_775),
    .CI(u5_mul_69_18_n_707),
    .CON(UNCONNECTED102));
 FAx1_ASAP7_75t_R g235102 (.SN(n_14400),
    .A(u5_mul_69_18_n_896),
    .B(u5_mul_69_18_n_768),
    .CI(u5_mul_69_18_n_807),
    .CON(UNCONNECTED103));
 FAx1_ASAP7_75t_R g235103 (.SN(n_14401),
    .A(u5_mul_69_18_n_900),
    .B(u5_mul_69_18_n_841),
    .CI(u5_mul_69_18_n_170),
    .CON(UNCONNECTED104));
 FAx1_ASAP7_75t_R g235104 (.SN(n_14402),
    .A(u5_mul_69_18_n_848),
    .B(u5_mul_69_18_n_893),
    .CI(u5_mul_69_18_n_967),
    .CON(UNCONNECTED105));
 FAx1_ASAP7_75t_R g235105 (.SN(n_14403),
    .A(u5_mul_69_18_n_880),
    .B(u5_mul_69_18_n_899),
    .CI(u5_mul_69_18_n_980),
    .CON(UNCONNECTED106));
 FAx1_ASAP7_75t_R g235106 (.SN(n_14404),
    .A(u5_mul_69_18_n_906),
    .B(u5_mul_69_18_n_748),
    .CI(u5_mul_69_18_n_1003),
    .CON(UNCONNECTED107));
 FAx1_ASAP7_75t_R g235107 (.SN(n_14405),
    .A(u5_mul_69_18_n_696),
    .B(u5_mul_69_18_n_977),
    .CI(u5_mul_69_18_n_189),
    .CON(UNCONNECTED108));
 FAx1_ASAP7_75t_R g235108 (.SN(n_14406),
    .A(u5_mul_69_18_n_787),
    .B(u5_mul_69_18_n_869),
    .CI(u5_mul_69_18_n_973),
    .CON(UNCONNECTED109));
 FAx1_ASAP7_75t_R g235109 (.SN(n_14407),
    .A(u5_mul_69_18_n_718),
    .B(u5_mul_69_18_n_797),
    .CI(u5_mul_69_18_n_928),
    .CON(UNCONNECTED110));
 FAx1_ASAP7_75t_R g235110 (.SN(n_14408),
    .A(u5_mul_69_18_n_970),
    .B(u5_mul_69_18_n_212),
    .CI(u5_mul_69_18_n_695),
    .CON(UNCONNECTED111));
 FAx1_ASAP7_75t_R g235111 (.SN(n_14409),
    .A(u5_mul_69_18_n_802),
    .B(u5_mul_69_18_n_709),
    .CI(u5_mul_69_18_n_631),
    .CON(UNCONNECTED112));
 FAx1_ASAP7_75t_R g235112 (.SN(n_14410),
    .A(u5_mul_69_18_n_910),
    .B(u5_mul_69_18_n_674),
    .CI(u5_mul_69_18_n_810),
    .CON(UNCONNECTED113));
 FAx1_ASAP7_75t_R g235113 (.SN(n_14411),
    .A(u5_mul_69_18_n_925),
    .B(u5_mul_69_18_n_879),
    .CI(u5_mul_69_18_n_946),
    .CON(UNCONNECTED114));
 FAx1_ASAP7_75t_R g235114 (.SN(n_14412),
    .A(u5_mul_69_18_n_908),
    .B(u5_mul_69_18_n_758),
    .CI(u5_mul_69_18_n_805),
    .CON(UNCONNECTED115));
 FAx1_ASAP7_75t_R g235115 (.SN(n_14413),
    .A(u5_mul_69_18_n_876),
    .B(u5_mul_69_18_n_923),
    .CI(u5_mul_69_18_n_840),
    .CON(UNCONNECTED116));
 FAx1_ASAP7_75t_R g235116 (.SN(n_14414),
    .A(u5_mul_69_18_n_723),
    .B(u5_mul_69_18_n_969),
    .CI(u5_mul_69_18_n_209),
    .CON(UNCONNECTED117));
 FAx1_ASAP7_75t_R g235117 (.SN(n_14415),
    .A(u5_mul_69_18_n_889),
    .B(u5_mul_69_18_n_661),
    .CI(u5_mul_69_18_n_957),
    .CON(UNCONNECTED118));
 FAx1_ASAP7_75t_R g235118 (.SN(n_14416),
    .A(u5_mul_69_18_n_737),
    .B(u5_mul_69_18_n_790),
    .CI(u5_mul_69_18_n_665),
    .CON(UNCONNECTED119));
 FAx1_ASAP7_75t_R g235119 (.SN(n_14417),
    .A(u5_mul_69_18_n_864),
    .B(u5_mul_69_18_n_656),
    .CI(u5_mul_69_18_n_937),
    .CON(UNCONNECTED120));
 FAx1_ASAP7_75t_R g235120 (.SN(n_14418),
    .A(u5_mul_69_18_n_752),
    .B(u5_mul_69_18_n_668),
    .CI(u5_mul_69_18_n_836),
    .CON(UNCONNECTED121));
 FAx1_ASAP7_75t_R g235121 (.SN(n_14419),
    .A(u5_mul_69_18_n_762),
    .B(u5_mul_69_18_n_664),
    .CI(u5_mul_69_18_n_806),
    .CON(UNCONNECTED122));
 FAx1_ASAP7_75t_R g235122 (.SN(n_14420),
    .A(u5_mul_69_18_n_782),
    .B(u5_mul_69_18_n_657),
    .CI(u5_mul_69_18_n_792),
    .CON(UNCONNECTED123));
 FAx1_ASAP7_75t_R g235123 (.SN(n_14421),
    .A(u5_mul_69_18_n_971),
    .B(u5_mul_69_18_n_187),
    .CI(u5_mul_69_18_n_706),
    .CON(UNCONNECTED124));
 FAx1_ASAP7_75t_R g235124 (.SN(n_14422),
    .A(u5_mul_69_18_n_711),
    .B(u5_mul_69_18_n_663),
    .CI(u5_mul_69_18_n_830),
    .CON(UNCONNECTED125));
 FAx1_ASAP7_75t_R g235125 (.SN(n_14423),
    .A(u5_mul_69_18_n_966),
    .B(u5_mul_69_18_n_205),
    .CI(u5_mul_69_18_n_845),
    .CON(UNCONNECTED126));
 FAx1_ASAP7_75t_R g235126 (.SN(n_14424),
    .A(u5_mul_69_18_n_920),
    .B(u5_mul_69_18_n_732),
    .CI(u5_mul_69_18_n_825),
    .CON(UNCONNECTED127));
 FAx1_ASAP7_75t_R g235127 (.SN(n_14425),
    .A(u5_mul_69_18_n_742),
    .B(u5_mul_69_18_n_789),
    .CI(u5_mul_69_18_n_834),
    .CON(UNCONNECTED128));
 FAx1_ASAP7_75t_R g235128 (.SN(n_14426),
    .A(u5_mul_69_18_n_749),
    .B(u5_mul_69_18_n_751),
    .CI(u5_mul_69_18_n_816),
    .CON(UNCONNECTED129));
 FAx1_ASAP7_75t_R g235129 (.SN(n_14427),
    .A(u5_mul_69_18_n_909),
    .B(u5_mul_69_18_n_858),
    .CI(u5_mul_69_18_n_954),
    .CON(UNCONNECTED130));
 FAx1_ASAP7_75t_R g235130 (.SN(n_14428),
    .A(u5_mul_69_18_n_796),
    .B(u5_mul_69_18_n_645),
    .CI(u5_mul_69_18_n_753),
    .CON(UNCONNECTED131));
 FAx1_ASAP7_75t_R g235131 (.SN(n_14429),
    .A(u5_mul_69_18_n_714),
    .B(u5_mul_69_18_n_650),
    .CI(u5_mul_69_18_n_794),
    .CON(UNCONNECTED132));
 FAx1_ASAP7_75t_R g235132 (.SN(n_14430),
    .A(u5_mul_69_18_n_919),
    .B(u5_mul_69_18_n_652),
    .CI(u5_mul_69_18_n_831),
    .CON(UNCONNECTED133));
 FAx1_ASAP7_75t_R g235133 (.SN(n_14431),
    .A(u5_mul_69_18_n_733),
    .B(u5_mul_69_18_n_735),
    .CI(u5_mul_69_18_n_944),
    .CON(UNCONNECTED134));
 FAx1_ASAP7_75t_R g235134 (.SN(n_14432),
    .A(u5_mul_69_18_n_839),
    .B(u5_mul_69_18_n_921),
    .CI(u5_mul_69_18_n_882),
    .CON(UNCONNECTED135));
 FAx1_ASAP7_75t_R g235135 (.SN(n_14433),
    .A(u5_mul_69_18_n_780),
    .B(u5_mul_69_18_n_757),
    .CI(u5_mul_69_18_n_963),
    .CON(UNCONNECTED136));
 FAx1_ASAP7_75t_R g235136 (.SN(n_14434),
    .A(u5_mul_69_18_n_866),
    .B(u5_mul_69_18_n_870),
    .CI(u5_mul_69_18_n_955),
    .CON(UNCONNECTED137));
 FAx1_ASAP7_75t_R g235137 (.SN(n_14435),
    .A(u5_mul_69_18_n_877),
    .B(u5_mul_69_18_n_885),
    .CI(u5_mul_69_18_n_817),
    .CON(UNCONNECTED138));
 FAx1_ASAP7_75t_R g235138 (.SN(n_14436),
    .A(u5_mul_69_18_n_857),
    .B(u5_mul_69_18_n_856),
    .CI(u5_mul_69_18_n_932),
    .CON(UNCONNECTED139));
 FAx1_ASAP7_75t_R g235139 (.SN(n_14437),
    .A(u5_mul_69_18_n_888),
    .B(u5_mul_69_18_n_729),
    .CI(u5_mul_69_18_n_809),
    .CON(UNCONNECTED140));
 FAx1_ASAP7_75t_R g235140 (.SN(n_14438),
    .A(u5_mul_69_18_n_776),
    .B(u5_mul_69_18_n_712),
    .CI(u5_mul_69_18_n_838),
    .CON(UNCONNECTED141));
 FAx1_ASAP7_75t_R g235141 (.SN(n_14439),
    .A(u5_mul_69_18_n_852),
    .B(u5_mul_69_18_n_854),
    .CI(u5_mul_69_18_n_953),
    .CON(UNCONNECTED142));
 FAx1_ASAP7_75t_R g235142 (.SN(n_14440),
    .A(u5_mul_69_18_n_739),
    .B(u5_mul_69_18_n_821),
    .CI(u5_mul_69_18_n_734),
    .CON(UNCONNECTED143));
 FAx1_ASAP7_75t_R g235143 (.SN(n_14441),
    .A(u5_mul_69_18_n_788),
    .B(u5_mul_69_18_n_743),
    .CI(u5_mul_69_18_n_791),
    .CON(UNCONNECTED144));
 FAx1_ASAP7_75t_R g235144 (.SN(n_14442),
    .A(u5_mul_69_18_n_798),
    .B(u5_mul_69_18_n_778),
    .CI(u5_mul_69_18_n_850),
    .CON(UNCONNECTED145));
 FAx1_ASAP7_75t_R g235145 (.SN(n_14443),
    .A(u5_mul_69_18_n_902),
    .B(u5_mul_69_18_n_746),
    .CI(u5_mul_69_18_n_814),
    .CON(UNCONNECTED146));
 FAx1_ASAP7_75t_R g235146 (.SN(n_14444),
    .A(u5_mul_69_18_n_781),
    .B(u5_mul_69_18_n_892),
    .CI(u5_mul_69_18_n_799),
    .CON(UNCONNECTED147));
 FAx1_ASAP7_75t_R g235147 (.SN(n_14445),
    .A(u5_mul_69_18_n_837),
    .B(u5_mul_69_18_n_853),
    .CI(u5_mul_69_18_n_849),
    .CON(UNCONNECTED148));
 FAx1_ASAP7_75t_R g235148 (.SN(n_14446),
    .A(u5_mul_69_18_n_771),
    .B(u5_mul_69_18_n_769),
    .CI(u5_mul_69_18_n_803),
    .CON(UNCONNECTED149));
 FAx1_ASAP7_75t_R g235149 (.SN(n_14447),
    .A(u5_mul_69_18_n_756),
    .B(u5_mul_69_18_n_726),
    .CI(u5_mul_69_18_n_818),
    .CON(UNCONNECTED150));
 FAx1_ASAP7_75t_R g235150 (.SN(n_14448),
    .A(u5_mul_69_18_n_736),
    .B(u5_mul_69_18_n_904),
    .CI(u5_mul_69_18_n_822),
    .CON(UNCONNECTED151));
 FAx1_ASAP7_75t_R g235151 (.SN(n_14449),
    .A(u5_mul_69_18_n_741),
    .B(u5_mul_69_18_n_926),
    .CI(u5_mul_69_18_n_819),
    .CON(UNCONNECTED152));
 FAx1_ASAP7_75t_R g235152 (.SN(n_14450),
    .A(u5_mul_69_18_n_965),
    .B(u5_mul_69_18_n_755),
    .CI(u5_mul_69_18_n_914),
    .CON(UNCONNECTED153));
 FAx1_ASAP7_75t_R g235153 (.SN(n_14451),
    .A(u5_mul_69_18_n_750),
    .B(u5_mul_69_18_n_903),
    .CI(u5_mul_69_18_n_960),
    .CON(UNCONNECTED154));
 FAx1_ASAP7_75t_R g235154 (.SN(n_14452),
    .A(u5_mul_69_18_n_721),
    .B(u5_mul_69_18_n_722),
    .CI(u5_mul_69_18_n_959),
    .CON(UNCONNECTED155));
 FAx1_ASAP7_75t_R g235155 (.SN(n_14453),
    .A(u5_mul_69_18_n_720),
    .B(u5_mul_69_18_n_12),
    .CI(u5_mul_69_18_n_941),
    .CON(UNCONNECTED156));
 FAx1_ASAP7_75t_R g235156 (.SN(n_14454),
    .A(u5_mul_69_18_n_865),
    .B(u5_mul_69_18_n_777),
    .CI(u5_mul_69_18_n_949),
    .CON(UNCONNECTED157));
 FAx1_ASAP7_75t_R g235157 (.SN(n_14455),
    .A(u5_mul_69_18_n_958),
    .B(u5_mul_69_18_n_648),
    .CI(u5_mul_69_18_n_924),
    .CON(UNCONNECTED158));
 FAx1_ASAP7_75t_R g235158 (.SN(n_14456),
    .A(u5_mul_69_18_n_943),
    .B(u5_mul_69_18_n_646),
    .CI(u5_mul_69_18_n_765),
    .CON(UNCONNECTED159));
 FAx1_ASAP7_75t_R g235159 (.SN(n_14457),
    .A(u5_mul_69_18_n_677),
    .B(u5_mul_69_18_n_651),
    .CI(u5_mul_69_18_n_800),
    .CON(UNCONNECTED160));
 FAx1_ASAP7_75t_R g235160 (.SN(n_14458),
    .A(u5_mul_69_18_n_659),
    .B(u5_mul_69_18_n_649),
    .CI(u5_mul_69_18_n_936),
    .CON(UNCONNECTED161));
 FAx1_ASAP7_75t_R g235161 (.SN(n_14459),
    .A(u5_mul_69_18_n_662),
    .B(u5_mul_69_18_n_654),
    .CI(u5_mul_69_18_n_811),
    .CON(UNCONNECTED162));
 FAx1_ASAP7_75t_R g235162 (.SN(n_14460),
    .A(u5_mul_69_18_n_675),
    .B(u5_mul_69_18_n_647),
    .CI(u5_mul_69_18_n_935),
    .CON(UNCONNECTED163));
 FAx1_ASAP7_75t_R g235163 (.SN(n_14461),
    .A(u5_mul_69_18_n_1705),
    .B(u5_mul_69_18_n_1616),
    .CI(n_14328),
    .CON(UNCONNECTED164));
 FAx1_ASAP7_75t_R g235164 (.SN(n_14462),
    .A(u5_mul_69_18_n_1700),
    .B(n_14347),
    .CI(u5_mul_69_18_n_1614),
    .CON(UNCONNECTED165));
 FAx1_ASAP7_75t_R g235165 (.SN(n_14463),
    .A(u5_mul_69_18_n_1487),
    .B(u5_mul_69_18_n_1361),
    .CI(u5_mul_69_18_n_1326),
    .CON(UNCONNECTED166));
 FAx1_ASAP7_75t_R g235166 (.SN(n_14464),
    .A(u5_mul_69_18_n_1420),
    .B(u5_mul_69_18_n_1236),
    .CI(u5_mul_69_18_n_1196),
    .CON(UNCONNECTED167));
 O2A1O1Ixp33_ASAP7_75t_L g235167 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2339),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13118),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .Y(n_14465));
 A2O1A1Ixp33_ASAP7_75t_L g235168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12301),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12553),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .Y(n_14466));
 INVxp33_ASAP7_75t_R g235169 (.A(n_14467),
    .Y(n_14468));
 A2O1A1Ixp33_ASAP7_75t_R g235170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10999),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11077),
    .Y(n_14467));
 FAx1_ASAP7_75t_R g235171 (.SN(n_14469),
    .A(u6_rem_96_22_Y_u6_div_90_17_n_10337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .CI(u6_rem_96_22_Y_u6_div_90_17_n_10375),
    .CON(UNCONNECTED168));
 INVxp33_ASAP7_75t_R g235173 (.A(n_14471),
    .Y(n_14472));
 A2O1A1Ixp33_ASAP7_75t_R g235174 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1949),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9921),
    .Y(n_14471));
 OA211x2_ASAP7_75t_R g235175 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1930),
    .Y(n_14473));
 AOI31xp33_ASAP7_75t_SL g235176 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1835),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9044),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_8904),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1846),
    .Y(n_14474));
 INVxp67_ASAP7_75t_R g235177 (.A(n_14475),
    .Y(n_14476));
 A2O1A1Ixp33_ASAP7_75t_L g235178 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8127),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8332),
    .Y(n_14475));
 OA211x2_ASAP7_75t_R g235179 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1730),
    .Y(n_14477));
 O2A1O1Ixp33_ASAP7_75t_L g235180 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7904),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .Y(n_14478));
 A2O1A1Ixp33_ASAP7_75t_R g235181 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7121),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7318),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .Y(n_14479));
 AOI211xp5_ASAP7_75t_SL g235182 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1607),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7196),
    .Y(n_14480));
 AO21x1_ASAP7_75t_R g235183 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7019),
    .Y(n_14481));
 AOI31xp33_ASAP7_75t_SL g235184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1560),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1532),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_6478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1557),
    .Y(n_14482));
 INVxp33_ASAP7_75t_R g235185 (.A(n_14483),
    .Y(n_14484));
 A2O1A1Ixp33_ASAP7_75t_R g235186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5834),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5948),
    .Y(n_14483));
 A2O1A1Ixp33_ASAP7_75t_L g235187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4959),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5080),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(n_14485));
 A2O1A1Ixp33_ASAP7_75t_R g235188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5014),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5133),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(n_14486));
 A2O1A1Ixp33_ASAP7_75t_L g235189 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4500),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4648),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4691),
    .Y(n_14487));
 OA21x2_ASAP7_75t_L g235190 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4297),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4358),
    .Y(n_14488));
 AO221x1_ASAP7_75t_L g235191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3644),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2761),
    .Y(n_14489));
 AO221x1_ASAP7_75t_R g235192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3644),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2586),
    .Y(n_14490));
 AOI32xp33_ASAP7_75t_SL g235193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .A2(n_3647),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_788),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_712),
    .B2(n_14290),
    .Y(n_14491));
 AOI21xp33_ASAP7_75t_SL g235194 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_708),
    .Y(n_14492));
 A2O1A1Ixp33_ASAP7_75t_SL g235195 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2101),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11186),
    .C(n_14024),
    .Y(n_14493));
 FAx1_ASAP7_75t_R g235196 (.SN(n_14494),
    .A(u3_sub_52_45_Y_add_52_31_n_702),
    .B(u3_sub_52_45_Y_add_52_31_n_792),
    .CI(fracta[3]),
    .CON(UNCONNECTED169));
 FAx1_ASAP7_75t_R g235197 (.SN(n_14495),
    .A(u3_sub_52_45_Y_add_52_31_n_639),
    .B(u3_sub_52_45_Y_add_52_31_n_786),
    .CI(fracta[24]),
    .CON(UNCONNECTED170));
 FAx1_ASAP7_75t_R g235198 (.SN(n_14496),
    .A(u3_sub_52_45_Y_add_52_31_n_693),
    .B(u3_sub_52_45_Y_add_52_31_n_796),
    .CI(fracta[6]),
    .CON(UNCONNECTED171));
 FAx1_ASAP7_75t_R g235199 (.SN(n_14497),
    .A(u3_sub_52_45_Y_add_52_31_n_681),
    .B(u3_sub_52_45_Y_add_52_31_n_777),
    .CI(fracta[10]),
    .CON(UNCONNECTED172));
 FAx1_ASAP7_75t_L g235200 (.SN(n_14498),
    .A(u3_sub_52_45_Y_add_52_31_n_672),
    .B(u3_sub_52_45_Y_add_52_31_n_778),
    .CI(fracta[13]),
    .CON(UNCONNECTED173));
 FAx1_ASAP7_75t_R g235201 (.SN(n_14499),
    .A(u3_sub_52_45_Y_add_52_31_n_675),
    .B(u3_sub_52_45_Y_add_52_31_n_772),
    .CI(fracta[12]),
    .CON(UNCONNECTED174));
 FAx1_ASAP7_75t_L g235202 (.SN(n_14500),
    .A(u3_sub_52_45_Y_add_52_31_n_690),
    .B(u3_sub_52_45_Y_add_52_31_n_780),
    .CI(fracta[7]),
    .CON(UNCONNECTED175));
 FAx1_ASAP7_75t_R g235203 (.SN(n_14501),
    .A(u3_sub_52_45_Y_add_52_31_n_642),
    .B(u3_sub_52_45_Y_add_52_31_n_773),
    .CI(fracta[23]),
    .CON(UNCONNECTED176));
 FAx1_ASAP7_75t_R g235204 (.SN(n_14502),
    .A(u3_sub_52_45_Y_add_52_31_n_645),
    .B(u3_sub_52_45_Y_add_52_31_n_793),
    .CI(fracta[22]),
    .CON(UNCONNECTED177));
 FAx1_ASAP7_75t_R g235205 (.SN(n_14503),
    .A(u3_sub_52_45_Y_add_52_31_n_651),
    .B(u3_sub_52_45_Y_add_52_31_n_782),
    .CI(fracta[20]),
    .CON(UNCONNECTED178));
 FAx1_ASAP7_75t_R g235206 (.SN(n_14504),
    .A(u3_sub_52_45_Y_add_52_31_n_666),
    .B(u3_sub_52_45_Y_add_52_31_n_791),
    .CI(fracta[15]),
    .CON(UNCONNECTED179));
 FAx1_ASAP7_75t_R g235207 (.SN(n_14505),
    .A(u3_sub_52_45_Y_add_52_31_n_663),
    .B(u3_sub_52_45_Y_add_52_31_n_794),
    .CI(fracta[16]),
    .CON(UNCONNECTED180));
 FAx1_ASAP7_75t_R g235208 (.SN(n_14506),
    .A(u3_sub_52_45_Y_add_52_31_n_657),
    .B(u3_sub_52_45_Y_add_52_31_n_770),
    .CI(fracta[18]),
    .CON(UNCONNECTED181));
 FAx1_ASAP7_75t_R g235209 (.SN(n_14507),
    .A(u3_sub_52_45_Y_add_52_31_n_654),
    .B(u3_sub_52_45_Y_add_52_31_n_775),
    .CI(fracta[19]),
    .CON(UNCONNECTED182));
 FAx1_ASAP7_75t_R g235210 (.SN(n_14508),
    .A(u3_sub_52_45_Y_add_52_31_n_669),
    .B(u3_sub_52_45_Y_add_52_31_n_795),
    .CI(fracta[14]),
    .CON(UNCONNECTED183));
 FAx1_ASAP7_75t_R g235211 (.SN(n_14509),
    .A(u3_sub_52_45_Y_add_52_31_n_633),
    .B(u3_sub_52_45_Y_add_52_31_n_790),
    .CI(fracta[26]),
    .CON(UNCONNECTED184));
 FAx1_ASAP7_75t_R g235212 (.SN(n_14510),
    .A(u3_sub_52_45_Y_add_52_31_n_684),
    .B(u3_sub_52_45_Y_add_52_31_n_779),
    .CI(fracta[9]),
    .CON(UNCONNECTED185));
 FAx1_ASAP7_75t_R g235213 (.SN(n_14511),
    .A(u3_sub_52_45_Y_add_52_31_n_687),
    .B(u3_sub_52_45_Y_add_52_31_n_776),
    .CI(fracta[8]),
    .CON(UNCONNECTED186));
 FAx1_ASAP7_75t_R g235214 (.SN(n_14512),
    .A(u3_sub_52_45_Y_add_52_31_n_648),
    .B(u3_sub_52_45_Y_add_52_31_n_789),
    .CI(fracta[21]),
    .CON(UNCONNECTED187));
 FAx1_ASAP7_75t_R g235215 (.SN(n_14513),
    .A(u3_sub_52_45_Y_add_52_31_n_636),
    .B(u3_sub_52_45_Y_add_52_31_n_771),
    .CI(fracta[25]),
    .CON(UNCONNECTED188));
 FAx1_ASAP7_75t_R g235216 (.SN(n_14514),
    .A(u3_sub_52_45_Y_add_52_31_n_660),
    .B(u3_sub_52_45_Y_add_52_31_n_774),
    .CI(fracta[17]),
    .CON(UNCONNECTED189));
 FAx1_ASAP7_75t_R g235217 (.SN(n_14515),
    .A(u3_sub_52_45_Y_add_52_31_n_678),
    .B(u3_sub_52_45_Y_add_52_31_n_781),
    .CI(fracta[11]),
    .CON(UNCONNECTED190));
 FAx1_ASAP7_75t_R g235218 (.SN(n_14516),
    .A(u3_sub_52_45_Y_add_52_31_n_696),
    .B(u3_sub_52_45_Y_add_52_31_n_787),
    .CI(fracta[5]),
    .CON(UNCONNECTED191));
 OAI21xp33_ASAP7_75t_R g235219 (.A1(n_1401),
    .A2(n_1402),
    .B(n_14517),
    .Y(n_14518));
 MAJx2_ASAP7_75t_R g235220 (.A(n_1349),
    .B(n_1387),
    .C(u1_n_1045),
    .Y(n_14517));
 NAND2xp5_ASAP7_75t_L g235221 (.A(n_14519),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(n_14520));
 XOR2xp5_ASAP7_75t_R g235222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8211),
    .Y(n_14519));
 AO21x1_ASAP7_75t_L g235223 (.A1(n_14521),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7000),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7178),
    .Y(n_14522));
 NOR2xp33_ASAP7_75t_L g235224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1636),
    .Y(n_14521));
 OAI21xp33_ASAP7_75t_R g235225 (.A1(n_14523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(n_14524));
 AO21x1_ASAP7_75t_R g235226 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1586),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .Y(n_14523));
 NAND2xp33_ASAP7_75t_R g235227 (.A(n_14525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(n_14526));
 XOR2xp5_ASAP7_75t_R g235228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1458),
    .Y(n_14525));
 NOR2xp33_ASAP7_75t_SL g235229 (.A(n_14527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(n_14528));
 XNOR2xp5_ASAP7_75t_R g235230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5102),
    .Y(n_14527));
 OAI21xp33_ASAP7_75t_SL g235231 (.A1(n_14529),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4050),
    .Y(n_14530));
 MAJIxp5_ASAP7_75t_SL g235232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1029),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4013),
    .Y(n_14529));
 OA21x2_ASAP7_75t_SL g235233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3934),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3928),
    .B(n_14531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3969));
 AOI21xp5_ASAP7_75t_L g235234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3957),
    .Y(n_14531));
 NAND2xp33_ASAP7_75t_L g235235 (.A(n_14533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(n_14534));
 XOR2xp5_ASAP7_75t_L g235236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3535),
    .Y(n_14533));
 HAxp5_ASAP7_75t_R g235237 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2507),
    .CON(n_14536),
    .SN(n_14535));
 NOR2xp33_ASAP7_75t_R g235239 (.A(opa_r1[2]),
    .B(sub_327_16_n_589),
    .Y(n_14564));
 A2O1A1Ixp33_ASAP7_75t_L g235241 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7632),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7812),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(n_14575));
 INVxp33_ASAP7_75t_R g235246 (.A(u5_mul_69_18_n_673),
    .Y(u5_mul_69_18_n_843));
 INVxp33_ASAP7_75t_R g27155 (.A(u4_n_1439),
    .Y(n_3490));
 INVxp33_ASAP7_75t_R g27156 (.A(u4_n_1091),
    .Y(n_3489));
 INVxp33_ASAP7_75t_R g27157 (.A(n_3813),
    .Y(n_3488));
 INVxp33_ASAP7_75t_R g27158 (.A(n_3571),
    .Y(n_3487));
 INVxp33_ASAP7_75t_R g27160 (.A(u4_n_1438),
    .Y(n_3491));
 INVxp33_ASAP7_75t_R g27162 (.A(u1_n_980),
    .Y(n_3481));
 INVxp33_ASAP7_75t_R g27164 (.A(n_3759),
    .Y(n_3480));
 INVxp33_ASAP7_75t_R g27166 (.A(n_3824),
    .Y(n_3483));
 INVxp67_ASAP7_75t_R g27168 (.A(fasu_op),
    .Y(u3_sub_52_45_Y_add_52_31_n_841));
 INVxp33_ASAP7_75t_R g27198 (.A(fpu_op[0]),
    .Y(n_3287));
 HB1xp67_ASAP7_75t_R g27210 (.A(n_3297),
    .Y(n_3444));
 HB1xp67_ASAP7_75t_R g27212 (.A(n_14120),
    .Y(n_3297));
 HB1xp67_ASAP7_75t_R g27218 (.A(n_3353),
    .Y(n_3476));
 HB1xp67_ASAP7_75t_R g27220 (.A(n_14114),
    .Y(n_3353));
 HB1xp67_ASAP7_75t_R g27222 (.A(n_3350),
    .Y(n_3438));
 HB1xp67_ASAP7_75t_R g27224 (.A(n_14106),
    .Y(n_3350));
 HB1xp67_ASAP7_75t_R g27226 (.A(n_3355),
    .Y(n_3436));
 HB1xp67_ASAP7_75t_R g27228 (.A(n_14090),
    .Y(n_3355));
 HB1xp67_ASAP7_75t_R g27230 (.A(n_3344),
    .Y(n_3434));
 HB1xp67_ASAP7_75t_R g27232 (.A(n_14102),
    .Y(n_3344));
 INVxp33_ASAP7_75t_R g27233 (.A(u5_mul_69_18_n_106),
    .Y(n_3432));
 HB1xp67_ASAP7_75t_R g27237 (.A(n_14108),
    .Y(n_3337));
 HB1xp67_ASAP7_75t_R g27243 (.A(n_3294),
    .Y(n_3427));
 HB1xp67_ASAP7_75t_R g27245 (.A(n_14092),
    .Y(n_3294));
 HB1xp67_ASAP7_75t_R g27271 (.A(n_3311),
    .Y(n_3415));
 HB1xp67_ASAP7_75t_R g27273 (.A(n_14116),
    .Y(n_3311));
 HB1xp67_ASAP7_75t_R g27279 (.A(n_3306),
    .Y(n_3411));
 HB1xp67_ASAP7_75t_R g27281 (.A(n_14094),
    .Y(n_3306));
 HB1xp67_ASAP7_75t_R g27283 (.A(n_3305),
    .Y(n_3409));
 HB1xp67_ASAP7_75t_R g27285 (.A(n_14100),
    .Y(n_3305));
 HB1xp67_ASAP7_75t_R g27289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .Y(n_3303));
 HB1xp67_ASAP7_75t_R g27332 (.A(n_3310),
    .Y(n_3401));
 HB1xp67_ASAP7_75t_R g27334 (.A(n_14174),
    .Y(n_3310));
 HB1xp67_ASAP7_75t_R g27342 (.A(n_14088),
    .Y(n_3302));
 HB1xp67_ASAP7_75t_R g27344 (.A(n_3299),
    .Y(n_3395));
 HB1xp67_ASAP7_75t_R g27346 (.A(n_14098),
    .Y(n_3299));
 HB1xp67_ASAP7_75t_R g27357 (.A(n_3292),
    .Y(n_3386));
 HB1xp67_ASAP7_75t_R g27359 (.A(n_14176),
    .Y(n_3292));
 HB1xp67_ASAP7_75t_R g27362 (.A(n_2896),
    .Y(n_3336));
 HB1xp67_ASAP7_75t_R g27365 (.A(n_3345),
    .Y(n_3440));
 HB1xp67_ASAP7_75t_R g27367 (.A(n_14096),
    .Y(n_3345));
 HB1xp67_ASAP7_75t_R g27369 (.A(n_3349),
    .Y(n_3474));
 HB1xp67_ASAP7_75t_R g27371 (.A(n_14118),
    .Y(n_3349));
 HB1xp67_ASAP7_75t_R g27373 (.A(n_3351),
    .Y(n_3472));
 HB1xp67_ASAP7_75t_R g27375 (.A(n_14172),
    .Y(n_3351));
 HB1xp67_ASAP7_75t_R g27381 (.A(n_3358),
    .Y(n_3468));
 HB1xp67_ASAP7_75t_R g27383 (.A(n_14110),
    .Y(n_3358));
 HB1xp67_ASAP7_75t_R g27385 (.A(n_3341),
    .Y(n_3466));
 HB1xp67_ASAP7_75t_R g27387 (.A(n_14112),
    .Y(n_3341));
 HB1xp67_ASAP7_75t_R g27409 (.A(n_3347),
    .Y(n_3456));
 HB1xp67_ASAP7_75t_R g27411 (.A(n_14170),
    .Y(n_3347));
 HB1xp67_ASAP7_75t_R g27413 (.A(n_3354),
    .Y(n_3452));
 HB1xp67_ASAP7_75t_R g27415 (.A(n_14168),
    .Y(n_3354));
 HB1xp67_ASAP7_75t_R g27421 (.A(n_3348),
    .Y(n_3454));
 HB1xp67_ASAP7_75t_R g27423 (.A(n_14166),
    .Y(n_3348));
 AO21x1_ASAP7_75t_R g27424__2398 (.A1(n_3802),
    .A2(n_3222),
    .B(n_3760),
    .Y(u4_exp_zero));
 NAND3xp33_ASAP7_75t_R g27425__5107 (.A(n_3800),
    .B(rmode_r3[1]),
    .C(u4_n_1792),
    .Y(n_3222));
 NAND2xp33_ASAP7_75t_R g27426__6260 (.A(u4_n_1792),
    .B(n_3800),
    .Y(n_3579));
 INVxp33_ASAP7_75t_R g27427 (.A(n_3221),
    .Y(n_3800));
 AOI31xp33_ASAP7_75t_R g27428__4319 (.A1(n_3220),
    .A2(n_3596),
    .A3(u4_n_1446),
    .B(n_3577),
    .Y(n_3221));
 NAND2xp33_ASAP7_75t_R g27429__8428 (.A(u4_exp_out[7]),
    .B(u4_round2a_BAR),
    .Y(n_3220));
 NAND3xp33_ASAP7_75t_R g27430__5526 (.A(n_15699_BAR),
    .B(n_3219),
    .C(n_3578),
    .Y(u4_exp_out[7]));
 NAND2xp33_ASAP7_75t_R g27431__6783 (.A(n_3597),
    .B(n_3750),
    .Y(n_3219));
 AOI221xp5_ASAP7_75t_R g27571 (.A1(n_621),
    .A2(opa_r1[28]),
    .B1(n_620),
    .B2(exp_mul[5]),
    .C(n_628),
    .Y(n_639));
 AOI221xp5_ASAP7_75t_R g27572 (.A1(n_621),
    .A2(opa_r1[27]),
    .B1(n_620),
    .B2(exp_mul[4]),
    .C(n_631),
    .Y(n_638));
 AOI221xp5_ASAP7_75t_R g27573 (.A1(n_621),
    .A2(opa_r1[26]),
    .B1(n_620),
    .B2(exp_mul[3]),
    .C(n_630),
    .Y(n_637));
 AOI221xp5_ASAP7_75t_R g27574 (.A1(n_621),
    .A2(opa_r1[29]),
    .B1(n_620),
    .B2(exp_mul[6]),
    .C(n_625),
    .Y(n_636));
 AOI221xp5_ASAP7_75t_R g27575 (.A1(n_621),
    .A2(opa_r1[23]),
    .B1(n_620),
    .B2(exp_mul[0]),
    .C(n_629),
    .Y(n_635));
 AOI221xp5_ASAP7_75t_R g27576 (.A1(n_621),
    .A2(opa_r1[30]),
    .B1(n_620),
    .B2(exp_mul[7]),
    .C(n_626),
    .Y(n_634));
 AOI221xp5_ASAP7_75t_R g27577 (.A1(n_621),
    .A2(opa_r1[24]),
    .B1(n_620),
    .B2(exp_mul[1]),
    .C(n_627),
    .Y(n_633));
 AOI221xp5_ASAP7_75t_R g27578 (.A1(n_621),
    .A2(opa_r1[25]),
    .B1(n_620),
    .B2(exp_mul[2]),
    .C(n_624),
    .Y(n_632));
 AO22x1_ASAP7_75t_R g27579 (.A1(exp_fasu[4]),
    .A2(n_622),
    .B1(exp_r[4]),
    .B2(n_623),
    .Y(n_631));
 AO22x1_ASAP7_75t_R g27580 (.A1(exp_fasu[3]),
    .A2(n_622),
    .B1(exp_r[3]),
    .B2(n_623),
    .Y(n_630));
 AO22x1_ASAP7_75t_R g27581 (.A1(exp_fasu[0]),
    .A2(n_622),
    .B1(exp_r[0]),
    .B2(n_623),
    .Y(n_629));
 AO22x1_ASAP7_75t_R g27582 (.A1(exp_fasu[5]),
    .A2(n_622),
    .B1(exp_r[5]),
    .B2(n_623),
    .Y(n_628));
 AO22x1_ASAP7_75t_R g27583 (.A1(exp_fasu[1]),
    .A2(n_622),
    .B1(exp_r[1]),
    .B2(n_623),
    .Y(n_627));
 AO22x1_ASAP7_75t_R g27584 (.A1(exp_fasu[7]),
    .A2(n_622),
    .B1(exp_r[7]),
    .B2(n_623),
    .Y(n_626));
 AO22x1_ASAP7_75t_R g27585 (.A1(exp_fasu[6]),
    .A2(n_622),
    .B1(exp_r[6]),
    .B2(n_623),
    .Y(n_625));
 AO22x1_ASAP7_75t_R g27586 (.A1(exp_fasu[2]),
    .A2(n_622),
    .B1(exp_r[2]),
    .B2(n_623),
    .Y(n_624));
 AND2x2_ASAP7_75t_R g27587 (.A(fpu_op_r2[1]),
    .B(n_3557),
    .Y(n_623));
 NOR2xp33_ASAP7_75t_R g27588 (.A(fpu_op_r2[2]),
    .B(fpu_op_r2[1]),
    .Y(n_622));
 INVxp33_ASAP7_75t_R g27589 (.A(n_3499),
    .Y(n_621));
 INVxp33_ASAP7_75t_R g27590 (.A(n_3557),
    .Y(n_620));
 XOR2xp5_ASAP7_75t_R g3 (.A(exp_r[3]),
    .B(n_3716),
    .Y(n_13841));
 OR2x2_ASAP7_75t_SL g35524__3680 (.A(n_3212),
    .B(n_3218),
    .Y(n_3646));
 A2O1A1Ixp33_ASAP7_75t_SL g35525__1617 (.A1(n_3203),
    .A2(n_3177),
    .B(n_2942),
    .C(n_3180),
    .Y(n_3839));
 A2O1A1Ixp33_ASAP7_75t_SL g35526__2802 (.A1(n_3208),
    .A2(n_3181),
    .B(n_2942),
    .C(n_3176),
    .Y(n_3838));
 OAI22xp33_ASAP7_75t_R g35527__1705 (.A1(n_2942),
    .A2(n_3214),
    .B1(n_2941),
    .B2(n_83),
    .Y(n_3643));
 A2O1A1Ixp33_ASAP7_75t_R g35528__5122 (.A1(n_3186),
    .A2(n_3167),
    .B(n_2942),
    .C(n_3201),
    .Y(n_3642));
 NAND3xp33_ASAP7_75t_SL g35529__8246 (.A(n_3196),
    .B(n_13835),
    .C(n_13834),
    .Y(n_3645));
 OAI221xp5_ASAP7_75t_R g35531__6131 (.A1(n_3210),
    .A2(n_2942),
    .B1(n_3541),
    .B2(n_3084),
    .C(n_3141),
    .Y(n_3641));
 OAI221xp5_ASAP7_75t_R g35532__1881 (.A1(n_3543),
    .A2(n_3084),
    .B1(n_72),
    .B2(n_2941),
    .C(n_3216),
    .Y(n_3640));
 OAI22xp33_ASAP7_75t_R g35533__5115 (.A1(fracta_mul[23]),
    .A2(n_3207),
    .B1(n_3049),
    .B2(n_73),
    .Y(n_3639));
 OAI311xp33_ASAP7_75t_SL g35534__7482 (.A1(n_3847),
    .A2(n_88),
    .A3(n_2944),
    .B1(n_3217),
    .C1(n_3189),
    .Y(n_3218));
 OAI221xp5_ASAP7_75t_R g35535__4733 (.A1(n_14294),
    .A2(n_3084),
    .B1(n_84),
    .B2(n_3049),
    .C(n_3215),
    .Y(n_3636));
 OAI22xp33_ASAP7_75t_R g35536__6161 (.A1(fracta_mul[23]),
    .A2(n_3206),
    .B1(n_3049),
    .B2(n_90),
    .Y(n_3633));
 AOI21xp5_ASAP7_75t_SL g35537__9315 (.A1(n_3182),
    .A2(n_2940),
    .B(n_3202),
    .Y(n_3217));
 OAI31xp33_ASAP7_75t_R g35538__9945 (.A1(n_3166),
    .A2(n_3135),
    .A3(n_3152),
    .B(n_2941),
    .Y(n_3216));
 A2O1A1Ixp33_ASAP7_75t_R g35539__2883 (.A1(n_14096),
    .A2(n_2936),
    .B(n_3190),
    .C(n_3049),
    .Y(n_3215));
 OAI221xp5_ASAP7_75t_R g35540__2346 (.A1(n_3188),
    .A2(n_13883),
    .B1(n_3045),
    .B2(n_3091),
    .C(n_3140),
    .Y(n_3637));
 NOR4xp25_ASAP7_75t_R g35541__1666 (.A(n_3204),
    .B(n_3168),
    .C(n_3156),
    .D(n_3115),
    .Y(n_3214));
 AO21x1_ASAP7_75t_R g35542__7410 (.A1(n_13883),
    .A2(n_14112),
    .B(n_3209),
    .Y(n_3638));
 OAI22xp33_ASAP7_75t_R g35543__6417 (.A1(n_13884),
    .A2(n_3184),
    .B1(n_3049),
    .B2(n_80),
    .Y(n_3634));
 OAI22xp33_ASAP7_75t_R g35544__5477 (.A1(n_13884),
    .A2(n_3193),
    .B1(n_3049),
    .B2(n_79),
    .Y(n_3635));
 NOR3xp33_ASAP7_75t_L g35545__2398 (.A(n_3199),
    .B(n_3160),
    .C(n_3158),
    .Y(n_3213));
 NAND3xp33_ASAP7_75t_SL g35546__5107 (.A(n_13836),
    .B(n_3178),
    .C(n_3185),
    .Y(n_3212));
 AND4x1_ASAP7_75t_R g35548__4319 (.A(n_3155),
    .B(n_3092),
    .C(n_3132),
    .D(n_3150),
    .Y(n_3210));
 AOI31xp33_ASAP7_75t_R g35549__8428 (.A1(n_3171),
    .A2(n_3093),
    .A3(n_3117),
    .B(n_13883),
    .Y(n_3209));
 OAI221xp5_ASAP7_75t_R g35550__5526 (.A1(n_3840),
    .A2(n_3084),
    .B1(n_3020),
    .B2(n_3089),
    .C(n_3174),
    .Y(n_3630));
 AOI211xp5_ASAP7_75t_R g35551__6783 (.A1(n_2951),
    .A2(n_14092),
    .B(n_3192),
    .C(n_3097),
    .Y(n_3208));
 AND4x1_ASAP7_75t_R g35552__3680 (.A(n_3162),
    .B(n_3126),
    .C(n_3112),
    .D(n_3094),
    .Y(n_3207));
 AOI221xp5_ASAP7_75t_R g35553__1617 (.A1(n_2934),
    .A2(n_14092),
    .B1(n_2930),
    .B2(n_14096),
    .C(n_3179),
    .Y(n_3206));
 OAI221xp5_ASAP7_75t_R g35555__1705 (.A1(n_3849),
    .A2(n_88),
    .B1(n_3541),
    .B2(n_78),
    .C(n_3145),
    .Y(n_3204));
 NOR2xp33_ASAP7_75t_L g35556__5122 (.A(n_3187),
    .B(n_3169),
    .Y(n_3203));
 A2O1A1O1Ixp25_ASAP7_75t_SL g35557__8246 (.A1(n_14293),
    .A2(n_3077),
    .B(n_79),
    .C(n_3149),
    .D(n_13838),
    .Y(n_3202));
 OAI221xp5_ASAP7_75t_R g35558__7098 (.A1(n_3125),
    .A2(n_13883),
    .B1(n_3034),
    .B2(n_3084),
    .C(n_3139),
    .Y(n_3631));
 A2O1A1Ixp33_ASAP7_75t_R g35559__6131 (.A1(n_3060),
    .A2(n_3120),
    .B(fracta_mul[23]),
    .C(n_3082),
    .Y(n_3632));
 AOI221xp5_ASAP7_75t_R g35560__1881 (.A1(n_2951),
    .A2(n_3083),
    .B1(n_2953),
    .B2(n_3088),
    .C(n_3142),
    .Y(n_3201));
 OAI21xp5_ASAP7_75t_SL g35561__5115 (.A1(n_2944),
    .A2(n_3165),
    .B(n_3194),
    .Y(n_3200));
 OAI21xp33_ASAP7_75t_SL g35562__7482 (.A1(n_2944),
    .A2(n_3164),
    .B(n_3191),
    .Y(n_3199));
 AOI31xp33_ASAP7_75t_L g35563__4733 (.A1(n_2953),
    .A2(n_14098),
    .A3(n_2940),
    .B(n_3183),
    .Y(n_3198));
 AOI21xp5_ASAP7_75t_SL g35565__9315 (.A1(n_3173),
    .A2(n_2940),
    .B(n_3175),
    .Y(n_3196));
 OAI21xp33_ASAP7_75t_L g35567__2883 (.A1(n_3058),
    .A2(n_3133),
    .B(n_2940),
    .Y(n_3194));
 AOI211xp5_ASAP7_75t_R g35568__2346 (.A1(n_2947),
    .A2(n_14090),
    .B(n_3127),
    .C(n_3161),
    .Y(n_3193));
 NAND3xp33_ASAP7_75t_R g35569__1666 (.A(n_3110),
    .B(n_3114),
    .C(n_3069),
    .Y(n_3192));
 OAI21xp33_ASAP7_75t_L g35570__7410 (.A1(n_3065),
    .A2(n_3113),
    .B(n_2940),
    .Y(n_3191));
 NAND3xp33_ASAP7_75t_R g35571__6417 (.A(n_3105),
    .B(n_3121),
    .C(n_3064),
    .Y(n_3190));
 A2O1A1Ixp33_ASAP7_75t_SL g35572__5477 (.A1(n_14096),
    .A2(n_3071),
    .B(n_3109),
    .C(n_2940),
    .Y(n_3189));
 AOI221xp5_ASAP7_75t_R g35573__2398 (.A1(n_2947),
    .A2(n_2907),
    .B1(n_2946),
    .B2(n_14096),
    .C(n_3170),
    .Y(n_3188));
 NAND3xp33_ASAP7_75t_R g35574__5107 (.A(n_3111),
    .B(n_3106),
    .C(n_3130),
    .Y(n_3187));
 AOI221xp5_ASAP7_75t_R g35575__6260 (.A1(n_3047),
    .A2(n_2907),
    .B1(n_2938),
    .B2(n_14102),
    .C(n_3159),
    .Y(n_3186));
 NAND4xp25_ASAP7_75t_R g35576__4319 (.A(n_2952),
    .B(n_14090),
    .C(n_14092),
    .D(n_2940),
    .Y(n_3185));
 AOI21xp33_ASAP7_75t_R g35577__8428 (.A1(n_2947),
    .A2(n_14088),
    .B(n_3172),
    .Y(n_3184));
 A2O1A1Ixp33_ASAP7_75t_L g35578__5526 (.A1(n_3079),
    .A2(n_3068),
    .B(n_2944),
    .C(n_3080),
    .Y(n_3183));
 OAI21xp33_ASAP7_75t_SL g35579__6783 (.A1(n_82),
    .A2(n_3849),
    .B(n_3157),
    .Y(n_3182));
 OAI221xp5_ASAP7_75t_R g35580__3680 (.A1(n_2928),
    .A2(n_3089),
    .B1(n_3091),
    .B2(n_76),
    .C(n_3138),
    .Y(n_3629));
 AOI21xp33_ASAP7_75t_R g35581__1617 (.A1(n_2907),
    .A2(n_2953),
    .B(n_3153),
    .Y(n_3181));
 NOR2xp33_ASAP7_75t_R g35582__2802 (.A(n_3148),
    .B(n_3147),
    .Y(n_3180));
 OAI211xp5_ASAP7_75t_R g35583__1705 (.A1(n_91),
    .A2(n_2935),
    .B(n_3099),
    .C(n_3026),
    .Y(n_3179));
 NAND3xp33_ASAP7_75t_R g35584__5122 (.A(n_14102),
    .B(n_2940),
    .C(n_2953),
    .Y(n_3178));
 AOI21xp33_ASAP7_75t_R g35585__8246 (.A1(n_2953),
    .A2(n_14096),
    .B(n_3143),
    .Y(n_3177));
 OAI222xp33_ASAP7_75t_R g35586__7098 (.A1(n_2928),
    .A2(n_3084),
    .B1(n_3089),
    .B2(n_76),
    .C1(n_78),
    .C2(n_3049),
    .Y(n_3628));
 AOI221xp5_ASAP7_75t_R g35587__6131 (.A1(n_3071),
    .A2(n_3083),
    .B1(n_3087),
    .B2(n_3088),
    .C(n_3081),
    .Y(n_3176));
 OAI31xp33_ASAP7_75t_L g35588__1881 (.A1(n_3849),
    .A2(n_74),
    .A3(n_2944),
    .B(n_3078),
    .Y(n_3175));
 AOI322xp5_ASAP7_75t_R g35589__5115 (.A1(n_2882),
    .A2(n_2907),
    .A3(n_3049),
    .B1(n_3090),
    .B2(n_2877),
    .C1(n_14096),
    .C2(n_13884),
    .Y(n_3174));
 NAND3xp33_ASAP7_75t_R g35590__7482 (.A(n_2952),
    .B(n_3014),
    .C(n_2940),
    .Y(n_3647));
 NOR3xp33_ASAP7_75t_R g35591__4733 (.A(n_3848),
    .B(n_88),
    .C(n_78),
    .Y(n_3173));
 OAI211xp5_ASAP7_75t_R g35592__6161 (.A1(n_91),
    .A2(n_2945),
    .B(n_3118),
    .C(n_3063),
    .Y(n_3172));
 AOI221xp5_ASAP7_75t_R g35593__9315 (.A1(n_2938),
    .A2(n_2907),
    .B1(n_2947),
    .B2(n_14096),
    .C(n_3129),
    .Y(n_3171));
 OAI211xp5_ASAP7_75t_R g35594__9945 (.A1(n_90),
    .A2(n_2932),
    .B(n_3116),
    .C(n_3040),
    .Y(n_3170));
 OAI221xp5_ASAP7_75t_R g35595__2883 (.A1(n_3055),
    .A2(n_90),
    .B1(n_3053),
    .B2(n_80),
    .C(n_3124),
    .Y(n_3169));
 OAI221xp5_ASAP7_75t_R g35596__2346 (.A1(n_3055),
    .A2(n_82),
    .B1(n_3053),
    .B2(n_2887),
    .C(n_3123),
    .Y(n_3168));
 AOI221xp5_ASAP7_75t_R g35597__1666 (.A1(n_2949),
    .A2(n_14096),
    .B1(n_2948),
    .B2(n_14098),
    .C(n_3122),
    .Y(n_3167));
 OAI221xp5_ASAP7_75t_R g35598__7410 (.A1(n_3055),
    .A2(n_78),
    .B1(n_3053),
    .B2(n_2908),
    .C(n_3119),
    .Y(n_3166));
 NOR2xp33_ASAP7_75t_SL g35599__6417 (.A(n_3101),
    .B(n_3104),
    .Y(n_3165));
 NOR2xp33_ASAP7_75t_L g35600__5477 (.A(n_3098),
    .B(n_3102),
    .Y(n_3164));
 OAI21xp33_ASAP7_75t_L g35601__2398 (.A1(n_2908),
    .A2(n_3070),
    .B(n_3107),
    .Y(n_3163));
 AOI221xp5_ASAP7_75t_R g35602__5107 (.A1(n_2948),
    .A2(n_14092),
    .B1(n_2939),
    .B2(n_2907),
    .C(n_3128),
    .Y(n_3162));
 OAI221xp5_ASAP7_75t_R g35603__6260 (.A1(n_3034),
    .A2(n_74),
    .B1(n_3020),
    .B2(n_2887),
    .C(n_3103),
    .Y(n_3161));
 NOR3xp33_ASAP7_75t_R g35604__4319 (.A(n_3070),
    .B(n_78),
    .C(n_2944),
    .Y(n_3160));
 OAI211xp5_ASAP7_75t_R g35605__8428 (.A1(n_80),
    .A2(n_3052),
    .B(n_3100),
    .C(n_3062),
    .Y(n_3159));
 NOR3xp33_ASAP7_75t_R g35606__5526 (.A(n_3849),
    .B(n_2908),
    .C(n_2944),
    .Y(n_3158));
 AOI221xp5_ASAP7_75t_R g35607__6783 (.A1(n_2947),
    .A2(n_14116),
    .B1(n_2946),
    .B2(n_14166),
    .C(n_3067),
    .Y(n_3157));
 OAI21xp33_ASAP7_75t_R g35608__3680 (.A1(n_74),
    .A2(n_14293),
    .B(n_3108),
    .Y(n_3156));
 AOI222xp33_ASAP7_75t_R g35609__1617 (.A1(n_3047),
    .A2(n_14092),
    .B1(n_2946),
    .B2(n_2896),
    .C1(n_2930),
    .C2(n_14112),
    .Y(n_3155));
 OAI22xp33_ASAP7_75t_R g35610__2802 (.A1(n_88),
    .A2(n_3845),
    .B1(n_91),
    .B2(n_3844),
    .Y(n_3154));
 OAI21xp33_ASAP7_75t_R g35611__1705 (.A1(n_74),
    .A2(n_3543),
    .B(n_3096),
    .Y(n_3153));
 OAI221xp5_ASAP7_75t_R g35612__5122 (.A1(n_82),
    .A2(n_3045),
    .B1(n_2887),
    .B2(n_3052),
    .C(n_3059),
    .Y(n_3152));
 OAI21xp33_ASAP7_75t_SL g35613__8246 (.A1(n_78),
    .A2(n_3845),
    .B(n_3095),
    .Y(n_3151));
 AOI221xp5_ASAP7_75t_R g35614__7098 (.A1(n_2938),
    .A2(n_2888),
    .B1(n_2947),
    .B2(n_14102),
    .C(n_3061),
    .Y(n_3150));
 AOI221xp5_ASAP7_75t_L g35615__6131 (.A1(n_2934),
    .A2(n_14170),
    .B1(n_3035),
    .B2(n_14168),
    .C(n_2944),
    .Y(n_3149));
 OAI22xp33_ASAP7_75t_R g35616__1881 (.A1(n_3084),
    .A2(n_3844),
    .B1(n_2941),
    .B2(n_85),
    .Y(n_3148));
 OAI22xp33_ASAP7_75t_R g35617__5115 (.A1(n_3089),
    .A2(n_3070),
    .B1(n_3091),
    .B2(n_3849),
    .Y(n_3147));
 OAI22xp5_ASAP7_75t_R g35618__7482 (.A1(n_82),
    .A2(n_2950),
    .B1(n_90),
    .B2(n_3543),
    .Y(n_3146));
 AOI22xp33_ASAP7_75t_R g35619__4733 (.A1(n_14090),
    .A2(n_2951),
    .B1(n_2907),
    .B2(n_3086),
    .Y(n_3145));
 OAI22xp33_ASAP7_75t_R g35620__6161 (.A1(n_74),
    .A2(n_2950),
    .B1(n_2887),
    .B2(n_3543),
    .Y(n_3144));
 OAI22xp33_ASAP7_75t_R g35621__9315 (.A1(n_2908),
    .A2(n_2950),
    .B1(n_82),
    .B2(n_3543),
    .Y(n_3143));
 OAI22xp33_ASAP7_75t_R g35622__9945 (.A1(n_3091),
    .A2(n_3543),
    .B1(n_2941),
    .B2(n_95),
    .Y(n_3142));
 AOI22xp33_ASAP7_75t_R g35623__2883 (.A1(n_3088),
    .A2(n_3086),
    .B1(n_2942),
    .B2(n_14166),
    .Y(n_3141));
 OAI22xp33_ASAP7_75t_R g35624__2346 (.A1(n_76),
    .A2(n_3084),
    .B1(n_3049),
    .B2(n_91),
    .Y(n_3627));
 AOI22xp33_ASAP7_75t_R g35625__1666 (.A1(n_3083),
    .A2(n_2948),
    .B1(n_13883),
    .B2(n_14110),
    .Y(n_3140));
 AOI22xp33_ASAP7_75t_R g35626__7410 (.A1(n_3090),
    .A2(n_2930),
    .B1(fracta_mul[23]),
    .B2(n_14098),
    .Y(n_3139));
 AOI22xp33_ASAP7_75t_R g35627__6417 (.A1(n_3083),
    .A2(n_2930),
    .B1(n_13883),
    .B2(n_2907),
    .Y(n_3138));
 OAI22xp33_ASAP7_75t_R g35628__5477 (.A1(n_91),
    .A2(n_3845),
    .B1(n_78),
    .B2(n_3844),
    .Y(n_3137));
 OAI22xp5_ASAP7_75t_L g35629__2398 (.A1(n_2908),
    .A2(n_3844),
    .B1(n_2887),
    .B2(n_2950),
    .Y(n_3136));
 OAI222xp33_ASAP7_75t_R g35630__5107 (.A1(n_2945),
    .A2(n_90),
    .B1(n_14293),
    .B2(n_91),
    .C1(n_3020),
    .C2(n_77),
    .Y(n_3135));
 INVxp33_ASAP7_75t_R g35635 (.A(n_2953),
    .Y(n_3541));
 OAI22xp33_ASAP7_75t_L g35638__6260 (.A1(n_73),
    .A2(n_3052),
    .B1(n_72),
    .B2(n_2945),
    .Y(n_3133));
 AOI222xp33_ASAP7_75t_R g35640__4319 (.A1(n_2949),
    .A2(n_2907),
    .B1(n_2936),
    .B2(n_14106),
    .C1(n_2934),
    .C2(n_14108),
    .Y(n_3132));
 AOI221xp5_ASAP7_75t_R g35642__5526 (.A1(n_2931),
    .A2(n_14166),
    .B1(n_2938),
    .B2(n_14108),
    .C(n_3025),
    .Y(n_3130));
 OAI221xp5_ASAP7_75t_R g35643__6783 (.A1(n_2945),
    .A2(n_82),
    .B1(n_2932),
    .B2(n_80),
    .C(n_3042),
    .Y(n_3129));
 OAI221xp5_ASAP7_75t_R g35644__3680 (.A1(n_3045),
    .A2(n_74),
    .B1(n_2932),
    .B2(n_79),
    .C(n_3028),
    .Y(n_3128));
 OAI221xp5_ASAP7_75t_R g35645__1617 (.A1(n_2945),
    .A2(n_78),
    .B1(n_2932),
    .B2(n_82),
    .C(n_3027),
    .Y(n_3127));
 AOI222xp33_ASAP7_75t_R g35646__2802 (.A1(n_2949),
    .A2(n_14090),
    .B1(n_2936),
    .B2(n_14102),
    .C1(n_2934),
    .C2(n_2896),
    .Y(n_3126));
 AOI222xp33_ASAP7_75t_R g35647__1705 (.A1(n_2882),
    .A2(n_14096),
    .B1(n_2931),
    .B2(n_14090),
    .C1(n_2877),
    .C2(n_2907),
    .Y(n_3125));
 AOI21xp33_ASAP7_75t_R g35648__5122 (.A1(n_2939),
    .A2(n_14106),
    .B(n_3066),
    .Y(n_3124));
 AOI222xp33_ASAP7_75t_R g35649__8246 (.A1(n_2939),
    .A2(n_14102),
    .B1(n_2936),
    .B2(n_14110),
    .C1(n_2934),
    .C2(n_14112),
    .Y(n_3123));
 OAI222xp33_ASAP7_75t_R g35650__7098 (.A1(n_2935),
    .A2(n_84),
    .B1(n_14294),
    .B2(n_2887),
    .C1(n_3034),
    .C2(n_77),
    .Y(n_3122));
 AOI222xp33_ASAP7_75t_R g35651__6131 (.A1(n_2938),
    .A2(n_14090),
    .B1(n_2934),
    .B2(n_14098),
    .C1(n_2930),
    .C2(n_14102),
    .Y(n_3121));
 AOI222xp33_ASAP7_75t_R g35652__1881 (.A1(n_2934),
    .A2(n_14090),
    .B1(n_2936),
    .B2(n_14088),
    .C1(n_2930),
    .C2(n_2907),
    .Y(n_3120));
 AOI222xp33_ASAP7_75t_R g35653__5115 (.A1(n_2936),
    .A2(n_2896),
    .B1(n_2934),
    .B2(n_14106),
    .C1(n_2939),
    .C2(n_14096),
    .Y(n_3119));
 AOI222xp33_ASAP7_75t_R g35654__7482 (.A1(n_2936),
    .A2(n_14092),
    .B1(n_2930),
    .B2(n_14098),
    .C1(n_2934),
    .C2(n_2907),
    .Y(n_3118));
 AOI222xp33_ASAP7_75t_R g35655__4733 (.A1(n_2939),
    .A2(n_14092),
    .B1(n_2936),
    .B2(n_2888),
    .C1(n_2934),
    .C2(n_14102),
    .Y(n_3117));
 AOI222xp33_ASAP7_75t_R g35656__6161 (.A1(n_2939),
    .A2(n_14090),
    .B1(n_2936),
    .B2(n_14098),
    .C1(n_2934),
    .C2(n_2888),
    .Y(n_3116));
 NAND2xp33_ASAP7_75t_R g35657__9315 (.A(n_3014),
    .B(n_2952),
    .Y(n_3545));
 NAND2xp33_ASAP7_75t_R g35658__9945 (.A(n_2988),
    .B(n_2952),
    .Y(n_3847));
 NAND2xp33_ASAP7_75t_R g35659__2883 (.A(n_14092),
    .B(n_2952),
    .Y(n_3846));
 AND4x1_ASAP7_75t_R g35660__2346 (.A(n_3037),
    .B(n_2937),
    .C(n_79),
    .D(n_2896),
    .Y(n_2953));
 OAI221xp5_ASAP7_75t_R g35661__1666 (.A1(n_3045),
    .A2(n_80),
    .B1(n_2932),
    .B2(n_73),
    .C(n_3039),
    .Y(n_3115));
 AOI221xp5_ASAP7_75t_R g35662__7410 (.A1(n_2938),
    .A2(n_14106),
    .B1(n_2931),
    .B2(n_14116),
    .C(n_3041),
    .Y(n_3114));
 OAI22xp33_ASAP7_75t_R g35663__6417 (.A1(n_89),
    .A2(n_3052),
    .B1(n_73),
    .B2(n_2945),
    .Y(n_3113));
 AOI22xp33_ASAP7_75t_R g35664__5477 (.A1(n_3047),
    .A2(n_14088),
    .B1(n_2947),
    .B2(n_14098),
    .Y(n_3112));
 AOI22xp33_ASAP7_75t_R g35665__2398 (.A1(n_2888),
    .A2(n_3047),
    .B1(n_14110),
    .B2(n_2947),
    .Y(n_3111));
 AOI22xp33_ASAP7_75t_R g35666__5107 (.A1(n_14108),
    .A2(n_2947),
    .B1(n_14110),
    .B2(n_2946),
    .Y(n_3110));
 OAI22xp33_ASAP7_75t_L g35667__6260 (.A1(n_89),
    .A2(n_14294),
    .B1(n_73),
    .B2(n_3045),
    .Y(n_3109));
 AOI22xp33_ASAP7_75t_R g35668__4319 (.A1(n_14106),
    .A2(n_2947),
    .B1(n_14108),
    .B2(n_2946),
    .Y(n_3108));
 AOI221xp5_ASAP7_75t_SL g35669__8428 (.A1(n_2931),
    .A2(n_14170),
    .B1(n_2938),
    .B2(n_14112),
    .C(n_3043),
    .Y(n_3107));
 AOI22xp33_ASAP7_75t_R g35670__5526 (.A1(n_14112),
    .A2(n_2946),
    .B1(n_14168),
    .B2(n_2930),
    .Y(n_3106));
 AOI22xp33_ASAP7_75t_R g35671__6783 (.A1(n_14092),
    .A2(n_2947),
    .B1(n_2907),
    .B2(n_2946),
    .Y(n_3105));
 OAI22xp5_ASAP7_75t_L g35672__3680 (.A1(n_80),
    .A2(n_14293),
    .B1(n_84),
    .B2(n_3053),
    .Y(n_3104));
 AOI22xp33_ASAP7_75t_R g35673__1617 (.A1(n_14088),
    .A2(n_2938),
    .B1(n_2907),
    .B2(n_2936),
    .Y(n_3103));
 OAI22xp33_ASAP7_75t_R g35674__2802 (.A1(n_90),
    .A2(n_14293),
    .B1(n_80),
    .B2(n_3055),
    .Y(n_3102));
 OAI22xp5_ASAP7_75t_L g35675__1705 (.A1(n_79),
    .A2(n_3055),
    .B1(n_77),
    .B2(n_14294),
    .Y(n_3101));
 AOI22xp33_ASAP7_75t_R g35676__5122 (.A1(n_14106),
    .A2(n_2946),
    .B1(n_14114),
    .B2(n_2930),
    .Y(n_3100));
 AOI22xp33_ASAP7_75t_R g35677__8246 (.A1(n_14088),
    .A2(n_2946),
    .B1(n_2907),
    .B2(n_2931),
    .Y(n_3099));
 OAI22xp5_ASAP7_75t_L g35678__7098 (.A1(n_79),
    .A2(n_3053),
    .B1(n_84),
    .B2(n_14294),
    .Y(n_3098));
 OAI22xp33_ASAP7_75t_R g35679__6131 (.A1(n_82),
    .A2(n_14293),
    .B1(n_90),
    .B2(n_3053),
    .Y(n_3097));
 AOI22xp33_ASAP7_75t_R g35680__1881 (.A1(n_2888),
    .A2(n_2949),
    .B1(n_2896),
    .B2(n_2939),
    .Y(n_3096));
 AOI22xp5_ASAP7_75t_SL g35681__5115 (.A1(n_14108),
    .A2(n_2949),
    .B1(n_14110),
    .B2(n_3054),
    .Y(n_3095));
 AOI22xp33_ASAP7_75t_R g35682__7482 (.A1(n_2888),
    .A2(n_2946),
    .B1(n_14108),
    .B2(n_2930),
    .Y(n_3094));
 AOI22xp33_ASAP7_75t_R g35683__4733 (.A1(n_2949),
    .A2(n_14088),
    .B1(n_2948),
    .B2(n_14090),
    .Y(n_3093));
 AOI22xp33_ASAP7_75t_R g35684__6161 (.A1(n_2948),
    .A2(n_14096),
    .B1(n_2939),
    .B2(n_14098),
    .Y(n_3092));
 INVx1_ASAP7_75t_R g35690 (.A(n_2952),
    .Y(n_3848));
 INVxp33_ASAP7_75t_R g35691 (.A(n_3091),
    .Y(n_3090));
 INVxp67_ASAP7_75t_R g35692 (.A(n_3089),
    .Y(n_3088));
 INVxp33_ASAP7_75t_R g35695 (.A(n_3849),
    .Y(n_3087));
 INVxp33_ASAP7_75t_R g35699 (.A(n_2950),
    .Y(n_2951));
 INVxp33_ASAP7_75t_R g35702 (.A(n_3543),
    .Y(n_3086));
 INVx1_ASAP7_75t_R g35707 (.A(n_3084),
    .Y(n_3083));
 NOR2xp33_ASAP7_75t_R g35708__9315 (.A(n_3049),
    .B(n_88),
    .Y(n_3626));
 NAND2xp33_ASAP7_75t_R g35709__9945 (.A(n_2888),
    .B(fracta_mul[23]),
    .Y(n_3082));
 NOR2xp33_ASAP7_75t_R g35710__2883 (.A(n_2941),
    .B(n_86),
    .Y(n_3081));
 NAND2xp33_ASAP7_75t_R g35711__2346 (.A(n_2944),
    .B(n_14118),
    .Y(n_3080));
 NAND2xp33_ASAP7_75t_R g35712__1666 (.A(n_14110),
    .B(n_2938),
    .Y(n_3079));
 NAND2xp33_ASAP7_75t_R g35713__7410 (.A(n_2944),
    .B(n_14120),
    .Y(n_3078));
 NAND3xp33_ASAP7_75t_R g35714__6417 (.A(n_3037),
    .B(n_2937),
    .C(n_2896),
    .Y(n_3077));
 AND2x2_ASAP7_75t_L g35716__5477 (.A(n_3021),
    .B(n_3057),
    .Y(n_2952));
 NAND2xp5_ASAP7_75t_R g35717__2398 (.A(n_2941),
    .B(n_14092),
    .Y(n_3091));
 NAND2xp5_ASAP7_75t_R g35718__5107 (.A(n_2941),
    .B(n_14090),
    .Y(n_3089));
 NAND2xp5_ASAP7_75t_L g35719__6260 (.A(n_2888),
    .B(n_3057),
    .Y(n_3849));
 NAND3xp33_ASAP7_75t_SL g35720__4319 (.A(n_3037),
    .B(n_2937),
    .C(n_3019),
    .Y(n_2950));
 NAND3xp33_ASAP7_75t_L g35721__234781 (.A(n_3037),
    .B(n_2937),
    .C(n_14106),
    .Y(n_3543));
 NAND2xp5_ASAP7_75t_SL g35723__6783 (.A(n_2941),
    .B(n_14088),
    .Y(n_3084));
 INVxp33_ASAP7_75t_R g35724 (.A(u1_n_590),
    .Y(n_3074));
 INVxp67_ASAP7_75t_L g35732 (.A(n_3070),
    .Y(n_3071));
 AOI22xp33_ASAP7_75t_R g35733__3680 (.A1(n_14112),
    .A2(n_2936),
    .B1(n_14114),
    .B2(n_2934),
    .Y(n_3069));
 AOI221xp5_ASAP7_75t_L g35734__1617 (.A1(n_2930),
    .A2(n_14170),
    .B1(n_2931),
    .B2(n_14168),
    .C(n_3031),
    .Y(n_3068));
 OAI221xp5_ASAP7_75t_R g35735__2802 (.A1(n_2932),
    .A2(n_86),
    .B1(n_13839),
    .B2(n_85),
    .C(n_3022),
    .Y(n_3067));
 OAI22xp33_ASAP7_75t_R g35736__1705 (.A1(n_73),
    .A2(n_2935),
    .B1(n_72),
    .B2(n_3034),
    .Y(n_3066));
 OAI22xp33_ASAP7_75t_R g35737__5122 (.A1(n_72),
    .A2(n_2935),
    .B1(n_81),
    .B2(n_3034),
    .Y(n_3065));
 AOI222xp33_ASAP7_75t_R g35738__8246 (.A1(n_2931),
    .A2(n_2888),
    .B1(n_2877),
    .B2(n_2896),
    .C1(n_2882),
    .C2(n_14106),
    .Y(n_3064));
 AOI222xp33_ASAP7_75t_R g35739__7098 (.A1(n_2931),
    .A2(n_14096),
    .B1(n_2877),
    .B2(n_2888),
    .C1(n_2882),
    .C2(n_14102),
    .Y(n_3063));
 AOI222xp33_ASAP7_75t_R g35740__6131 (.A1(n_2931),
    .A2(n_14112),
    .B1(n_2877),
    .B2(n_14116),
    .C1(n_2882),
    .C2(n_14166),
    .Y(n_3062));
 OAI222xp33_ASAP7_75t_R g35741__1881 (.A1(n_73),
    .A2(n_2928),
    .B1(n_77),
    .B2(n_2932),
    .C1(n_72),
    .C2(n_76),
    .Y(n_3061));
 AOI222xp33_ASAP7_75t_R g35742__5115 (.A1(n_2931),
    .A2(n_14092),
    .B1(n_2877),
    .B2(n_14096),
    .C1(n_2882),
    .C2(n_14098),
    .Y(n_3060));
 AOI222xp33_ASAP7_75t_R g35743__7482 (.A1(n_2931),
    .A2(n_14108),
    .B1(n_2877),
    .B2(n_14112),
    .C1(n_2882),
    .C2(n_14114),
    .Y(n_3059));
 OAI22xp33_ASAP7_75t_R g35744__4733 (.A1(n_81),
    .A2(n_2935),
    .B1(n_95),
    .B2(n_3034),
    .Y(n_3058));
 XNOR2xp5_ASAP7_75t_R g35745__6161 (.A(u1_n_5382),
    .B(opa_r[31]),
    .Y(u1_n_590));
 NAND2xp5_ASAP7_75t_L g35746__9315 (.A(n_3009),
    .B(n_3057),
    .Y(n_3845));
 NAND2xp5_ASAP7_75t_L g35747__9945 (.A(n_3016),
    .B(n_3057),
    .Y(n_3844));
 NAND2xp5_ASAP7_75t_SL g35748__2883 (.A(n_2990),
    .B(n_3057),
    .Y(n_3070));
 INVxp33_ASAP7_75t_R g35749 (.A(n_3057),
    .Y(u0_n_321));
 INVxp67_ASAP7_75t_R g35759 (.A(n_3055),
    .Y(n_2949));
 INVxp67_ASAP7_75t_L g35762 (.A(n_3053),
    .Y(n_3054));
 INVxp33_ASAP7_75t_R g35766 (.A(n_3053),
    .Y(n_2948));
 INVx1_ASAP7_75t_R g35787 (.A(n_2947),
    .Y(n_3052));
 INVxp67_ASAP7_75t_R g35806 (.A(n_3049),
    .Y(fracta_mul[23]));
 HB1xp67_ASAP7_75t_R g35821 (.A(n_2941),
    .Y(n_3049));
 INVxp67_ASAP7_75t_R g35822 (.A(n_2941),
    .Y(n_2942));
 BUFx2_ASAP7_75t_L g35829 (.A(n_2940),
    .Y(n_2941));
 OR5x1_ASAP7_75t_L g35842__2346 (.A(n_3029),
    .B(opb_r[23]),
    .C(opb_r[30]),
    .D(opb_r[26]),
    .E(opb_r[29]),
    .Y(fractb_mul[23]));
 AND2x2_ASAP7_75t_SL g35843__1666 (.A(n_3030),
    .B(n_3037),
    .Y(n_3057));
 NAND2x1p5_ASAP7_75t_SL g35844__7410 (.A(n_3010),
    .B(n_3037),
    .Y(n_3055));
 NAND2xp5_ASAP7_75t_L g35845__6417 (.A(n_3018),
    .B(n_3037),
    .Y(n_3053));
 AND3x2_ASAP7_75t_SL g35846__5477 (.A(n_3012),
    .B(n_3005),
    .C(n_2983),
    .Y(n_2947));
 AND3x1_ASAP7_75t_R g35847__2398 (.A(n_3012),
    .B(n_3005),
    .C(n_14168),
    .Y(n_2946));
 NAND4xp25_ASAP7_75t_R g35848__5107 (.A(n_3001),
    .B(n_3007),
    .C(n_3005),
    .D(n_14168),
    .Y(n_2945));
 NOR5xp2_ASAP7_75t_SL g35849__6260 (.A(n_3024),
    .B(opa_r[28]),
    .C(opa_r[29]),
    .D(opa_r[23]),
    .E(opa_r[27]),
    .Y(n_2943));
 INVxp33_ASAP7_75t_R g35850 (.A(n_14293),
    .Y(n_3047));
 INVxp67_ASAP7_75t_R g35869 (.A(n_14294),
    .Y(n_2939));
 INVxp67_ASAP7_75t_R g35881 (.A(n_2938),
    .Y(n_3045));
 OAI221xp5_ASAP7_75t_R g35883__4319 (.A1(n_3020),
    .A2(n_86),
    .B1(n_2928),
    .B2(n_85),
    .C(n_2992),
    .Y(n_3043));
 AOI222xp33_ASAP7_75t_R g35884__8428 (.A1(n_2930),
    .A2(n_14106),
    .B1(n_2877),
    .B2(n_14108),
    .C1(n_2882),
    .C2(n_14110),
    .Y(n_3042));
 OAI221xp5_ASAP7_75t_R g35885__5526 (.A1(n_3020),
    .A2(n_81),
    .B1(n_2928),
    .B2(n_95),
    .C(n_2989),
    .Y(n_3041));
 AOI222xp33_ASAP7_75t_R g35886__6783 (.A1(n_2930),
    .A2(n_2896),
    .B1(n_2877),
    .B2(n_14106),
    .C1(n_2882),
    .C2(n_14108),
    .Y(n_3040));
 AOI222xp33_ASAP7_75t_R g35887__3680 (.A1(n_2930),
    .A2(n_14116),
    .B1(n_2877),
    .B2(n_14166),
    .C1(n_2882),
    .C2(n_14168),
    .Y(n_3039));
 AND2x2_ASAP7_75t_L g35890__1705 (.A(n_3008),
    .B(n_3023),
    .Y(n_2938));
 INVxp67_ASAP7_75t_R g35907 (.A(n_2935),
    .Y(n_2936));
 INVxp67_ASAP7_75t_R g35909 (.A(n_3035),
    .Y(n_2935));
 INVxp67_ASAP7_75t_L g35928 (.A(n_2934),
    .Y(n_3034));
 INVxp33_ASAP7_75t_R g35930 (.A(n_2931),
    .Y(n_3840));
 INVxp67_ASAP7_75t_SL g35944 (.A(n_2932),
    .Y(n_2931));
 AND3x1_ASAP7_75t_L g35945__5122 (.A(n_2997),
    .B(n_2999),
    .C(n_84),
    .Y(n_2937));
 OAI21xp33_ASAP7_75t_R g35946__8246 (.A1(n_86),
    .A2(n_2928),
    .B(n_2993),
    .Y(n_3031));
 NOR3xp33_ASAP7_75t_L g35948__7098 (.A(n_3011),
    .B(n_2879),
    .C(n_2878),
    .Y(n_3030));
 AND2x4_ASAP7_75t_SL g35949__6131 (.A(n_3017),
    .B(n_3012),
    .Y(n_3037));
 NOR3xp33_ASAP7_75t_R g35950__1881 (.A(n_2984),
    .B(n_2991),
    .C(n_3002),
    .Y(n_3035));
 AND5x1_ASAP7_75t_SL g35951__5115 (.A(n_96),
    .B(n_76),
    .C(n_85),
    .D(n_93),
    .E(n_14172),
    .Y(n_2934));
 NAND4xp25_ASAP7_75t_SL g35952__7482 (.A(n_96),
    .B(n_76),
    .C(n_14174),
    .D(n_93),
    .Y(n_2932));
 OR4x1_ASAP7_75t_L g35953__4733 (.A(opb_r[27]),
    .B(opb_r[25]),
    .C(opb_r[28]),
    .D(opb_r[24]),
    .Y(n_3029));
 AOI22xp33_ASAP7_75t_R g35954__6161 (.A1(n_14110),
    .A2(n_2877),
    .B1(n_14112),
    .B2(n_2882),
    .Y(n_3028));
 AOI22xp33_ASAP7_75t_R g35955__9315 (.A1(n_14102),
    .A2(n_2877),
    .B1(n_2896),
    .B2(n_2882),
    .Y(n_3027));
 AOI22xp33_ASAP7_75t_R g35956__9945 (.A1(n_14098),
    .A2(n_2877),
    .B1(n_2882),
    .B2(n_2888),
    .Y(n_3026));
 OAI22xp33_ASAP7_75t_R g35957__2883 (.A1(n_83),
    .A2(n_2928),
    .B1(n_86),
    .B2(n_76),
    .Y(n_3025));
 OR4x1_ASAP7_75t_L g35958__2346 (.A(opa_r[30]),
    .B(opa_r[25]),
    .C(opa_r[26]),
    .D(opa_r[24]),
    .Y(n_3024));
 NOR3xp33_ASAP7_75t_L g35959__1666 (.A(n_3002),
    .B(n_2982),
    .C(n_14176),
    .Y(n_3023));
 AOI21xp33_ASAP7_75t_R g35960__7410 (.A1(n_14120),
    .A2(n_14118),
    .B(n_2986),
    .Y(n_3022));
 XOR2xp5_ASAP7_75t_R g35961__6417 (.A(opb_r[31]),
    .B(fpu_op_r1[0]),
    .Y(u1_n_5382));
 INVxp33_ASAP7_75t_R g35962 (.A(n_3021),
    .Y(n_3544));
 INVx1_ASAP7_75t_R g35981 (.A(n_3020),
    .Y(n_2930));
 NOR2xp33_ASAP7_75t_R g35982__5477 (.A(n_90),
    .B(n_3570),
    .Y(n_3019));
 NOR2xp33_ASAP7_75t_R g35983__2398 (.A(n_89),
    .B(n_2879),
    .Y(n_3018));
 NOR2xp33_ASAP7_75t_SL g35984__5107 (.A(n_2995),
    .B(n_3003),
    .Y(n_3017));
 NOR2xp33_ASAP7_75t_R g35985__6260 (.A(n_74),
    .B(n_2998),
    .Y(n_3016));
 NOR2xp33_ASAP7_75t_L g35986__4319 (.A(n_3566),
    .B(n_2998),
    .Y(n_3021));
 NAND3xp33_ASAP7_75t_L g35988__5526 (.A(n_96),
    .B(n_76),
    .C(n_14118),
    .Y(n_3020));
 NAND2xp33_ASAP7_75t_R g35990__6783 (.A(n_2929),
    .B(n_2996),
    .Y(n_3011));
 AND3x1_ASAP7_75t_R g35991__3680 (.A(n_78),
    .B(n_88),
    .C(n_91),
    .Y(n_3014));
 NOR2xp33_ASAP7_75t_L g35992__1617 (.A(n_2987),
    .B(n_2879),
    .Y(n_3010));
 NOR2xp33_ASAP7_75t_R g35993__2802 (.A(n_2994),
    .B(n_2998),
    .Y(n_3009));
 NOR4xp25_ASAP7_75t_R g35994__1705 (.A(n_14166),
    .B(n_14118),
    .C(n_14170),
    .D(n_14172),
    .Y(n_3008));
 NOR2xp67_ASAP7_75t_SL g35995__5122 (.A(n_3000),
    .B(n_2880),
    .Y(n_3012));
 INVxp33_ASAP7_75t_R g35996 (.A(n_2880),
    .Y(n_3007));
 INVx1_ASAP7_75t_R g35998 (.A(n_3003),
    .Y(n_3005));
 NAND2xp5_ASAP7_75t_SL g36003__8246 (.A(n_86),
    .B(n_83),
    .Y(n_3003));
 NAND2xp5_ASAP7_75t_R g36014__7098 (.A(n_96),
    .B(n_85),
    .Y(n_3002));
 INVxp33_ASAP7_75t_R g36022 (.A(n_3000),
    .Y(n_3001));
 INVxp67_ASAP7_75t_L g36023 (.A(n_2878),
    .Y(n_2999));
 INVxp33_ASAP7_75t_R g36026 (.A(n_2929),
    .Y(n_3570));
 INVx1_ASAP7_75t_R g36029 (.A(n_2879),
    .Y(n_2997));
 INVxp33_ASAP7_75t_R g36045 (.A(n_2928),
    .Y(n_2877));
 NOR2xp33_ASAP7_75t_R g36051__6131 (.A(n_14102),
    .B(n_14108),
    .Y(n_2996));
 NAND2xp5_ASAP7_75t_SL g36052__1881 (.A(n_95),
    .B(n_81),
    .Y(n_2995));
 NAND2xp33_ASAP7_75t_R g36053__5115 (.A(n_14094),
    .B(n_74),
    .Y(n_2994));
 NAND2xp33_ASAP7_75t_R g36054__7482 (.A(n_14174),
    .B(n_2882),
    .Y(n_2993));
 NAND2xp5_ASAP7_75t_SL g36055__4733 (.A(n_85),
    .B(n_76),
    .Y(n_3000));
 NAND2xp33_ASAP7_75t_R g36056__6161 (.A(n_14118),
    .B(n_14176),
    .Y(n_2992));
 NAND2xp33_ASAP7_75t_R g36057__9315 (.A(n_76),
    .B(n_93),
    .Y(n_2991));
 NOR2xp33_ASAP7_75t_R g36058__9945 (.A(n_2888),
    .B(n_82),
    .Y(n_2990));
 NAND2xp33_ASAP7_75t_R g36059__2883 (.A(n_14170),
    .B(n_2882),
    .Y(n_2989));
 NOR2xp33_ASAP7_75t_R g36060__2346 (.A(n_91),
    .B(n_14092),
    .Y(n_2988));
 NAND2xp5_ASAP7_75t_R g36061__1666 (.A(n_14110),
    .B(n_89),
    .Y(n_2987));
 NOR2xp33_ASAP7_75t_R g36062__7410 (.A(n_96),
    .B(n_76),
    .Y(n_2986));
 NAND2xp33_ASAP7_75t_R g36064__5477 (.A(n_86),
    .B(n_14170),
    .Y(n_2984));
 NOR2xp33_ASAP7_75t_R g36065__2398 (.A(n_81),
    .B(n_14168),
    .Y(n_2983));
 NAND2xp33_ASAP7_75t_R g36066__5107 (.A(n_14116),
    .B(n_95),
    .Y(n_2982));
 NAND2xp5_ASAP7_75t_R g36067__6260 (.A(n_74),
    .B(n_87),
    .Y(n_3566));
 NOR2xp33_ASAP7_75t_L g36069__4319 (.A(n_2896),
    .B(n_14106),
    .Y(n_2929));
 OR2x2_ASAP7_75t_R g36070__8428 (.A(n_14100),
    .B(n_14098),
    .Y(n_2998));
 INVxp33_ASAP7_75t_R g36074 (.A(opb[30]),
    .Y(n_2980));
 INVxp33_ASAP7_75t_R g36075 (.A(opa[27]),
    .Y(n_2979));
 INVxp33_ASAP7_75t_R g36076 (.A(opa[30]),
    .Y(n_2978));
 INVxp33_ASAP7_75t_R g36077 (.A(opa[28]),
    .Y(n_2977));
 INVxp33_ASAP7_75t_R g36078 (.A(opa[29]),
    .Y(n_2976));
 INVxp33_ASAP7_75t_R g36079 (.A(opa[26]),
    .Y(n_2975));
 INVxp33_ASAP7_75t_R g36080 (.A(opb[28]),
    .Y(n_2974));
 INVxp33_ASAP7_75t_R g36081 (.A(opb[24]),
    .Y(n_2973));
 INVxp33_ASAP7_75t_R g36082 (.A(opb[23]),
    .Y(n_2972));
 INVxp33_ASAP7_75t_R g36083 (.A(opb[27]),
    .Y(n_2971));
 INVx1_ASAP7_75t_L g36087 (.A(n_14120),
    .Y(n_96));
 INVx1_ASAP7_75t_L g36099 (.A(n_14170),
    .Y(n_83));
 INVx1_ASAP7_75t_R g36103 (.A(n_14172),
    .Y(n_86));
 INVx1_ASAP7_75t_L g36121 (.A(n_14168),
    .Y(n_95));
 INVxp33_ASAP7_75t_R g36130 (.A(n_14114),
    .Y(n_73));
 INVxp67_ASAP7_75t_R g36142 (.A(n_14116),
    .Y(n_72));
 INVxp67_ASAP7_75t_R g36145 (.A(n_14088),
    .Y(n_88));
 INVxp67_ASAP7_75t_L g36169 (.A(n_14112),
    .Y(n_89));
 INVx1_ASAP7_75t_R g36170 (.A(n_14092),
    .Y(n_78));
 INVxp67_ASAP7_75t_R g36190 (.A(n_14098),
    .Y(n_82));
 INVxp33_ASAP7_75t_R g36208 (.A(n_2907),
    .Y(n_2908));
 HB1xp67_ASAP7_75t_L g36209 (.A(n_14094),
    .Y(n_2907));
 INVxp33_ASAP7_75t_R g36210 (.A(opa[31]),
    .Y(n_2964));
 INVxp33_ASAP7_75t_R g36211 (.A(opa[25]),
    .Y(n_2963));
 INVxp33_ASAP7_75t_R g36212 (.A(opa[24]),
    .Y(n_2962));
 INVxp33_ASAP7_75t_R g36213 (.A(opb[31]),
    .Y(n_2961));
 INVxp33_ASAP7_75t_R g36214 (.A(opb[26]),
    .Y(n_2960));
 INVxp33_ASAP7_75t_R g36215 (.A(opb[25]),
    .Y(n_2959));
 INVxp33_ASAP7_75t_R g36216 (.A(opa[23]),
    .Y(n_2958));
 INVxp33_ASAP7_75t_R g36217 (.A(opb[29]),
    .Y(n_2957));
 INVxp67_ASAP7_75t_SL g36220 (.A(n_14174),
    .Y(n_85));
 INVx1_ASAP7_75t_L g36230 (.A(n_14118),
    .Y(n_93));
 INVx1_ASAP7_75t_L g36245 (.A(n_14166),
    .Y(n_81));
 INVxp33_ASAP7_75t_R g36246 (.A(n_14110),
    .Y(n_77));
 INVxp67_ASAP7_75t_R g36270 (.A(n_2896),
    .Y(n_80));
 INVx1_ASAP7_75t_L g36289 (.A(n_14108),
    .Y(n_84));
 INVxp67_ASAP7_75t_R g36302 (.A(n_14106),
    .Y(n_79));
 INVxp33_ASAP7_75t_R g36322 (.A(n_14090),
    .Y(n_91));
 INVxp67_ASAP7_75t_R g36338 (.A(n_14102),
    .Y(n_90));
 INVxp33_ASAP7_75t_R g36359 (.A(n_2888),
    .Y(n_2887));
 HB1xp67_ASAP7_75t_SL g36360 (.A(n_14100),
    .Y(n_2888));
 INVx1_ASAP7_75t_L g36379 (.A(n_14096),
    .Y(n_74));
 INVx1_ASAP7_75t_R g36404 (.A(n_76),
    .Y(n_2882));
 INVx2_ASAP7_75t_SL g36405 (.A(n_14176),
    .Y(n_76));
 OR2x2_ASAP7_75t_R g36419__6783 (.A(n_96),
    .B(n_14176),
    .Y(n_2928));
 OR2x2_ASAP7_75t_R g36420__3680 (.A(n_14118),
    .B(n_14120),
    .Y(n_2880));
 OR2x2_ASAP7_75t_L g36421__1617 (.A(n_14116),
    .B(n_14114),
    .Y(n_2879));
 OR2x2_ASAP7_75t_L g36422__2802 (.A(n_14112),
    .B(n_14110),
    .Y(n_2878));
 AOI311xp33_ASAP7_75t_R g36596 (.A1(n_604),
    .A2(n_3755),
    .A3(opas_r2),
    .B(n_615),
    .C(n_618),
    .Y(n_619));
 OAI321xp33_ASAP7_75t_R g36597 (.A1(n_617),
    .A2(n_599),
    .A3(n_230),
    .B1(sign_mul_r),
    .B2(n_345),
    .C(n_367),
    .Y(n_618));
 OR3x1_ASAP7_75t_R g36599 (.A(n_611),
    .B(n_612),
    .C(n_379),
    .Y(n_617));
 O2A1O1Ixp33_ASAP7_75t_R g36600 (.A1(n_253),
    .A2(n_360),
    .B(n_533),
    .C(n_614),
    .Y(n_616));
 AO22x1_ASAP7_75t_R g36601 (.A1(n_608),
    .A2(n_611),
    .B1(nan_sign_d),
    .B2(n_612),
    .Y(n_615));
 AOI211xp5_ASAP7_75t_R g36604 (.A1(n_607),
    .A2(n_603),
    .B(n_231),
    .C(inf_mul_r),
    .Y(n_614));
 AOI221xp5_ASAP7_75t_R g36606 (.A1(n_602),
    .A2(n_3596),
    .B1(n_296),
    .B2(opb_inf),
    .C(n_605),
    .Y(n_613));
 A2O1A1Ixp33_ASAP7_75t_R g36607 (.A1(n_114),
    .A2(n_600),
    .B(n_258),
    .C(n_47),
    .Y(n_610));
 OAI22xp33_ASAP7_75t_R g36608 (.A1(n_70),
    .A2(n_606),
    .B1(n_114),
    .B2(n_599),
    .Y(n_612));
 NOR3xp33_ASAP7_75t_R g36609 (.A(n_606),
    .B(n_113),
    .C(ind_d),
    .Y(n_611));
 AOI322xp5_ASAP7_75t_R g36610 (.A1(n_598),
    .A2(n_275),
    .A3(n_149),
    .B1(n_360),
    .B2(n_537),
    .C1(n_509),
    .C2(fpu_op_r3[2]),
    .Y(n_609));
 AO22x1_ASAP7_75t_R g36611 (.A1(result_zero_sign_d),
    .A2(n_602),
    .B1(sign_fasu_r),
    .B2(n_601),
    .Y(n_608));
 NAND4xp25_ASAP7_75t_R g36612 (.A(n_596),
    .B(n_473),
    .C(u4_op_dn),
    .D(sign),
    .Y(n_607));
 AO21x1_ASAP7_75t_R g36613 (.A1(n_333),
    .A2(n_596),
    .B(n_604),
    .Y(n_605));
 OR3x1_ASAP7_75t_R g36614 (.A(n_599),
    .B(n_22),
    .C(n_23),
    .Y(n_606));
 O2A1O1Ixp33_ASAP7_75t_R g36615 (.A1(n_531),
    .A2(n_594),
    .B(underflow_fmul_r[2]),
    .C(underflow_fmul_r[0]),
    .Y(n_603));
 AND2x2_ASAP7_75t_R g36616 (.A(n_114),
    .B(n_599),
    .Y(n_604));
 INVxp33_ASAP7_75t_R g36617 (.A(n_602),
    .Y(n_601));
 OAI311xp33_ASAP7_75t_R g36618 (.A1(fpu_op_r3[1]),
    .A2(n_35),
    .A3(n_148),
    .B1(n_595),
    .C1(n_363),
    .Y(n_600));
 NOR3xp33_ASAP7_75t_R g36619 (.A(n_597),
    .B(n_113),
    .C(inf_d),
    .Y(n_602));
 NOR2xp33_ASAP7_75t_R g36620 (.A(n_3803),
    .B(n_597),
    .Y(n_599));
 NAND3xp33_ASAP7_75t_R g36621 (.A(n_597),
    .B(n_540),
    .C(n_363),
    .Y(n_598));
 INVxp33_ASAP7_75t_R g36622 (.A(n_597),
    .Y(n_596));
 NAND2xp33_ASAP7_75t_R g36623 (.A(n_531),
    .B(n_594),
    .Y(n_597));
 NAND2xp33_ASAP7_75t_R g36624 (.A(n_530),
    .B(n_594),
    .Y(n_595));
 NOR5xp2_ASAP7_75t_R g36625 (.A(n_593),
    .B(n_592),
    .C(n_587),
    .D(n_588),
    .E(n_589),
    .Y(n_594));
 NAND5xp2_ASAP7_75t_R g36628 (.A(n_591),
    .B(n_551),
    .C(n_552),
    .D(n_554),
    .E(n_550),
    .Y(n_593));
 NAND4xp25_ASAP7_75t_R g36642 (.A(n_545),
    .B(n_562),
    .C(n_564),
    .D(n_560),
    .Y(n_592));
 AND3x1_ASAP7_75t_R g36650 (.A(n_546),
    .B(n_548),
    .C(n_547),
    .Y(n_591));
 AOI21xp33_ASAP7_75t_R g36651 (.A1(n_544),
    .A2(n_13),
    .B(n_395),
    .Y(n_590));
 NAND4xp25_ASAP7_75t_R g36652 (.A(n_542),
    .B(n_559),
    .C(n_557),
    .D(n_558),
    .Y(n_589));
 NAND4xp25_ASAP7_75t_R g36653 (.A(n_556),
    .B(n_555),
    .C(n_553),
    .D(n_549),
    .Y(n_588));
 NAND4xp25_ASAP7_75t_R g36654 (.A(n_563),
    .B(n_543),
    .C(n_565),
    .D(n_561),
    .Y(n_587));
 OR2x2_ASAP7_75t_R g36656 (.A(n_8),
    .B(n_557),
    .Y(n_586));
 OR2x2_ASAP7_75t_R g36657 (.A(n_381),
    .B(n_549),
    .Y(n_585));
 OR2x2_ASAP7_75t_R g36658 (.A(n_8),
    .B(n_554),
    .Y(n_584));
 OR2x2_ASAP7_75t_R g36659 (.A(n_8),
    .B(n_546),
    .Y(n_583));
 OR2x2_ASAP7_75t_R g36660 (.A(n_381),
    .B(n_550),
    .Y(n_582));
 OR2x2_ASAP7_75t_R g36661 (.A(n_8),
    .B(n_552),
    .Y(n_581));
 OR2x2_ASAP7_75t_R g36662 (.A(n_381),
    .B(n_561),
    .Y(n_580));
 OR2x2_ASAP7_75t_R g36663 (.A(n_8),
    .B(n_555),
    .Y(n_579));
 OR2x2_ASAP7_75t_R g36664 (.A(n_8),
    .B(n_562),
    .Y(n_578));
 OR2x2_ASAP7_75t_R g36665 (.A(n_381),
    .B(n_556),
    .Y(n_577));
 OR2x2_ASAP7_75t_R g36666 (.A(n_8),
    .B(n_563),
    .Y(n_576));
 OR2x2_ASAP7_75t_R g36667 (.A(n_8),
    .B(n_560),
    .Y(n_575));
 OR2x2_ASAP7_75t_R g36668 (.A(n_381),
    .B(n_565),
    .Y(n_574));
 OR2x2_ASAP7_75t_R g36669 (.A(n_381),
    .B(n_547),
    .Y(n_573));
 OR2x2_ASAP7_75t_R g36670 (.A(n_381),
    .B(n_548),
    .Y(n_572));
 OR2x2_ASAP7_75t_R g36671 (.A(n_8),
    .B(n_558),
    .Y(n_571));
 OR2x2_ASAP7_75t_R g36672 (.A(n_381),
    .B(n_551),
    .Y(n_570));
 OR2x2_ASAP7_75t_R g36673 (.A(n_8),
    .B(n_559),
    .Y(n_569));
 OR2x2_ASAP7_75t_R g36674 (.A(n_381),
    .B(n_564),
    .Y(n_568));
 OR2x2_ASAP7_75t_R g36675 (.A(n_381),
    .B(n_545),
    .Y(n_567));
 AO21x1_ASAP7_75t_R g36676 (.A1(n_15),
    .A2(n_542),
    .B(n_8),
    .Y(n_566));
 AOI221xp5_ASAP7_75t_R g36677 (.A1(n_541),
    .A2(u4_fract_out[15]),
    .B1(n_538),
    .B2(n_3792),
    .C(n_539),
    .Y(n_565));
 AOI221xp5_ASAP7_75t_R g36678 (.A1(n_541),
    .A2(u4_fract_out[20]),
    .B1(n_538),
    .B2(n_3797),
    .C(n_539),
    .Y(n_564));
 AOI221xp5_ASAP7_75t_R g36679 (.A1(n_541),
    .A2(u4_fract_out[17]),
    .B1(n_2),
    .B2(n_3794),
    .C(n_3),
    .Y(n_563));
 AOI221xp5_ASAP7_75t_R g36680 (.A1(n_5),
    .A2(u4_fract_out[10]),
    .B1(n_2),
    .B2(n_3787),
    .C(n_3),
    .Y(n_562));
 AOI221xp5_ASAP7_75t_R g36681 (.A1(n_5),
    .A2(u4_fract_out[8]),
    .B1(n_2),
    .B2(n_3785),
    .C(n_3),
    .Y(n_561));
 AOI221xp5_ASAP7_75t_R g36682 (.A1(n_5),
    .A2(u4_fract_out[14]),
    .B1(n_538),
    .B2(n_3791),
    .C(n_539),
    .Y(n_560));
 AOI221xp5_ASAP7_75t_R g36683 (.A1(n_5),
    .A2(u4_fract_out[19]),
    .B1(n_2),
    .B2(n_3796),
    .C(n_3),
    .Y(n_559));
 AOI221xp5_ASAP7_75t_R g36684 (.A1(n_5),
    .A2(u4_fract_out[13]),
    .B1(n_2),
    .B2(n_3790),
    .C(n_3),
    .Y(n_558));
 AOI221xp5_ASAP7_75t_R g36685 (.A1(n_5),
    .A2(u4_fract_out[2]),
    .B1(n_2),
    .B2(n_3779),
    .C(n_3),
    .Y(n_557));
 AOI221xp5_ASAP7_75t_R g36686 (.A1(n_5),
    .A2(u4_fract_out[11]),
    .B1(n_538),
    .B2(n_3788),
    .C(n_539),
    .Y(n_556));
 AOI221xp5_ASAP7_75t_R g36687 (.A1(n_541),
    .A2(u4_fract_out[9]),
    .B1(n_2),
    .B2(n_3786),
    .C(n_539),
    .Y(n_555));
 INVxp33_ASAP7_75t_R g36688 (.A(n_543),
    .Y(n_544));
 AOI221xp5_ASAP7_75t_R g36689 (.A1(n_5),
    .A2(u4_fract_out[1]),
    .B1(n_538),
    .B2(n_3778),
    .C(n_539),
    .Y(n_554));
 AOI221xp5_ASAP7_75t_R g36690 (.A1(n_541),
    .A2(u4_fract_out[22]),
    .B1(n_538),
    .B2(n_3799),
    .C(n_539),
    .Y(n_553));
 AOI221xp5_ASAP7_75t_R g36691 (.A1(n_541),
    .A2(u4_fract_out[6]),
    .B1(n_2),
    .B2(n_3783),
    .C(n_3),
    .Y(n_552));
 AOI221xp5_ASAP7_75t_R g36692 (.A1(n_5),
    .A2(u4_fract_out[18]),
    .B1(n_538),
    .B2(n_3795),
    .C(n_539),
    .Y(n_551));
 AOI221xp5_ASAP7_75t_R g36693 (.A1(n_541),
    .A2(u4_fract_out[5]),
    .B1(n_2),
    .B2(n_3782),
    .C(n_3),
    .Y(n_550));
 AOI221xp5_ASAP7_75t_R g36694 (.A1(n_541),
    .A2(u4_fract_out[3]),
    .B1(n_538),
    .B2(n_3780),
    .C(n_539),
    .Y(n_549));
 AOI221xp5_ASAP7_75t_R g36695 (.A1(n_541),
    .A2(u4_fract_out[16]),
    .B1(n_538),
    .B2(n_3793),
    .C(n_539),
    .Y(n_548));
 AOI221xp5_ASAP7_75t_R g36696 (.A1(n_541),
    .A2(u4_fract_out[12]),
    .B1(n_538),
    .B2(n_3789),
    .C(n_539),
    .Y(n_547));
 AOI221xp5_ASAP7_75t_R g36697 (.A1(n_541),
    .A2(u4_fract_out[4]),
    .B1(n_538),
    .B2(n_3781),
    .C(n_539),
    .Y(n_546));
 AOI221xp5_ASAP7_75t_R g36698 (.A1(n_5),
    .A2(u4_fract_out[21]),
    .B1(n_538),
    .B2(n_3798),
    .C(n_3),
    .Y(n_545));
 AOI221xp5_ASAP7_75t_R g36699 (.A1(n_541),
    .A2(u4_g),
    .B1(n_2),
    .B2(n_39),
    .C(n_3),
    .Y(n_543));
 AOI22xp33_ASAP7_75t_R g36700 (.A1(u4_fract_out[7]),
    .A2(n_541),
    .B1(n_3784),
    .B2(n_538),
    .Y(n_542));
 AOI21xp33_ASAP7_75t_R g36703 (.A1(n_250),
    .A2(n_117),
    .B(n_537),
    .Y(n_540));
 AND2x2_ASAP7_75t_R g36704 (.A(n_534),
    .B(n_14),
    .Y(n_541));
 AOI31xp33_ASAP7_75t_R g36709 (.A1(n_498),
    .A2(n_450),
    .A3(n_3513),
    .B(n_535),
    .Y(n_539));
 O2A1O1Ixp33_ASAP7_75t_R g36710 (.A1(n_3756),
    .A2(n_245),
    .B(n_106),
    .C(n_535),
    .Y(n_538));
 O2A1O1Ixp33_ASAP7_75t_R g36711 (.A1(n_275),
    .A2(n_360),
    .B(n_532),
    .C(n_315),
    .Y(n_536));
 OR3x1_ASAP7_75t_R g36712 (.A(n_533),
    .B(n_532),
    .C(n_509),
    .Y(n_537));
 INVxp33_ASAP7_75t_R g36713 (.A(n_534),
    .Y(n_535));
 AOI311xp33_ASAP7_75t_R g36714 (.A1(n_530),
    .A2(n_3803),
    .A3(n_118),
    .B(n_289),
    .C(n_501),
    .Y(n_534));
 OAI32xp33_ASAP7_75t_R g36715 (.A1(n_530),
    .A2(n_511),
    .A3(n_13919),
    .B1(n_3850),
    .B2(n_294),
    .Y(n_533));
 OAI322xp33_ASAP7_75t_R g36716 (.A1(n_529),
    .A2(n_132),
    .A3(n_117),
    .B1(n_510),
    .B2(n_13919),
    .C1(n_401),
    .C2(n_22),
    .Y(n_532));
 NOR5xp2_ASAP7_75t_R g36717 (.A(n_527),
    .B(n_514),
    .C(n_513),
    .D(n_518),
    .E(n_515),
    .Y(n_531));
 INVxp33_ASAP7_75t_R g36718 (.A(n_529),
    .Y(n_530));
 NAND5xp2_ASAP7_75t_R g36719 (.A(n_528),
    .B(n_513),
    .C(n_519),
    .D(n_514),
    .E(n_508),
    .Y(n_529));
 AND4x1_ASAP7_75t_R g36720 (.A(n_515),
    .B(n_517),
    .C(n_512),
    .D(n_518),
    .Y(n_528));
 OR4x1_ASAP7_75t_R g36721 (.A(n_517),
    .B(n_512),
    .C(n_519),
    .D(n_508),
    .Y(n_527));
 NOR2xp33_ASAP7_75t_R g36729 (.A(n_8),
    .B(n_519),
    .Y(n_526));
 NOR2xp33_ASAP7_75t_R g36730 (.A(n_381),
    .B(n_518),
    .Y(n_525));
 NOR2xp33_ASAP7_75t_R g36732 (.A(n_381),
    .B(n_514),
    .Y(n_524));
 NOR2xp33_ASAP7_75t_R g36733 (.A(n_8),
    .B(n_512),
    .Y(n_523));
 NOR2xp33_ASAP7_75t_R g36734 (.A(n_381),
    .B(n_513),
    .Y(n_522));
 NOR2xp33_ASAP7_75t_R g36735 (.A(n_8),
    .B(n_515),
    .Y(n_521));
 NOR2xp33_ASAP7_75t_R g36736 (.A(n_8),
    .B(n_517),
    .Y(n_520));
 NOR2xp33_ASAP7_75t_R g36737 (.A(n_381),
    .B(n_508),
    .Y(n_516));
 A2O1A1Ixp33_ASAP7_75t_R g36738 (.A1(n_435),
    .A2(n_478),
    .B(n_502),
    .C(n_507),
    .Y(n_519));
 OAI21xp33_ASAP7_75t_R g36739 (.A1(n_491),
    .A2(n_502),
    .B(n_507),
    .Y(n_518));
 A2O1A1Ixp33_ASAP7_75t_R g36740 (.A1(n_435),
    .A2(n_487),
    .B(n_502),
    .C(n_507),
    .Y(n_517));
 OAI21xp33_ASAP7_75t_R g36741 (.A1(n_492),
    .A2(n_502),
    .B(n_507),
    .Y(n_515));
 OAI21xp33_ASAP7_75t_R g36742 (.A1(n_490),
    .A2(n_502),
    .B(n_507),
    .Y(n_514));
 OAI21xp33_ASAP7_75t_R g36743 (.A1(n_485),
    .A2(n_502),
    .B(n_507),
    .Y(n_513));
 OAI21xp33_ASAP7_75t_R g36744 (.A1(n_480),
    .A2(n_502),
    .B(n_507),
    .Y(n_512));
 NAND3xp33_ASAP7_75t_R g36745 (.A(n_505),
    .B(n_474),
    .C(n_123),
    .Y(n_511));
 OA211x2_ASAP7_75t_R g36746 (.A1(n_204),
    .A2(n_401),
    .B(n_505),
    .C(n_123),
    .Y(n_510));
 OAI221xp5_ASAP7_75t_R g36747 (.A1(n_38),
    .A2(n_3594),
    .B1(n_302),
    .B2(n_3803),
    .C(n_503),
    .Y(n_509));
 OAI22xp33_ASAP7_75t_R g36748 (.A1(n_305),
    .A2(n_506),
    .B1(n_475),
    .B2(n_502),
    .Y(n_508));
 OAI21xp33_ASAP7_75t_R g36749 (.A1(n_292),
    .A2(n_504),
    .B(n_304),
    .Y(n_507));
 NOR2xp33_ASAP7_75t_R g36750 (.A(n_292),
    .B(n_501),
    .Y(n_506));
 INVxp33_ASAP7_75t_R g36751 (.A(n_504),
    .Y(n_505));
 NAND2xp33_ASAP7_75t_R g36752 (.A(n_3497),
    .B(n_499),
    .Y(n_503));
 NAND2xp33_ASAP7_75t_R g36753 (.A(n_498),
    .B(n_500),
    .Y(n_504));
 NAND2xp33_ASAP7_75t_R g36754 (.A(n_304),
    .B(n_498),
    .Y(n_502));
 INVxp33_ASAP7_75t_R g36755 (.A(n_500),
    .Y(n_501));
 NAND3xp33_ASAP7_75t_R g36756 (.A(n_498),
    .B(n_109),
    .C(n_3555),
    .Y(n_499));
 AOI331xp33_ASAP7_75t_R g36757 (.A1(n_358),
    .A2(n_22),
    .A3(n_67),
    .B1(n_496),
    .B2(u4_op_dn),
    .B3(rmode_r3[1]),
    .C1(n_445),
    .Y(n_500));
 AOI32xp33_ASAP7_75t_R g36758 (.A1(n_347),
    .A2(n_3801),
    .A3(n_3756),
    .B1(n_497),
    .B2(n_22),
    .Y(n_498));
 OAI221xp5_ASAP7_75t_R g36759 (.A1(n_414),
    .A2(exp_ovf_r[1]),
    .B1(n_357),
    .B2(n_118),
    .C(n_495),
    .Y(n_497));
 NOR5xp2_ASAP7_75t_R g36760 (.A(n_494),
    .B(n_3573),
    .C(n_3508),
    .D(n_13920),
    .E(sign),
    .Y(n_496));
 A2O1A1Ixp33_ASAP7_75t_R g36761 (.A1(n_137),
    .A2(n_493),
    .B(n_403),
    .C(sign),
    .Y(n_495));
 NOR4xp25_ASAP7_75t_R g36762 (.A(n_492),
    .B(n_489),
    .C(n_491),
    .D(n_490),
    .Y(n_494));
 OAI321xp33_ASAP7_75t_R g36763 (.A1(n_417),
    .A2(n_3502),
    .A3(n_3508),
    .B1(n_24),
    .B2(n_13845),
    .C(n_398),
    .Y(n_493));
 AND5x1_ASAP7_75t_R g36764 (.A(n_471),
    .B(n_429),
    .C(n_376),
    .D(n_356),
    .E(n_435),
    .Y(n_492));
 AOI211xp5_ASAP7_75t_R g36766 (.A1(n_353),
    .A2(n_3762),
    .B(n_481),
    .C(n_436),
    .Y(n_491));
 NAND3xp33_ASAP7_75t_R g36767 (.A(n_484),
    .B(n_479),
    .C(n_475),
    .Y(n_489));
 AOI211xp5_ASAP7_75t_R g36769 (.A1(n_353),
    .A2(n_3761),
    .B(n_483),
    .C(n_436),
    .Y(n_490));
 AND4x1_ASAP7_75t_R g36770 (.A(n_467),
    .B(n_380),
    .C(n_356),
    .D(n_402),
    .Y(n_487));
 AOI211xp5_ASAP7_75t_R g36771 (.A1(u1_n_852),
    .A2(n_143),
    .B(n_477),
    .C(n_419),
    .Y(n_486));
 INVxp33_ASAP7_75t_R g36772 (.A(n_484),
    .Y(n_485));
 NAND2xp33_ASAP7_75t_R g36773 (.A(n_325),
    .B(n_476),
    .Y(n_483));
 OAI211xp5_ASAP7_75t_R g36774 (.A1(n_3805),
    .A2(n_354),
    .B(n_469),
    .C(n_435),
    .Y(n_484));
 A2O1A1Ixp33_ASAP7_75t_R g36776 (.A1(n_270),
    .A2(n_3776),
    .B(n_356),
    .C(n_472),
    .Y(n_481));
 INVxp33_ASAP7_75t_R g36777 (.A(n_479),
    .Y(n_480));
 OAI221xp5_ASAP7_75t_R g36778 (.A1(n_99),
    .A2(u1_n_1593),
    .B1(n_378),
    .B2(u1_n_5054),
    .C(n_464),
    .Y(n_477));
 AOI221xp5_ASAP7_75t_R g36779 (.A1(n_352),
    .A2(n_263),
    .B1(n_415),
    .B2(exp_r[3]),
    .C(n_468),
    .Y(n_476));
 NAND3xp33_ASAP7_75t_R g36780 (.A(n_422),
    .B(n_462),
    .C(n_435),
    .Y(n_479));
 AOI221xp5_ASAP7_75t_R g36781 (.A1(n_353),
    .A2(n_3765),
    .B1(n_457),
    .B2(u4_exp_out[7]),
    .C(n_439),
    .Y(n_478));
 OAI332xp33_ASAP7_75t_R g36782 (.A1(n_456),
    .A2(exp_ovf_r[1]),
    .A3(exp_ovf_r[0]),
    .B1(n_38),
    .B2(n_104),
    .B3(opb_dn),
    .C1(n_421),
    .C2(n_3496),
    .Y(n_474));
 OR5x1_ASAP7_75t_R g36783 (.A(n_465),
    .B(prod[26]),
    .C(prod[1]),
    .D(prod[25]),
    .E(prod[2]),
    .Y(n_473));
 AOI221xp5_ASAP7_75t_R g36784 (.A1(n_461),
    .A2(n_3724),
    .B1(n_415),
    .B2(exp_r[4]),
    .C(n_392),
    .Y(n_472));
 AOI22xp33_ASAP7_75t_R g36785 (.A1(n_3725),
    .A2(n_466),
    .B1(n_269),
    .B2(n_344),
    .Y(n_471));
 AOI21xp33_ASAP7_75t_R g36786 (.A1(n_415),
    .A2(n_13972),
    .B(n_470),
    .Y(n_475));
 OAI21xp33_ASAP7_75t_R g36787 (.A1(n_3727),
    .A2(n_354),
    .B(n_463),
    .Y(n_470));
 AOI211xp5_ASAP7_75t_R g36788 (.A1(n_458),
    .A2(n_3722),
    .B(n_430),
    .C(n_388),
    .Y(n_469));
 OAI22xp33_ASAP7_75t_R g36789 (.A1(n_37),
    .A2(n_459),
    .B1(n_3767),
    .B2(n_356),
    .Y(n_468));
 AOI221xp5_ASAP7_75t_R g36790 (.A1(n_460),
    .A2(n_3726),
    .B1(n_415),
    .B2(exp_r[6]),
    .C(n_391),
    .Y(n_467));
 AO221x1_ASAP7_75t_R g36791 (.A1(n_352),
    .A2(n_324),
    .B1(n_3724),
    .B2(n_269),
    .C(n_461),
    .Y(n_466));
 NAND4xp25_ASAP7_75t_R g36792 (.A(n_451),
    .B(n_332),
    .C(n_164),
    .D(n_201),
    .Y(n_465));
 AOI21xp33_ASAP7_75t_R g36793 (.A1(n_454),
    .A2(u1_n_2218),
    .B(n_412),
    .Y(n_464));
 AOI221xp5_ASAP7_75t_R g36794 (.A1(n_452),
    .A2(u4_exp_out[0]),
    .B1(n_355),
    .B2(n_337),
    .C(n_393),
    .Y(n_463));
 AOI22xp33_ASAP7_75t_R g36795 (.A1(n_452),
    .A2(n_3721),
    .B1(n_415),
    .B2(exp_r[1]),
    .Y(n_462));
 OAI221xp5_ASAP7_75t_R g36796 (.A1(n_351),
    .A2(n_362),
    .B1(n_344),
    .B2(n_268),
    .C(n_453),
    .Y(n_460));
 AOI221xp5_ASAP7_75t_R g36797 (.A1(n_352),
    .A2(n_242),
    .B1(n_241),
    .B2(n_269),
    .C(n_452),
    .Y(n_459));
 OAI21xp33_ASAP7_75t_R g36798 (.A1(n_268),
    .A2(n_277),
    .B(n_453),
    .Y(n_461));
 OAI221xp5_ASAP7_75t_R g36799 (.A1(n_351),
    .A2(n_126),
    .B1(n_138),
    .B2(n_268),
    .C(n_453),
    .Y(n_458));
 OAI221xp5_ASAP7_75t_R g36800 (.A1(n_351),
    .A2(n_382),
    .B1(n_384),
    .B2(n_268),
    .C(n_453),
    .Y(n_457));
 AOI21xp33_ASAP7_75t_R g36801 (.A1(n_36),
    .A2(n_3556),
    .B(n_455),
    .Y(n_456));
 AOI21xp33_ASAP7_75t_R g36802 (.A1(n_440),
    .A2(n_329),
    .B(u4_n_1722),
    .Y(n_455));
 NAND4xp25_ASAP7_75t_R g36803 (.A(n_432),
    .B(n_14279),
    .C(n_291),
    .D(n_14278),
    .Y(n_454));
 INVxp33_ASAP7_75t_R g36804 (.A(n_453),
    .Y(n_452));
 NOR5xp2_ASAP7_75t_R g36805 (.A(n_428),
    .B(n_163),
    .C(prod[42]),
    .D(prod[0]),
    .E(prod[36]),
    .Y(n_451));
 AOI332xp33_ASAP7_75t_R g36806 (.A1(n_288),
    .A2(n_411),
    .A3(n_117),
    .B1(n_427),
    .B2(n_3579),
    .B3(rmode_r3[1]),
    .C1(n_287),
    .C2(n_67),
    .Y(n_453));
 AOI22xp33_ASAP7_75t_R g36816 (.A1(n_131),
    .A2(n_415),
    .B1(n_13919),
    .B2(n_436),
    .Y(n_450));
 NAND2xp33_ASAP7_75t_R g36817 (.A(u1_exp_large[3]),
    .B(n_437),
    .Y(n_449));
 NAND2xp33_ASAP7_75t_R g36820 (.A(u1_exp_large[0]),
    .B(n_437),
    .Y(n_448));
 NAND2xp33_ASAP7_75t_R g36821 (.A(u1_exp_large[1]),
    .B(n_437),
    .Y(n_447));
 NAND2xp33_ASAP7_75t_R g36822 (.A(u1_exp_large[2]),
    .B(n_437),
    .Y(n_446));
 O2A1O1Ixp33_ASAP7_75t_R g36824 (.A1(n_66),
    .A2(n_317),
    .B(n_423),
    .C(sign),
    .Y(n_445));
 NAND2xp33_ASAP7_75t_R g36825 (.A(u1_exp_large[5]),
    .B(n_437),
    .Y(n_444));
 NAND2xp33_ASAP7_75t_R g36826 (.A(u1_exp_large[6]),
    .B(n_437),
    .Y(n_443));
 NAND2xp33_ASAP7_75t_R g36827 (.A(u1_exp_large[7]),
    .B(n_437),
    .Y(n_442));
 NAND2xp33_ASAP7_75t_R g36828 (.A(u1_exp_large[4]),
    .B(n_437),
    .Y(n_441));
 NAND5xp2_ASAP7_75t_R g36829 (.A(n_399),
    .B(n_3524),
    .C(n_50),
    .D(n_43),
    .E(n_3556),
    .Y(n_440));
 OAI221xp5_ASAP7_75t_R g36830 (.A1(n_407),
    .A2(u4_exp_out[7]),
    .B1(n_414),
    .B2(n_24),
    .C(n_356),
    .Y(n_439));
 AOI211xp5_ASAP7_75t_R g36831 (.A1(n_120),
    .A2(n_334),
    .B(n_418),
    .C(n_370),
    .Y(n_438));
 INVxp33_ASAP7_75t_R g36832 (.A(n_436),
    .Y(n_435));
 OA211x2_ASAP7_75t_R g36835 (.A1(u2_exp_tmp1[5]),
    .A2(n_394),
    .B(n_409),
    .C(n_373),
    .Y(n_434));
 NAND5xp2_ASAP7_75t_R g36836 (.A(n_205),
    .B(n_371),
    .C(n_157),
    .D(n_156),
    .E(n_103),
    .Y(n_437));
 NOR2xp33_ASAP7_75t_R g36837 (.A(n_66),
    .B(n_427),
    .Y(n_436));
 AOI211xp5_ASAP7_75t_R g36838 (.A1(n_228),
    .A2(n_260),
    .B(n_410),
    .C(n_348),
    .Y(n_433));
 NOR3xp33_ASAP7_75t_R g36839 (.A(n_406),
    .B(u1_n_917),
    .C(u1_n_923),
    .Y(n_432));
 AOI21xp33_ASAP7_75t_R g36840 (.A1(n_365),
    .A2(n_199),
    .B(n_420),
    .Y(n_431));
 AO32x1_ASAP7_75t_R g36841 (.A1(n_352),
    .A2(n_126),
    .A3(n_40),
    .B1(n_415),
    .B2(exp_r[2]),
    .Y(n_430));
 AOI22xp33_ASAP7_75t_R g36842 (.A1(n_350),
    .A2(n_352),
    .B1(exp_r[5]),
    .B2(n_415),
    .Y(n_429));
 OR5x1_ASAP7_75t_R g36843 (.A(n_405),
    .B(prod[46]),
    .C(prod[38]),
    .D(prod[45]),
    .E(prod[39]),
    .Y(n_428));
 A2O1A1O1Ixp25_ASAP7_75t_R g36844 (.A1(u2_n_1398),
    .A2(n_127),
    .B(n_225),
    .C(n_120),
    .D(n_404),
    .Y(n_426));
 AO21x1_ASAP7_75t_R g36845 (.A1(n_3487),
    .A2(n_326),
    .B(n_417),
    .Y(n_425));
 AOI221xp5_ASAP7_75t_R g36846 (.A1(n_312),
    .A2(n_33),
    .B1(n_280),
    .B2(n_243),
    .C(n_408),
    .Y(n_424));
 A2O1A1Ixp33_ASAP7_75t_R g36847 (.A1(n_68),
    .A2(n_386),
    .B(n_403),
    .C(n_22),
    .Y(n_423));
 NAND2xp33_ASAP7_75t_R g36848 (.A(n_3803),
    .B(n_416),
    .Y(n_427));
 AOI221xp5_ASAP7_75t_R g36849 (.A1(n_244),
    .A2(n_269),
    .B1(n_353),
    .B2(n_3808),
    .C(n_387),
    .Y(n_422));
 OA332x1_ASAP7_75t_R g36850 (.A1(n_342),
    .A2(n_112),
    .A3(u4_op_dn),
    .B1(n_160),
    .B2(n_3502),
    .B3(u4_op_dn),
    .C1(n_329),
    .C2(n_369),
    .Y(n_421));
 OAI31xp33_ASAP7_75t_R g36851 (.A1(n_115),
    .A2(n_199),
    .A3(n_14296),
    .B(n_413),
    .Y(n_420));
 AO32x1_ASAP7_75t_R g36852 (.A1(n_377),
    .A2(u1_n_850),
    .A3(u1_n_840),
    .B1(u1_n_969),
    .B2(n_94),
    .Y(n_419));
 OAI221xp5_ASAP7_75t_R g36853 (.A1(n_251),
    .A2(n_331),
    .B1(n_375),
    .B2(u2_exp_tmp1[6]),
    .C(n_341),
    .Y(n_418));
 INVxp33_ASAP7_75t_R g36854 (.A(n_417),
    .Y(n_416));
 INVxp33_ASAP7_75t_R g36855 (.A(n_415),
    .Y(n_414));
 A2O1A1Ixp33_ASAP7_75t_R g36856 (.A1(u2_exp_tmp1[6]),
    .A2(n_228),
    .B(n_374),
    .C(u2_exp_tmp1[7]),
    .Y(n_413));
 O2A1O1Ixp33_ASAP7_75t_R g36859 (.A1(n_27),
    .A2(n_14279),
    .B(n_310),
    .C(u1_n_4993),
    .Y(n_412));
 NAND2xp33_ASAP7_75t_R g36860 (.A(n_3803),
    .B(n_400),
    .Y(n_411));
 NAND2xp33_ASAP7_75t_R g36861 (.A(sign),
    .B(n_400),
    .Y(n_417));
 NOR2xp33_ASAP7_75t_R g36862 (.A(n_118),
    .B(n_401),
    .Y(n_415));
 OAI22xp33_ASAP7_75t_R g36863 (.A1(n_14295),
    .A2(n_368),
    .B1(n_267),
    .B2(n_119),
    .Y(n_410));
 AOI22xp33_ASAP7_75t_R g36864 (.A1(n_335),
    .A2(n_120),
    .B1(u2_exp_tmp1[5]),
    .B2(n_364),
    .Y(n_409));
 OAI221xp5_ASAP7_75t_R g36865 (.A1(n_119),
    .A2(n_303),
    .B1(u2_n_772),
    .B2(n_339),
    .C(n_340),
    .Y(n_408));
 OA21x2_ASAP7_75t_R g36866 (.A1(n_383),
    .A2(n_351),
    .B(n_402),
    .Y(n_407));
 OAI221xp5_ASAP7_75t_R g36867 (.A1(n_320),
    .A2(n_51),
    .B1(n_27),
    .B2(n_14277),
    .C(n_396),
    .Y(n_406));
 OR5x1_ASAP7_75t_R g36868 (.A(n_298),
    .B(n_161),
    .C(prod[47]),
    .D(prod[17]),
    .E(prod[8]),
    .Y(n_405));
 OAI21xp33_ASAP7_75t_R g36869 (.A1(n_240),
    .A2(u2_n_772),
    .B(n_389),
    .Y(n_404));
 INVxp33_ASAP7_75t_R g36870 (.A(n_401),
    .Y(n_400));
 NOR4xp25_ASAP7_75t_R g36871 (.A(n_3734),
    .B(n_319),
    .C(exp_r[2]),
    .D(exp_r[1]),
    .Y(n_399));
 A2O1A1Ixp33_ASAP7_75t_R g36872 (.A1(exp_ovf_r[0]),
    .A2(n_32),
    .B(n_358),
    .C(fract_denorm[47]),
    .Y(n_398));
 OR2x2_ASAP7_75t_R g36873 (.A(fpu_op_r3[2]),
    .B(n_385),
    .Y(n_397));
 A2O1A1O1Ixp25_ASAP7_75t_R g36874 (.A1(u1_n_852),
    .A2(n_285),
    .B(n_14297),
    .C(u1_n_840),
    .D(u1_n_921),
    .Y(n_396));
 AND2x2_ASAP7_75t_R g36875 (.A(n_36),
    .B(n_386),
    .Y(n_403));
 NOR2xp33_ASAP7_75t_R g36876 (.A(n_385),
    .B(n_13),
    .Y(n_395));
 NAND2xp33_ASAP7_75t_R g36877 (.A(n_384),
    .B(n_269),
    .Y(n_402));
 NAND2xp33_ASAP7_75t_R g36878 (.A(u4_exp_out[7]),
    .B(n_382),
    .Y(n_401));
 AOI211xp5_ASAP7_75t_R g36879 (.A1(n_25),
    .A2(n_322),
    .B(n_312),
    .C(n_280),
    .Y(n_394));
 AOI21xp33_ASAP7_75t_R g36880 (.A1(n_268),
    .A2(n_351),
    .B(u4_exp_out[0]),
    .Y(n_393));
 OAI22xp33_ASAP7_75t_R g36881 (.A1(n_336),
    .A2(n_351),
    .B1(n_3724),
    .B2(n_325),
    .Y(n_392));
 NOR3xp33_ASAP7_75t_R g36882 (.A(n_351),
    .B(n_361),
    .C(n_3726),
    .Y(n_391));
 AOI211xp5_ASAP7_75t_R g36883 (.A1(n_228),
    .A2(n_159),
    .B(n_366),
    .C(n_221),
    .Y(n_390));
 AOI221xp5_ASAP7_75t_R g36884 (.A1(n_116),
    .A2(n_266),
    .B1(n_286),
    .B2(n_122),
    .C(n_372),
    .Y(n_389));
 A2O1A1Ixp33_ASAP7_75t_R g36885 (.A1(n_3770),
    .A2(n_270),
    .B(n_356),
    .C(n_313),
    .Y(n_388));
 OAI22xp33_ASAP7_75t_R g36886 (.A1(n_356),
    .A2(n_13847),
    .B1(n_351),
    .B2(n_244),
    .Y(n_387));
 INVxp33_ASAP7_75t_R g36887 (.A(n_383),
    .Y(n_382));
 INVxp33_ASAP7_75t_R g36891 (.A(n_13),
    .Y(n_381));
 NAND2xp33_ASAP7_75t_R g36892 (.A(n_3764),
    .B(n_353),
    .Y(n_380));
 OAI21xp33_ASAP7_75t_R g36893 (.A1(sign_mul_r),
    .A2(n_130),
    .B(n_345),
    .Y(n_379));
 AOI211xp5_ASAP7_75t_R g36894 (.A1(u1_n_852),
    .A2(n_283),
    .B(u1_n_996),
    .C(u1_n_990),
    .Y(n_378));
 NAND2xp33_ASAP7_75t_R g36895 (.A(n_14279),
    .B(n_291),
    .Y(n_377));
 NAND2xp33_ASAP7_75t_R g36896 (.A(n_3763),
    .B(n_353),
    .Y(n_376));
 AND2x2_ASAP7_75t_R g36898 (.A(n_137),
    .B(n_358),
    .Y(n_386));
 NOR3xp33_ASAP7_75t_R g36899 (.A(n_299),
    .B(n_148),
    .C(n_113),
    .Y(n_385));
 NOR2xp33_ASAP7_75t_R g36900 (.A(n_3726),
    .B(n_343),
    .Y(n_384));
 NAND2xp33_ASAP7_75t_R g36901 (.A(n_3726),
    .B(n_362),
    .Y(n_383));
 OAI31xp33_ASAP7_75t_R g36902 (.A1(n_254),
    .A2(n_284),
    .A3(n_113),
    .B(n_3594),
    .Y(n_13));
 INVxp33_ASAP7_75t_R g36903 (.A(n_374),
    .Y(n_375));
 A2O1A1Ixp33_ASAP7_75t_R g36904 (.A1(n_290),
    .A2(n_234),
    .B(n_314),
    .C(n_116),
    .Y(n_373));
 O2A1O1Ixp33_ASAP7_75t_R g36905 (.A1(n_139),
    .A2(u2_n_772),
    .B(n_307),
    .C(u2_exp_tmp1[2]),
    .Y(n_372));
 NOR4xp25_ASAP7_75t_R g36906 (.A(u1_n_590),
    .B(n_293),
    .C(n_155),
    .D(n_165),
    .Y(n_371));
 NOR3xp33_ASAP7_75t_R g36907 (.A(u2_n_772),
    .B(u2_exp_tmp1[6]),
    .C(n_318),
    .Y(n_370));
 O2A1O1Ixp33_ASAP7_75t_R g36908 (.A1(exp_r[7]),
    .A2(n_256),
    .B(n_3501),
    .C(n_3556),
    .Y(n_369));
 AOI211xp5_ASAP7_75t_R g36909 (.A1(n_25),
    .A2(n_240),
    .B(n_306),
    .C(n_286),
    .Y(n_368));
 A2O1A1Ixp33_ASAP7_75t_R g36910 (.A1(sign_mul_r),
    .A2(n_282),
    .B(n_316),
    .C(n_230),
    .Y(n_367));
 OAI321xp33_ASAP7_75t_R g36911 (.A1(n_115),
    .A2(n_147),
    .A3(u2_exp_tmp1[0]),
    .B1(n_220),
    .B2(u2_n_772),
    .C(n_301),
    .Y(n_366));
 OAI32xp33_ASAP7_75t_R g36912 (.A1(n_119),
    .A2(n_273),
    .A3(n_134),
    .B1(n_309),
    .B2(n_115),
    .Y(n_365));
 OAI22xp33_ASAP7_75t_R g36913 (.A1(n_279),
    .A2(n_229),
    .B1(n_322),
    .B2(u2_n_772),
    .Y(n_364));
 OAI21xp33_ASAP7_75t_R g36914 (.A1(n_330),
    .A2(n_229),
    .B(n_125),
    .Y(n_374));
 INVxp33_ASAP7_75t_R g36915 (.A(n_361),
    .Y(n_362));
 INVxp33_ASAP7_75t_R g36916 (.A(n_358),
    .Y(n_357));
 INVxp33_ASAP7_75t_R g36917 (.A(n_356),
    .Y(n_355));
 INVxp33_ASAP7_75t_R g36918 (.A(n_354),
    .Y(n_353));
 INVxp33_ASAP7_75t_R g36919 (.A(n_352),
    .Y(n_351));
 NOR2xp33_ASAP7_75t_R g36921 (.A(n_3725),
    .B(n_324),
    .Y(n_350));
 AOI211xp5_ASAP7_75t_R g36922 (.A1(u1_n_909),
    .A2(u1_n_2218),
    .B(n_158),
    .C(n_300),
    .Y(n_349));
 OAI22xp33_ASAP7_75t_R g36923 (.A1(n_265),
    .A2(n_115),
    .B1(n_272),
    .B2(u2_n_772),
    .Y(n_348));
 OAI31xp33_ASAP7_75t_R g36924 (.A1(n_206),
    .A2(exp_ovf_r[1]),
    .A3(exp_ovf_r[0]),
    .B(n_123),
    .Y(n_347));
 A2O1A1Ixp33_ASAP7_75t_R g36925 (.A1(n_145),
    .A2(n_23),
    .B(n_284),
    .C(n_198),
    .Y(n_363));
 NAND2xp33_ASAP7_75t_R g36926 (.A(n_323),
    .B(n_3725),
    .Y(n_361));
 O2A1O1Ixp33_ASAP7_75t_R g36927 (.A1(n_113),
    .A2(n_3498),
    .B(n_281),
    .C(inf_d),
    .Y(n_360));
 NOR3xp33_ASAP7_75t_R g36929 (.A(n_327),
    .B(n_3804),
    .C(n_3527),
    .Y(n_358));
 NAND2xp33_ASAP7_75t_R g36930 (.A(n_22),
    .B(n_328),
    .Y(n_356));
 NAND2xp33_ASAP7_75t_R g36931 (.A(n_13919),
    .B(n_328),
    .Y(n_354));
 OAI22xp33_ASAP7_75t_R g36932 (.A1(n_3756),
    .A2(n_287),
    .B1(n_202),
    .B2(n_3579),
    .Y(n_352));
 INVxp33_ASAP7_75t_R g36934 (.A(n_344),
    .Y(n_343));
 A2O1A1Ixp33_ASAP7_75t_R g36935 (.A1(n_24),
    .A2(n_248),
    .B(n_3556),
    .C(n_297),
    .Y(n_342));
 A2O1A1Ixp33_ASAP7_75t_R g36936 (.A1(u2_n_140),
    .A2(n_237),
    .B(n_262),
    .C(n_116),
    .Y(n_341));
 A2O1A1Ixp33_ASAP7_75t_R g36937 (.A1(u2_n_1384),
    .A2(n_238),
    .B(n_264),
    .C(n_116),
    .Y(n_340));
 AOI21xp33_ASAP7_75t_R g36938 (.A1(n_272),
    .A2(n_33),
    .B(n_321),
    .Y(n_339));
 XOR2xp5_ASAP7_75t_R g36940 (.A(n_3595),
    .B(n_271),
    .Y(n_337));
 XOR2xp5_ASAP7_75t_R g36941 (.A(n_278),
    .B(n_3724),
    .Y(n_336));
 XNOR2xp5_ASAP7_75t_R g36942 (.A(n_234),
    .B(n_252),
    .Y(n_335));
 XOR2xp5_ASAP7_75t_R g36943 (.A(n_237),
    .B(n_273),
    .Y(n_334));
 OAI22xp33_ASAP7_75t_R g36944 (.A1(n_250),
    .A2(n_231),
    .B1(opb_inf),
    .B2(n_281),
    .Y(n_333));
 NOR5xp2_ASAP7_75t_R g36945 (.A(n_255),
    .B(prod[31]),
    .C(prod[30]),
    .D(prod[32]),
    .E(prod[33]),
    .Y(n_332));
 NAND4xp25_ASAP7_75t_R g36946 (.A(n_236),
    .B(opa_inf),
    .C(opb_inf),
    .D(sign_exe_r),
    .Y(n_345));
 NOR3xp33_ASAP7_75t_R g36947 (.A(n_276),
    .B(n_3724),
    .C(n_3725),
    .Y(n_344));
 INVxp33_ASAP7_75t_R g36948 (.A(n_330),
    .Y(n_331));
 INVxp33_ASAP7_75t_R g36949 (.A(n_326),
    .Y(n_327));
 INVxp33_ASAP7_75t_R g36950 (.A(n_323),
    .Y(n_324));
 INVxp33_ASAP7_75t_R g36951 (.A(n_321),
    .Y(n_322));
 NOR4xp25_ASAP7_75t_R g36952 (.A(n_285),
    .B(n_207),
    .C(u1_n_873),
    .D(u1_n_867),
    .Y(n_320));
 OA21x2_ASAP7_75t_R g36953 (.A1(n_200),
    .A2(n_3738),
    .B(n_3735),
    .Y(n_319));
 NOR2xp33_ASAP7_75t_R g36955 (.A(n_272),
    .B(u2_n_1487),
    .Y(n_318));
 A2O1A1Ixp33_ASAP7_75t_R g36956 (.A1(n_13919),
    .A2(n_32),
    .B(n_203),
    .C(n_3801),
    .Y(n_317));
 NOR2xp33_ASAP7_75t_R g36957 (.A(sign_mul_r),
    .B(n_282),
    .Y(n_316));
 NOR2xp33_ASAP7_75t_R g36958 (.A(n_128),
    .B(n_274),
    .Y(n_315));
 NOR2xp33_ASAP7_75t_R g36959 (.A(n_290),
    .B(n_234),
    .Y(n_314));
 OR2x2_ASAP7_75t_R g36960 (.A(n_268),
    .B(n_241),
    .Y(n_313));
 NOR2xp33_ASAP7_75t_R g36961 (.A(n_279),
    .B(u2_exp_tmp1[5]),
    .Y(n_330));
 NAND2xp33_ASAP7_75t_R g36962 (.A(u4_op_dn),
    .B(n_270),
    .Y(n_329));
 NOR2xp33_ASAP7_75t_R g36963 (.A(n_118),
    .B(n_288),
    .Y(n_328));
 NAND5xp2_ASAP7_75t_R g36964 (.A(n_3809),
    .B(n_105),
    .C(n_3814),
    .D(n_3806),
    .E(n_3805),
    .Y(n_326));
 NAND2xp33_ASAP7_75t_R g36965 (.A(n_269),
    .B(n_277),
    .Y(n_325));
 NOR2xp33_ASAP7_75t_R g36966 (.A(n_28),
    .B(n_278),
    .Y(n_323));
 NOR2xp33_ASAP7_75t_R g36967 (.A(n_33),
    .B(n_272),
    .Y(n_321));
 INVxp33_ASAP7_75t_R g36969 (.A(n_14296),
    .Y(n_309));
 INVxp33_ASAP7_75t_R g36970 (.A(n_306),
    .Y(n_307));
 INVxp33_ASAP7_75t_R g36971 (.A(n_304),
    .Y(n_305));
 XNOR2xp5_ASAP7_75t_R g36972 (.A(n_238),
    .B(n_233),
    .Y(n_303));
 AOI311xp33_ASAP7_75t_R g36973 (.A1(u4_f2i_zero),
    .A2(n_24),
    .A3(n_3532),
    .B(n_63),
    .C(u4_n_1248),
    .Y(n_302));
 A2O1A1Ixp33_ASAP7_75t_R g36974 (.A1(u2_exp_tmp1[0]),
    .A2(n_116),
    .B(n_120),
    .C(n_147),
    .Y(n_301));
 OAI32xp33_ASAP7_75t_R g36975 (.A1(u1_n_1592),
    .A2(u1_n_852),
    .A3(n_142),
    .B1(u1_n_1593),
    .B2(n_3481),
    .Y(n_300));
 OAI22xp33_ASAP7_75t_R g36976 (.A1(n_3850),
    .A2(n_198),
    .B1(n_13919),
    .B2(n_129),
    .Y(n_299));
 OR5x1_ASAP7_75t_R g36977 (.A(n_257),
    .B(prod[12]),
    .C(prod[7]),
    .D(prod[13]),
    .E(prod[6]),
    .Y(n_298));
 NAND3xp33_ASAP7_75t_R g36978 (.A(n_247),
    .B(n_24),
    .C(u4_exp_div[7]),
    .Y(n_297));
 NOR3xp33_ASAP7_75t_R g36979 (.A(n_235),
    .B(n_130),
    .C(opa_inf),
    .Y(n_296));
 AOI221xp5_ASAP7_75t_R g36980 (.A1(n_57),
    .A2(u1_n_937),
    .B1(n_14268),
    .B2(u1_n_997),
    .C(n_261),
    .Y(n_295));
 AOI33xp33_ASAP7_75t_R g36981 (.A1(n_3573),
    .A2(n_102),
    .A3(u4_n_1248),
    .B1(n_3532),
    .B2(exp_ovf_r[1]),
    .B3(n_65),
    .Y(n_294));
 NAND3xp33_ASAP7_75t_R g36982 (.A(u1_n_5489),
    .B(n_211),
    .C(n_196),
    .Y(n_293));
 OAI21xp33_ASAP7_75t_R g36983 (.A1(n_243),
    .A2(n_229),
    .B(n_125),
    .Y(n_312));
 NOR3xp33_ASAP7_75t_R g36984 (.A(n_283),
    .B(u1_n_966),
    .C(u1_n_972),
    .Y(n_310));
 OAI21xp33_ASAP7_75t_R g36986 (.A1(n_122),
    .A2(n_229),
    .B(n_125),
    .Y(n_306));
 AOI31xp33_ASAP7_75t_R g36987 (.A1(n_22),
    .A2(n_68),
    .A3(exp_ovf_r[1]),
    .B(n_289),
    .Y(n_304));
 INVxp33_ASAP7_75t_R g37030 (.A(n_277),
    .Y(n_276));
 INVxp33_ASAP7_75t_R g37031 (.A(n_274),
    .Y(n_275));
 INVxp33_ASAP7_75t_R g37032 (.A(n_271),
    .Y(n_270));
 INVxp33_ASAP7_75t_R g37033 (.A(n_269),
    .Y(n_268));
 XNOR2xp5_ASAP7_75t_R g37038 (.A(n_124),
    .B(n_140),
    .Y(n_267));
 XNOR2xp5_ASAP7_75t_R g37039 (.A(n_127),
    .B(u2_n_1392),
    .Y(n_266));
 XOR2xp5_ASAP7_75t_R g37040 (.A(n_124),
    .B(n_101),
    .Y(n_265));
 NOR2xp33_ASAP7_75t_R g37041 (.A(u2_n_1384),
    .B(n_238),
    .Y(n_264));
 NOR2xp33_ASAP7_75t_R g37042 (.A(n_3723),
    .B(n_242),
    .Y(n_263));
 NOR2xp33_ASAP7_75t_R g37043 (.A(u2_n_140),
    .B(n_237),
    .Y(n_262));
 OAI221xp5_ASAP7_75t_R g37044 (.A1(n_97),
    .A2(u1_n_1593),
    .B1(n_58),
    .B2(u1_n_4917),
    .C(n_110),
    .Y(n_261));
 AND3x1_ASAP7_75t_R g37046 (.A(n_14295),
    .B(n_69),
    .C(n_122),
    .Y(n_260));
 NAND3xp33_ASAP7_75t_R g37047 (.A(n_150),
    .B(n_30),
    .C(opa_nan_r),
    .Y(n_259));
 O2A1O1Ixp33_ASAP7_75t_R g37048 (.A1(opb_inf),
    .A2(n_30),
    .B(n_151),
    .C(n_235),
    .Y(n_258));
 OR3x1_ASAP7_75t_R g37049 (.A(n_162),
    .B(prod[15]),
    .C(prod[14]),
    .Y(n_257));
 OR4x1_ASAP7_75t_R g37050 (.A(n_59),
    .B(exp_r[3]),
    .C(exp_r[6]),
    .D(exp_r[5]),
    .Y(n_256));
 OR5x1_ASAP7_75t_R g37051 (.A(prod[27]),
    .B(prod[20]),
    .C(prod[23]),
    .D(prod[21]),
    .E(prod[22]),
    .Y(n_255));
 OAI22xp33_ASAP7_75t_R g37052 (.A1(n_13920),
    .A2(n_108),
    .B1(n_132),
    .B2(n_35),
    .Y(n_254));
 NOR3xp33_ASAP7_75t_R g37053 (.A(n_231),
    .B(n_100),
    .C(inf_mul_r),
    .Y(n_253));
 NOR2xp33_ASAP7_75t_R g37054 (.A(n_233),
    .B(n_136),
    .Y(n_252));
 OAI31xp33_ASAP7_75t_R g37055 (.A1(n_13920),
    .A2(n_3756),
    .A3(n_26),
    .B(n_3513),
    .Y(n_292));
 AOI211xp5_ASAP7_75t_R g37056 (.A1(u1_n_852),
    .A2(n_154),
    .B(u1_n_941),
    .C(u1_n_947),
    .Y(n_291));
 OAI21xp33_ASAP7_75t_R g37057 (.A1(n_136),
    .A2(n_48),
    .B(u2_n_1444),
    .Y(n_290));
 OAI22xp33_ASAP7_75t_R g37058 (.A1(n_107),
    .A2(n_13919),
    .B1(n_149),
    .B2(n_3850),
    .Y(n_289));
 NAND4xp25_ASAP7_75t_R g37059 (.A(n_3559),
    .B(n_53),
    .C(u4_g),
    .D(n_32),
    .Y(n_288));
 NAND2xp33_ASAP7_75t_R g37060 (.A(u4_fract_out_pl1[23]),
    .B(n_246),
    .Y(n_287));
 NOR2xp33_ASAP7_75t_R g37061 (.A(n_69),
    .B(n_229),
    .Y(n_286));
 OR3x1_ASAP7_75t_R g37062 (.A(n_14297),
    .B(u1_n_886),
    .C(u1_n_880),
    .Y(n_285));
 NAND2xp33_ASAP7_75t_R g37063 (.A(n_228),
    .B(u2_exp_tmp1[6]),
    .Y(n_251));
 NOR3xp33_ASAP7_75t_R g37064 (.A(n_3850),
    .B(n_3756),
    .C(n_128),
    .Y(n_284));
 OR4x1_ASAP7_75t_R g37065 (.A(u1_n_996),
    .B(u1_n_990),
    .C(u1_n_978),
    .D(u1_n_984),
    .Y(n_283));
 NAND2xp33_ASAP7_75t_R g37066 (.A(sign_exe_r),
    .B(n_197),
    .Y(n_282));
 NAND2xp33_ASAP7_75t_R g37067 (.A(n_236),
    .B(n_34),
    .Y(n_281));
 NOR2xp33_ASAP7_75t_R g37068 (.A(n_33),
    .B(n_229),
    .Y(n_280));
 NAND2xp33_ASAP7_75t_R g37069 (.A(n_33),
    .B(n_243),
    .Y(n_279));
 OR2x2_ASAP7_75t_R g37070 (.A(n_37),
    .B(n_242),
    .Y(n_278));
 NOR2xp33_ASAP7_75t_R g37071 (.A(n_3723),
    .B(n_241),
    .Y(n_277));
 NAND2xp33_ASAP7_75t_R g37072 (.A(n_35),
    .B(n_230),
    .Y(n_274));
 NAND2xp33_ASAP7_75t_R g37073 (.A(n_232),
    .B(u2_n_1399),
    .Y(n_273));
 NAND2xp33_ASAP7_75t_R g37074 (.A(n_14295),
    .B(n_239),
    .Y(n_272));
 A2O1A1Ixp33_ASAP7_75t_R g37075 (.A1(n_98),
    .A2(n_3565),
    .B(n_3516),
    .C(n_3523),
    .Y(n_271));
 NOR4xp25_ASAP7_75t_R g37076 (.A(n_3579),
    .B(n_3850),
    .C(n_66),
    .D(n_26),
    .Y(n_269));
 INVxp33_ASAP7_75t_R g37077 (.A(n_247),
    .Y(n_248));
 INVxp33_ASAP7_75t_R g37078 (.A(n_245),
    .Y(n_246));
 INVxp33_ASAP7_75t_R g37079 (.A(n_240),
    .Y(n_239));
 INVxp33_ASAP7_75t_R g37080 (.A(n_236),
    .Y(n_235));
 INVxp33_ASAP7_75t_R g37081 (.A(n_233),
    .Y(n_232));
 INVxp33_ASAP7_75t_R g37082 (.A(n_231),
    .Y(n_230));
 INVxp33_ASAP7_75t_R g37083 (.A(n_229),
    .Y(n_228));
 AOI22xp33_ASAP7_75t_R g37084 (.A1(u1_n_1049),
    .A2(n_20),
    .B1(u1_n_1022),
    .B2(u1_n_1066),
    .Y(n_227));
 AOI22xp33_ASAP7_75t_R g37085 (.A1(u1_n_1050),
    .A2(n_9),
    .B1(u1_n_1023),
    .B2(n_10),
    .Y(n_226));
 NOR2xp33_ASAP7_75t_R g37086 (.A(u2_n_1398),
    .B(n_127),
    .Y(n_225));
 AOI22xp33_ASAP7_75t_R g37087 (.A1(u1_n_1051),
    .A2(n_1),
    .B1(u1_n_1024),
    .B2(n_10),
    .Y(n_224));
 AOI22xp33_ASAP7_75t_R g37088 (.A1(u1_n_1052),
    .A2(n_7),
    .B1(u1_n_1025),
    .B2(n_11),
    .Y(n_223));
 AOI22xp33_ASAP7_75t_R g37089 (.A1(u1_n_1053),
    .A2(n_20),
    .B1(u1_n_1026),
    .B2(n_11),
    .Y(n_222));
 NOR2xp33_ASAP7_75t_R g37090 (.A(u2_exp_tmp1[1]),
    .B(n_125),
    .Y(n_221));
 NOR2xp33_ASAP7_75t_R g37091 (.A(n_122),
    .B(n_139),
    .Y(n_220));
 AOI22xp33_ASAP7_75t_R g37092 (.A1(u1_n_1055),
    .A2(n_20),
    .B1(u1_n_1028),
    .B2(n_17),
    .Y(n_219));
 AOI22xp33_ASAP7_75t_R g37093 (.A1(u1_n_1057),
    .A2(n_7),
    .B1(u1_n_1030),
    .B2(n_11),
    .Y(n_218));
 AOI22xp33_ASAP7_75t_R g37094 (.A1(u1_n_1059),
    .A2(n_20),
    .B1(u1_n_1032),
    .B2(n_12),
    .Y(n_217));
 AOI22xp33_ASAP7_75t_R g37095 (.A1(u1_n_1060),
    .A2(n_7),
    .B1(u1_n_1033),
    .B2(n_11),
    .Y(n_216));
 AOI22xp33_ASAP7_75t_R g37096 (.A1(u1_n_1061),
    .A2(n_20),
    .B1(u1_n_1034),
    .B2(n_11),
    .Y(n_215));
 AOI22xp33_ASAP7_75t_R g37097 (.A1(u1_n_1054),
    .A2(n_20),
    .B1(u1_n_1027),
    .B2(n_10),
    .Y(n_214));
 AOI22xp33_ASAP7_75t_R g37098 (.A1(u1_n_1056),
    .A2(n_7),
    .B1(u1_n_1029),
    .B2(u1_n_1066),
    .Y(n_213));
 AOI22xp33_ASAP7_75t_R g37099 (.A1(u1_n_1015),
    .A2(n_20),
    .B1(u1_n_1042),
    .B2(n_17),
    .Y(n_212));
 OAI21xp33_ASAP7_75t_R g37100 (.A1(opb_r[23]),
    .A2(opa_r[23]),
    .B(u1_n_8071),
    .Y(n_211));
 AOI22xp33_ASAP7_75t_R g37101 (.A1(u1_n_1014),
    .A2(n_7),
    .B1(u1_n_1041),
    .B2(u1_n_1066),
    .Y(n_210));
 AOI22xp33_ASAP7_75t_R g37102 (.A1(u1_n_1058),
    .A2(n_20),
    .B1(u1_n_1031),
    .B2(n_12),
    .Y(n_209));
 AOI22xp33_ASAP7_75t_R g37103 (.A1(u1_n_1016),
    .A2(n_7),
    .B1(u1_n_1043),
    .B2(n_10),
    .Y(n_208));
 AOI21xp33_ASAP7_75t_R g37104 (.A1(n_1163),
    .A2(u1_n_68),
    .B(n_27),
    .Y(n_207));
 NAND3xp33_ASAP7_75t_R g37105 (.A(u4_n_1438),
    .B(n_32),
    .C(n_46),
    .Y(n_206));
 AOI21xp33_ASAP7_75t_R g37106 (.A1(n_44),
    .A2(opb_r[25]),
    .B(u1_n_4702),
    .Y(n_205));
 AOI21xp33_ASAP7_75t_R g37107 (.A1(exp_r[7]),
    .A2(u4_op_dn),
    .B(exp_ovf_r[0]),
    .Y(n_204));
 AOI21xp33_ASAP7_75t_R g37108 (.A1(n_24),
    .A2(n_3502),
    .B(n_123),
    .Y(n_203));
 AOI21xp33_ASAP7_75t_R g37109 (.A1(n_3850),
    .A2(rmode_r3[1]),
    .B(n_137),
    .Y(n_202));
 NOR3xp33_ASAP7_75t_R g37110 (.A(prod[37]),
    .B(prod[24]),
    .C(prod[3]),
    .Y(n_201));
 AND3x1_ASAP7_75t_R g37111 (.A(n_3739),
    .B(n_3741),
    .C(n_3742),
    .Y(n_200));
 NAND2xp33_ASAP7_75t_R g37112 (.A(n_128),
    .B(n_144),
    .Y(n_250));
 OAI21xp33_ASAP7_75t_R g37114 (.A1(exp_r[6]),
    .A2(n_61),
    .B(n_3504),
    .Y(n_247));
 OAI21xp33_ASAP7_75t_R g37115 (.A1(u4_g),
    .A2(n_3559),
    .B(n_53),
    .Y(n_245));
 OR2x2_ASAP7_75t_R g37116 (.A(n_126),
    .B(n_138),
    .Y(n_244));
 NOR3xp33_ASAP7_75t_R g37117 (.A(n_14295),
    .B(n_121),
    .C(u2_exp_tmp1[2]),
    .Y(n_243));
 NAND2xp33_ASAP7_75t_R g37118 (.A(n_3722),
    .B(n_126),
    .Y(n_242));
 NAND2xp33_ASAP7_75t_R g37119 (.A(n_40),
    .B(n_138),
    .Y(n_241));
 NAND2xp33_ASAP7_75t_R g37120 (.A(u2_exp_tmp1[2]),
    .B(n_139),
    .Y(n_240));
 NAND2xp33_ASAP7_75t_R g37121 (.A(u2_n_1444),
    .B(n_135),
    .Y(n_238));
 NAND2xp33_ASAP7_75t_R g37122 (.A(n_152),
    .B(n_133),
    .Y(n_237));
 NOR2xp33_ASAP7_75t_R g37123 (.A(n_113),
    .B(n_13920),
    .Y(n_236));
 OAI21xp33_ASAP7_75t_R g37124 (.A1(n_31),
    .A2(u2_exp_tmp1[5]),
    .B(u2_n_1792),
    .Y(n_234));
 NAND2xp33_ASAP7_75t_R g37125 (.A(u2_n_1489),
    .B(n_141),
    .Y(n_233));
 NAND2xp33_ASAP7_75t_R g37126 (.A(n_114),
    .B(n_23),
    .Y(n_231));
 NAND3xp33_ASAP7_75t_R g37127 (.A(u2_exp_ovf_d[1]),
    .B(u2_n_775),
    .C(n_31),
    .Y(n_229));
 INVxp33_ASAP7_75t_R g37128 (.A(n_198),
    .Y(n_197));
 XNOR2xp5_ASAP7_75t_R g37129 (.A(opa_r[29]),
    .B(opb_r[29]),
    .Y(n_196));
 AOI22xp33_ASAP7_75t_R g37130 (.A1(u1_n_1045),
    .A2(n_20),
    .B1(u1_n_1018),
    .B2(n_10),
    .Y(n_195));
 AOI22xp33_ASAP7_75t_R g37131 (.A1(u1_n_1044),
    .A2(n_7),
    .B1(u1_n_1017),
    .B2(n_10),
    .Y(n_194));
 AOI22xp33_ASAP7_75t_R g37132 (.A1(u1_n_1043),
    .A2(n_1),
    .B1(u1_n_1016),
    .B2(n_12),
    .Y(n_193));
 AOI22xp33_ASAP7_75t_R g37133 (.A1(u1_n_1042),
    .A2(n_9),
    .B1(u1_n_1015),
    .B2(n_10),
    .Y(n_192));
 AOI22xp33_ASAP7_75t_R g37134 (.A1(u1_n_1041),
    .A2(n_7),
    .B1(u1_n_1014),
    .B2(n_12),
    .Y(n_191));
 AOI22xp33_ASAP7_75t_R g37135 (.A1(u1_n_1039),
    .A2(n_1),
    .B1(u1_n_1012),
    .B2(n_17),
    .Y(n_190));
 AOI22xp33_ASAP7_75t_R g37136 (.A1(u1_n_1026),
    .A2(n_9),
    .B1(u1_n_1053),
    .B2(n_17),
    .Y(n_189));
 AOI22xp33_ASAP7_75t_R g37137 (.A1(u1_n_1027),
    .A2(n_9),
    .B1(u1_n_1054),
    .B2(u1_n_1066),
    .Y(n_188));
 AOI22xp33_ASAP7_75t_R g37138 (.A1(u1_n_1047),
    .A2(n_1),
    .B1(u1_n_1020),
    .B2(n_17),
    .Y(n_187));
 AOI22xp33_ASAP7_75t_R g37139 (.A1(u1_n_1034),
    .A2(n_9),
    .B1(u1_n_1061),
    .B2(n_11),
    .Y(n_186));
 AOI22xp33_ASAP7_75t_R g37140 (.A1(u1_n_1033),
    .A2(n_1),
    .B1(u1_n_1060),
    .B2(n_12),
    .Y(n_185));
 AOI22xp33_ASAP7_75t_R g37141 (.A1(u1_n_1031),
    .A2(n_7),
    .B1(u1_n_1058),
    .B2(n_10),
    .Y(n_184));
 AOI22xp33_ASAP7_75t_R g37142 (.A1(u1_n_1029),
    .A2(n_20),
    .B1(u1_n_1056),
    .B2(n_10),
    .Y(n_183));
 AOI22xp33_ASAP7_75t_R g37143 (.A1(u1_n_1028),
    .A2(n_1),
    .B1(u1_n_1055),
    .B2(n_12),
    .Y(n_182));
 AOI22xp33_ASAP7_75t_R g37144 (.A1(u1_n_1032),
    .A2(n_9),
    .B1(u1_n_1059),
    .B2(n_17),
    .Y(n_181));
 AOI22xp33_ASAP7_75t_R g37145 (.A1(u1_n_1025),
    .A2(n_1),
    .B1(u1_n_1052),
    .B2(n_11),
    .Y(n_180));
 AOI22xp33_ASAP7_75t_R g37146 (.A1(u1_n_1021),
    .A2(n_9),
    .B1(u1_n_1048),
    .B2(u1_n_1066),
    .Y(n_179));
 AOI22xp33_ASAP7_75t_R g37147 (.A1(u1_n_1020),
    .A2(n_9),
    .B1(u1_n_1047),
    .B2(u1_n_1066),
    .Y(n_178));
 AOI22xp33_ASAP7_75t_R g37148 (.A1(u1_n_1017),
    .A2(n_1),
    .B1(u1_n_1044),
    .B2(n_12),
    .Y(n_177));
 AOI22xp33_ASAP7_75t_R g37149 (.A1(u1_n_1030),
    .A2(n_9),
    .B1(u1_n_1057),
    .B2(n_17),
    .Y(n_176));
 AOI22xp33_ASAP7_75t_R g37150 (.A1(u1_n_1013),
    .A2(n_9),
    .B1(u1_n_1040),
    .B2(n_17),
    .Y(n_175));
 AOI22xp33_ASAP7_75t_R g37151 (.A1(u1_n_1012),
    .A2(n_7),
    .B1(u1_n_1039),
    .B2(n_10),
    .Y(n_174));
 AOI22xp33_ASAP7_75t_R g37152 (.A1(u1_n_1024),
    .A2(n_20),
    .B1(u1_n_1051),
    .B2(u1_n_1066),
    .Y(n_173));
 AOI22xp33_ASAP7_75t_R g37153 (.A1(u1_n_1019),
    .A2(n_9),
    .B1(u1_n_1046),
    .B2(n_11),
    .Y(n_172));
 AOI22xp33_ASAP7_75t_R g37154 (.A1(u1_n_1023),
    .A2(n_1),
    .B1(u1_n_1050),
    .B2(u1_n_1066),
    .Y(n_171));
 AOI22xp33_ASAP7_75t_R g37155 (.A1(u1_n_1022),
    .A2(n_20),
    .B1(u1_n_1049),
    .B2(n_12),
    .Y(n_170));
 AOI22xp33_ASAP7_75t_R g37156 (.A1(u1_n_1046),
    .A2(n_7),
    .B1(u1_n_1019),
    .B2(u1_n_1066),
    .Y(n_169));
 AOI22xp33_ASAP7_75t_R g37157 (.A1(u1_n_1018),
    .A2(n_1),
    .B1(u1_n_1045),
    .B2(n_12),
    .Y(n_168));
 AOI22xp33_ASAP7_75t_R g37158 (.A1(u1_n_1040),
    .A2(n_9),
    .B1(u1_n_1013),
    .B2(n_11),
    .Y(n_167));
 AOI22xp33_ASAP7_75t_R g37159 (.A1(u1_n_1048),
    .A2(n_7),
    .B1(u1_n_1021),
    .B2(n_10),
    .Y(n_166));
 XOR2xp5_ASAP7_75t_R g37160 (.A(opa_r[28]),
    .B(opb_r[28]),
    .Y(n_165));
 NOR4xp25_ASAP7_75t_R g37161 (.A(prod[29]),
    .B(prod[34]),
    .C(prod[28]),
    .D(prod[35]),
    .Y(n_164));
 OR4x1_ASAP7_75t_R g37162 (.A(prod[44]),
    .B(prod[43]),
    .C(prod[41]),
    .D(prod[40]),
    .Y(n_163));
 OR4x1_ASAP7_75t_R g37163 (.A(prod[5]),
    .B(prod[4]),
    .C(prod[11]),
    .D(prod[10]),
    .Y(n_162));
 OR4x1_ASAP7_75t_R g37164 (.A(prod[19]),
    .B(prod[16]),
    .C(prod[18]),
    .D(prod[9]),
    .Y(n_161));
 NAND4xp25_ASAP7_75t_R g37165 (.A(u4_exp_div[1]),
    .B(u4_exp_div[2]),
    .C(u4_exp_div[3]),
    .D(u4_exp_div[4]),
    .Y(n_160));
 XOR2xp5_ASAP7_75t_R g37166 (.A(u2_exp_tmp1[1]),
    .B(u2_exp_tmp1[0]),
    .Y(n_159));
 AO22x1_ASAP7_75t_R g37167 (.A1(n_94),
    .A2(u1_n_4761),
    .B1(u1_n_3397),
    .B2(n_14268),
    .Y(n_158));
 XNOR2xp5_ASAP7_75t_R g37168 (.A(opa_r[24]),
    .B(opb_r[24]),
    .Y(n_157));
 XNOR2xp5_ASAP7_75t_R g37169 (.A(opa_r[26]),
    .B(opb_r[26]),
    .Y(n_156));
 XOR2xp5_ASAP7_75t_R g37170 (.A(opa_r[27]),
    .B(opb_r[27]),
    .Y(n_155));
 XNOR2xp5_ASAP7_75t_R g37171 (.A(u2_exp_tmp1[7]),
    .B(u2_n_606),
    .Y(n_199));
 AOI22xp33_ASAP7_75t_R g37172 (.A1(opb_inf),
    .A2(opa_00),
    .B1(opb_00),
    .B2(opa_inf),
    .Y(n_198));
 INVxp33_ASAP7_75t_R g37234 (.A(n_14278),
    .Y(n_154));
 INVxp33_ASAP7_75t_R g37235 (.A(n_150),
    .Y(n_151));
 INVxp33_ASAP7_75t_R g37236 (.A(n_144),
    .Y(n_145));
 INVxp33_ASAP7_75t_R g37237 (.A(n_142),
    .Y(n_143));
 INVxp33_ASAP7_75t_R g37238 (.A(n_140),
    .Y(n_141));
 INVxp33_ASAP7_75t_R g37239 (.A(n_135),
    .Y(n_136));
 INVxp33_ASAP7_75t_R g37240 (.A(n_134),
    .Y(n_133));
 INVxp33_ASAP7_75t_R g37241 (.A(n_132),
    .Y(n_131));
 INVxp33_ASAP7_75t_R g37242 (.A(n_129),
    .Y(n_130));
 INVxp33_ASAP7_75t_R g37243 (.A(n_122),
    .Y(n_121));
 INVxp33_ASAP7_75t_R g37244 (.A(n_120),
    .Y(n_119));
 INVxp33_ASAP7_75t_R g37245 (.A(n_118),
    .Y(n_117));
 INVxp33_ASAP7_75t_R g37246 (.A(n_116),
    .Y(n_115));
 INVxp33_ASAP7_75t_R g37247 (.A(n_114),
    .Y(n_113));
 NOR2xp33_ASAP7_75t_R g37248 (.A(n_24),
    .B(u4_exp_div[7]),
    .Y(n_112));
 NAND2xp33_ASAP7_75t_R g37259 (.A(u1_n_2218),
    .B(u1_n_915),
    .Y(n_110));
 NAND2xp33_ASAP7_75t_R g37263 (.A(n_3494),
    .B(u4_n_1442),
    .Y(n_109));
 NOR2xp33_ASAP7_75t_R g37265 (.A(opb_00),
    .B(opa_inf),
    .Y(n_108));
 NOR2xp33_ASAP7_75t_R g37269 (.A(opb_inf),
    .B(opa_00),
    .Y(n_107));
 NAND2xp33_ASAP7_75t_R g37270 (.A(rmode_r3[1]),
    .B(n_3800),
    .Y(n_106));
 NOR2xp33_ASAP7_75t_R g37272 (.A(n_3807),
    .B(n_3488),
    .Y(n_105));
 NOR2xp33_ASAP7_75t_R g37273 (.A(n_14180),
    .B(n_3567),
    .Y(n_104));
 OR2x2_ASAP7_75t_R g37274 (.A(n_44),
    .B(opb_r[25]),
    .Y(n_103));
 NAND2xp33_ASAP7_75t_R g37275 (.A(n_3495),
    .B(n_3489),
    .Y(n_102));
 NAND2xp33_ASAP7_75t_R g37278 (.A(u2_exp_tmp1[6]),
    .B(n_31),
    .Y(n_152));
 NOR2xp33_ASAP7_75t_R g37279 (.A(opa_00),
    .B(n_34),
    .Y(n_150));
 NAND2xp33_ASAP7_75t_R g37280 (.A(u2_n_1475),
    .B(u2_n_1448),
    .Y(n_101));
 NOR2xp33_ASAP7_75t_R g37281 (.A(opb_00),
    .B(opa_00),
    .Y(n_149));
 NOR2xp33_ASAP7_75t_R g37282 (.A(fasu_op_r2),
    .B(n_70),
    .Y(n_148));
 NAND2xp33_ASAP7_75t_R g37283 (.A(u2_n_1398),
    .B(u2_n_1756),
    .Y(n_147));
 NOR2xp33_ASAP7_75t_R g37285 (.A(opb_inf),
    .B(opa_inf),
    .Y(n_144));
 NAND2xp33_ASAP7_75t_R g37289 (.A(u1_n_853),
    .B(u1_n_996),
    .Y(n_142));
 NAND2xp33_ASAP7_75t_R g37290 (.A(u2_n_1398),
    .B(u2_n_1494),
    .Y(n_140));
 NOR2xp33_ASAP7_75t_R g37291 (.A(n_29),
    .B(u2_n_1493),
    .Y(n_139));
 NOR2xp33_ASAP7_75t_R g37292 (.A(n_3721),
    .B(u4_exp_out[0]),
    .Y(n_138));
 NOR2xp33_ASAP7_75t_R g37293 (.A(exp_ovf_r[1]),
    .B(n_66),
    .Y(n_137));
 NAND2xp33_ASAP7_75t_R g37294 (.A(n_33),
    .B(u2_n_606),
    .Y(n_135));
 NOR2xp33_ASAP7_75t_R g37295 (.A(n_31),
    .B(u2_exp_tmp1[6]),
    .Y(n_134));
 NAND2xp33_ASAP7_75t_R g37296 (.A(n_13920),
    .B(n_3803),
    .Y(n_132));
 NAND2xp33_ASAP7_75t_R g37297 (.A(opa_00),
    .B(opb_00),
    .Y(n_129));
 NOR2xp33_ASAP7_75t_R g37298 (.A(inf_mul2),
    .B(inf_mul_r),
    .Y(n_128));
 NAND2xp33_ASAP7_75t_R g37299 (.A(u2_n_1475),
    .B(u2_n_1494),
    .Y(n_127));
 AND2x2_ASAP7_75t_R g37300 (.A(u4_exp_out[0]),
    .B(n_3721),
    .Y(n_126));
 NAND2xp33_ASAP7_75t_R g37301 (.A(n_29),
    .B(u2_exp_ovf_d[1]),
    .Y(n_125));
 NAND2xp33_ASAP7_75t_R g37302 (.A(u2_n_1489),
    .B(u2_n_1777),
    .Y(n_124));
 NAND2xp33_ASAP7_75t_R g37303 (.A(exp_ovf_r[0]),
    .B(exp_ovf_r[1]),
    .Y(n_123));
 NOR2xp33_ASAP7_75t_R g37304 (.A(u2_exp_tmp1[0]),
    .B(u2_exp_tmp1[1]),
    .Y(n_122));
 NOR2xp33_ASAP7_75t_R g37305 (.A(n_29),
    .B(u2_exp_ovf_d[1]),
    .Y(n_120));
 NAND2xp33_ASAP7_75t_R g37306 (.A(rmode_r3[0]),
    .B(n_66),
    .Y(n_118));
 NOR2xp33_ASAP7_75t_R g37307 (.A(u2_n_775),
    .B(u2_exp_ovf_d[1]),
    .Y(n_116));
 NOR2xp33_ASAP7_75t_R g37308 (.A(qnan_d),
    .B(snan_d),
    .Y(n_114));
 INVxp33_ASAP7_75t_R g37309 (.A(underflow_fmul_r[1]),
    .Y(n_100));
 INVxp33_ASAP7_75t_R g37310 (.A(u1_n_992),
    .Y(n_99));
 INVxp33_ASAP7_75t_R g37312 (.A(u1_n_986),
    .Y(n_97));
 INVxp33_ASAP7_75t_R g37317 (.A(snan_d),
    .Y(n_92));
 INVxp33_ASAP7_75t_R g37322 (.A(n_14094),
    .Y(n_87));
 INVxp33_ASAP7_75t_R g37334 (.A(n_14100),
    .Y(n_75));
 INVxp33_ASAP7_75t_R g37339 (.A(ind_d),
    .Y(n_70));
 INVxp33_ASAP7_75t_R g37340 (.A(u2_exp_tmp1[2]),
    .Y(n_69));
 INVxp33_ASAP7_75t_R g37341 (.A(exp_ovf_r[0]),
    .Y(n_68));
 INVxp33_ASAP7_75t_R g37343 (.A(rmode_r3[1]),
    .Y(n_66));
 INVxp33_ASAP7_75t_R g37344 (.A(n_3530),
    .Y(n_65));
 INVxp33_ASAP7_75t_R g37345 (.A(fpu_op_r1[1]),
    .Y(n_64));
 INVxp33_ASAP7_75t_R g37346 (.A(n_3512),
    .Y(n_63));
 INVxp33_ASAP7_75t_R g37348 (.A(n_3564),
    .Y(n_61));
 INVxp33_ASAP7_75t_R g37350 (.A(n_3769),
    .Y(n_59));
 INVxp33_ASAP7_75t_R g37352 (.A(u1_n_4919),
    .Y(n_57));
 INVxp33_ASAP7_75t_R g37354 (.A(u1_fracta_s[26]),
    .Y(n_55));
 INVxp33_ASAP7_75t_R g37355 (.A(opa_r[23]),
    .Y(n_54));
 INVxp33_ASAP7_75t_R g37356 (.A(n_3558),
    .Y(n_53));
 INVxp33_ASAP7_75t_R g37359 (.A(n_3501),
    .Y(n_50));
 INVxp33_ASAP7_75t_R g37360 (.A(opa_r[28]),
    .Y(n_49));
 INVxp33_ASAP7_75t_R g37361 (.A(u2_n_1384),
    .Y(n_48));
 INVxp33_ASAP7_75t_R g37364 (.A(opa_r[27]),
    .Y(n_45));
 INVxp33_ASAP7_75t_R g37367 (.A(opa_r[29]),
    .Y(n_42));
 INVxp33_ASAP7_75t_R g37369 (.A(n_3722),
    .Y(n_40));
 INVxp33_ASAP7_75t_R g37370 (.A(u4_g),
    .Y(n_39));
 INVxp33_ASAP7_75t_R g37371 (.A(u4_n_1248),
    .Y(n_38));
 INVxp33_ASAP7_75t_R g37372 (.A(n_3723),
    .Y(n_37));
 INVxp33_ASAP7_75t_R g37374 (.A(inf_d),
    .Y(n_35));
 INVxp33_ASAP7_75t_R g37375 (.A(opb_00),
    .Y(n_34));
 INVxp33_ASAP7_75t_R g37376 (.A(u2_exp_tmp1[4]),
    .Y(n_33));
 INVxp33_ASAP7_75t_R g37377 (.A(n_3573),
    .Y(n_32));
 INVxp33_ASAP7_75t_R g37378 (.A(u2_n_606),
    .Y(n_31));
 INVxp33_ASAP7_75t_R g37379 (.A(opa_inf),
    .Y(n_30));
 INVxp33_ASAP7_75t_R g37380 (.A(u2_n_775),
    .Y(n_29));
 INVxp33_ASAP7_75t_R g37381 (.A(n_3724),
    .Y(n_28));
 INVxp33_ASAP7_75t_R g37384 (.A(u2_n_772),
    .Y(n_25));
 INVxp33_ASAP7_75t_R g37387 (.A(n_13920),
    .Y(n_22));
 INVxp33_ASAP7_75t_R g37389 (.A(u1_n_1066),
    .Y(n_20));
 HB1xp67_ASAP7_75t_R g37392 (.A(u1_n_1066),
    .Y(n_17));
 INVxp33_ASAP7_75t_R g37393 (.A(u1_n_1066),
    .Y(n_9));
 AOI221xp5_ASAP7_75t_R g42735 (.A1(u4_exp_div[7]),
    .A2(n_1029),
    .B1(n_3599),
    .B2(u4_n_1851),
    .C(n_1673),
    .Y(n_15699_BAR));
 OAI32xp33_ASAP7_75t_R g42736 (.A1(n_1655),
    .A2(n_3803),
    .A3(rmode_r3[0]),
    .B1(sign),
    .B2(n_1815),
    .Y(n_3577));
 A2O1A1Ixp33_ASAP7_75t_R g42737 (.A1(u4_n_1793),
    .A2(n_1812),
    .B(n_1814),
    .C(n_3801),
    .Y(n_1815));
 OAI21xp33_ASAP7_75t_R g42738 (.A1(n_1808),
    .A2(n_3531),
    .B(n_1813),
    .Y(u4_exp_div[7]));
 NAND4xp25_ASAP7_75t_R g42739 (.A(n_1809),
    .B(n_3592),
    .C(n_989),
    .D(opa_dn),
    .Y(n_3531));
 AOI211xp5_ASAP7_75t_R g42740 (.A1(n_1810),
    .A2(n_3530),
    .B(n_1663),
    .C(n_26),
    .Y(n_1814));
 AOI211xp5_ASAP7_75t_R g42741 (.A1(n_3804),
    .A2(n_1024),
    .B(n_1811),
    .C(n_1805),
    .Y(n_1813));
 OAI211xp5_ASAP7_75t_R g42742 (.A1(exp_ovf_r[0]),
    .A2(n_1801),
    .B(n_1308),
    .C(u4_n_1362),
    .Y(n_1812));
 O2A1O1Ixp33_ASAP7_75t_R g42743 (.A1(n_1803),
    .A2(n_3765),
    .B(n_1806),
    .C(n_3529),
    .Y(n_1811));
 AOI22xp33_ASAP7_75t_R g42744 (.A1(u4_n_1817),
    .A2(n_1804),
    .B1(n_1020),
    .B2(u4_n_1362),
    .Y(n_1810));
 NAND5xp2_ASAP7_75t_R g42745 (.A(n_1807),
    .B(n_3733),
    .C(n_3731),
    .D(n_3732),
    .E(n_1788),
    .Y(n_1809));
 INVxp33_ASAP7_75t_R g42746 (.A(n_1807),
    .Y(n_1808));
 XOR2xp5_ASAP7_75t_R g42747 (.A(n_1802),
    .B(n_3772),
    .Y(n_1807));
 NAND2xp33_ASAP7_75t_R g42748 (.A(n_3765),
    .B(n_1803),
    .Y(n_1806));
 O2A1O1Ixp33_ASAP7_75t_R g42749 (.A1(n_1679),
    .A2(n_1799),
    .B(n_1800),
    .C(n_3528),
    .Y(n_1805));
 NAND2xp33_ASAP7_75t_R g42750 (.A(n_1020),
    .B(u4_exp_out1_co),
    .Y(n_1804));
 NOR2xp33_ASAP7_75t_R g42751 (.A(n_3850),
    .B(n_1801),
    .Y(n_3760));
 AOI21xp33_ASAP7_75t_R g42752 (.A1(n_1785),
    .A2(n_1797),
    .B(n_1786),
    .Y(n_1802));
 OR3x1_ASAP7_75t_R g42753 (.A(n_3764),
    .B(n_3729),
    .C(n_3728),
    .Y(n_1803));
 INVxp33_ASAP7_75t_R g42754 (.A(u4_exp_out1_co),
    .Y(n_1801));
 XOR2xp5_ASAP7_75t_R g42755 (.A(n_1797),
    .B(n_1790),
    .Y(n_3731));
 XOR2xp5_ASAP7_75t_R g42756 (.A(n_1798),
    .B(n_3573),
    .Y(u4_exp_out1_co));
 NAND2xp33_ASAP7_75t_R g42757 (.A(n_1679),
    .B(n_1799),
    .Y(n_1800));
 XOR2xp5_ASAP7_75t_R g42758 (.A(n_1795),
    .B(n_1789),
    .Y(n_3733));
 OAI21xp33_ASAP7_75t_R g42759 (.A1(n_1076),
    .A2(n_1796),
    .B(n_1798),
    .Y(n_3765));
 A2O1A1Ixp33_ASAP7_75t_R g42760 (.A1(n_14181),
    .A2(n_3560),
    .B(n_1677),
    .C(n_3586),
    .Y(n_1799));
 NAND2xp33_ASAP7_75t_R g42761 (.A(n_1796),
    .B(n_1076),
    .Y(n_1798));
 AO21x1_ASAP7_75t_R g42762 (.A1(n_3773),
    .A2(n_1791),
    .B(n_1796),
    .Y(n_3764));
 XNOR2xp5_ASAP7_75t_R g42763 (.A(n_1787),
    .B(n_1667),
    .Y(n_3804));
 OAI21xp33_ASAP7_75t_R g42764 (.A1(n_1789),
    .A2(n_1793),
    .B(n_1794),
    .Y(n_1797));
 NAND2xp33_ASAP7_75t_R g42765 (.A(n_1794),
    .B(n_1792),
    .Y(n_1795));
 NOR2xp33_ASAP7_75t_R g42766 (.A(n_3773),
    .B(n_1791),
    .Y(n_1796));
 OR2x2_ASAP7_75t_R g42767 (.A(n_3762),
    .B(n_3763),
    .Y(n_3729));
 XOR2xp5_ASAP7_75t_R g42768 (.A(n_1783),
    .B(n_1778),
    .Y(n_3732));
 INVxp33_ASAP7_75t_R g42769 (.A(n_1792),
    .Y(n_1793));
 NOR2xp33_ASAP7_75t_R g42770 (.A(n_1784),
    .B(n_1786),
    .Y(n_1790));
 NAND2xp33_ASAP7_75t_R g42771 (.A(n_3775),
    .B(n_1782),
    .Y(n_1794));
 NAND2xp33_ASAP7_75t_R g42772 (.A(n_1069),
    .B(n_3734),
    .Y(n_1792));
 OAI21xp33_ASAP7_75t_R g42773 (.A1(n_1762),
    .A2(n_1777),
    .B(n_1759),
    .Y(n_1791));
 AND5x1_ASAP7_75t_R g42774 (.A(n_3737),
    .B(n_3736),
    .C(n_1743),
    .D(n_1742),
    .E(n_3740),
    .Y(n_1788));
 XNOR2xp5_ASAP7_75t_R g42775 (.A(n_1777),
    .B(n_1768),
    .Y(n_3763));
 A2O1A1Ixp33_ASAP7_75t_R g42776 (.A1(n_3812),
    .A2(n_3561),
    .B(n_1665),
    .C(n_3810),
    .Y(n_1787));
 AOI21xp33_ASAP7_75t_R g42777 (.A1(n_1780),
    .A2(n_1778),
    .B(n_1779),
    .Y(n_1789));
 INVxp33_ASAP7_75t_R g42778 (.A(n_1784),
    .Y(n_1785));
 AND2x2_ASAP7_75t_R g42779 (.A(n_3773),
    .B(n_3524),
    .Y(n_1786));
 NOR2xp33_ASAP7_75t_R g42780 (.A(n_3773),
    .B(n_3524),
    .Y(n_1784));
 NOR2xp33_ASAP7_75t_R g42781 (.A(n_1779),
    .B(n_1781),
    .Y(n_1783));
 INVxp33_ASAP7_75t_R g42782 (.A(n_1782),
    .Y(n_3734));
 NAND3xp33_ASAP7_75t_R g42783 (.A(n_3585),
    .B(n_3511),
    .C(n_3510),
    .Y(n_3560));
 XOR2xp5_ASAP7_75t_R g42784 (.A(n_1776),
    .B(n_1769),
    .Y(n_3737));
 OAI21xp33_ASAP7_75t_R g42785 (.A1(n_1643),
    .A2(n_1775),
    .B(n_3524),
    .Y(n_1782));
 INVxp33_ASAP7_75t_R g42786 (.A(n_1780),
    .Y(n_1781));
 NAND2xp33_ASAP7_75t_R g42787 (.A(n_14182),
    .B(n_3735),
    .Y(n_1780));
 NOR2xp33_ASAP7_75t_R g42788 (.A(n_14182),
    .B(n_3735),
    .Y(n_1779));
 NAND2xp33_ASAP7_75t_R g42789 (.A(n_1775),
    .B(n_1643),
    .Y(n_3524));
 OR3x1_ASAP7_75t_R g42790 (.A(n_3761),
    .B(n_3521),
    .C(n_1746),
    .Y(n_3728));
 XNOR2xp5_ASAP7_75t_R g42791 (.A(n_1767),
    .B(n_1770),
    .Y(n_3762));
 OAI21xp33_ASAP7_75t_R g42792 (.A1(n_1769),
    .A2(n_1772),
    .B(n_1774),
    .Y(n_1778));
 AOI21xp33_ASAP7_75t_R g42793 (.A1(n_1770),
    .A2(n_1755),
    .B(n_1761),
    .Y(n_1777));
 NAND2xp33_ASAP7_75t_R g42794 (.A(n_3589),
    .B(n_1771),
    .Y(n_3585));
 NAND2xp33_ASAP7_75t_R g42795 (.A(n_1774),
    .B(n_1773),
    .Y(n_1776));
 NAND3xp33_ASAP7_75t_R g42796 (.A(n_3574),
    .B(n_3817),
    .C(n_3509),
    .Y(n_3561));
 OAI21xp33_ASAP7_75t_R g42797 (.A1(n_1651),
    .A2(n_1765),
    .B(n_1653),
    .Y(n_1775));
 XOR2xp5_ASAP7_75t_R g42798 (.A(n_1763),
    .B(n_1754),
    .Y(n_3736));
 XNOR2xp5_ASAP7_75t_R g42799 (.A(n_1764),
    .B(n_1660),
    .Y(n_3735));
 INVxp33_ASAP7_75t_R g42800 (.A(n_1772),
    .Y(n_1773));
 A2O1A1Ixp33_ASAP7_75t_R g42801 (.A1(n_3518),
    .A2(n_3590),
    .B(n_1715),
    .C(n_3520),
    .Y(n_1771));
 NAND2xp33_ASAP7_75t_R g42802 (.A(n_3768),
    .B(n_1766),
    .Y(n_1774));
 NOR2xp33_ASAP7_75t_R g42803 (.A(n_3768),
    .B(n_1766),
    .Y(n_1772));
 XOR2xp5_ASAP7_75t_R g42804 (.A(n_1760),
    .B(n_1752),
    .Y(n_3761));
 OAI21xp33_ASAP7_75t_R g42805 (.A1(n_1753),
    .A2(n_1747),
    .B(n_1749),
    .Y(n_1770));
 AOI21xp33_ASAP7_75t_R g42806 (.A1(n_1757),
    .A2(n_1754),
    .B(n_1756),
    .Y(n_1769));
 AOI21xp33_ASAP7_75t_R g42807 (.A1(n_1748),
    .A2(n_3775),
    .B(n_1762),
    .Y(n_1768));
 NAND2xp33_ASAP7_75t_R g42808 (.A(n_3821),
    .B(n_1751),
    .Y(n_3817));
 OAI21xp33_ASAP7_75t_R g42809 (.A1(n_14182),
    .A2(n_3776),
    .B(n_1755),
    .Y(n_1767));
 INVxp33_ASAP7_75t_R g42810 (.A(n_1766),
    .Y(n_3738));
 INVxp33_ASAP7_75t_R g42811 (.A(n_1764),
    .Y(n_1765));
 NOR2xp33_ASAP7_75t_R g42812 (.A(n_1756),
    .B(n_1758),
    .Y(n_1763));
 XNOR2xp5_ASAP7_75t_R g42813 (.A(n_1745),
    .B(n_1662),
    .Y(n_1766));
 OAI21xp33_ASAP7_75t_R g42814 (.A1(n_1649),
    .A2(n_1745),
    .B(n_1654),
    .Y(n_1764));
 NAND2xp33_ASAP7_75t_R g42815 (.A(n_3598),
    .B(n_3757),
    .Y(n_3578));
 NOR2xp33_ASAP7_75t_R g42816 (.A(n_14182),
    .B(n_3776),
    .Y(n_1761));
 NOR2xp33_ASAP7_75t_R g42817 (.A(n_1747),
    .B(n_1750),
    .Y(n_1760));
 NOR2xp33_ASAP7_75t_R g42818 (.A(n_3775),
    .B(n_1748),
    .Y(n_1762));
 NAND2xp33_ASAP7_75t_R g42819 (.A(n_3775),
    .B(n_1748),
    .Y(n_1759));
 INVxp33_ASAP7_75t_R g42820 (.A(n_1757),
    .Y(n_1758));
 INVxp33_ASAP7_75t_R g42821 (.A(n_1752),
    .Y(n_1753));
 A2O1A1Ixp33_ASAP7_75t_R g42822 (.A1(n_3517),
    .A2(n_3818),
    .B(n_1686),
    .C(n_3519),
    .Y(n_1751));
 NAND2xp33_ASAP7_75t_R g42823 (.A(n_1014),
    .B(n_3739),
    .Y(n_1757));
 NOR2xp33_ASAP7_75t_R g42824 (.A(n_1014),
    .B(n_3739),
    .Y(n_1756));
 NAND2xp33_ASAP7_75t_R g42825 (.A(n_14182),
    .B(n_3776),
    .Y(n_1755));
 MAJIxp5_ASAP7_75t_R g42826 (.A(n_1737),
    .B(n_3820),
    .C(n_3741),
    .Y(n_1754));
 MAJIxp5_ASAP7_75t_R g42827 (.A(n_3770),
    .B(n_1014),
    .C(n_1740),
    .Y(n_1752));
 INVxp33_ASAP7_75t_R g42828 (.A(n_1749),
    .Y(n_1750));
 NAND2xp33_ASAP7_75t_R g42829 (.A(n_3768),
    .B(n_1741),
    .Y(n_1749));
 AND2x2_ASAP7_75t_R g42830 (.A(n_3523),
    .B(n_3568),
    .Y(n_3757));
 NAND2xp33_ASAP7_75t_R g42831 (.A(n_1643),
    .B(n_1744),
    .Y(n_1748));
 NOR2xp33_ASAP7_75t_R g42832 (.A(n_3768),
    .B(n_1741),
    .Y(n_1747));
 OAI21xp33_ASAP7_75t_R g42833 (.A1(n_1718),
    .A2(n_1736),
    .B(n_1717),
    .Y(n_3590));
 INVxp33_ASAP7_75t_R g42834 (.A(n_1746),
    .Y(n_3805));
 NAND2xp33_ASAP7_75t_R g42835 (.A(n_1742),
    .B(n_1743),
    .Y(n_3730));
 XOR2xp5_ASAP7_75t_R g42836 (.A(n_3818),
    .B(n_1692),
    .Y(n_1746));
 AOI21xp33_ASAP7_75t_R g42837 (.A1(n_1691),
    .A2(n_1739),
    .B(n_1690),
    .Y(n_1745));
 XNOR2xp5_ASAP7_75t_R g42838 (.A(n_1739),
    .B(n_1696),
    .Y(n_3739));
 OAI21xp33_ASAP7_75t_R g42839 (.A1(n_3516),
    .A2(n_1738),
    .B(n_1744),
    .Y(n_3776));
 NAND3xp33_ASAP7_75t_R g42840 (.A(n_3727),
    .B(n_1733),
    .C(n_1732),
    .Y(n_3521));
 NAND2xp33_ASAP7_75t_R g42841 (.A(n_3516),
    .B(n_1738),
    .Y(n_1744));
 OR2x2_ASAP7_75t_R g42842 (.A(n_3516),
    .B(n_3758),
    .Y(n_3568));
 INVxp33_ASAP7_75t_R g42843 (.A(n_1741),
    .Y(n_3767));
 NAND2xp33_ASAP7_75t_R g42844 (.A(n_1720),
    .B(n_1736),
    .Y(n_1743));
 OR2x2_ASAP7_75t_R g42845 (.A(n_1720),
    .B(n_1736),
    .Y(n_1742));
 MAJx2_ASAP7_75t_R g42846 (.A(n_3766),
    .B(n_3820),
    .C(n_1724),
    .Y(n_1740));
 AOI21xp33_ASAP7_75t_R g42847 (.A1(n_1734),
    .A2(n_3593),
    .B(n_1738),
    .Y(n_1741));
 NAND2xp33_ASAP7_75t_R g42848 (.A(n_3593),
    .B(n_1735),
    .Y(n_3758));
 NOR2xp33_ASAP7_75t_R g42849 (.A(u4_sll_315_50_n_29),
    .B(n_1731),
    .Y(n_1737));
 OAI21xp33_ASAP7_75t_R g42850 (.A1(n_1709),
    .A2(n_1729),
    .B(n_1708),
    .Y(n_1739));
 NOR2xp33_ASAP7_75t_R g42851 (.A(n_3593),
    .B(n_1734),
    .Y(n_1738));
 NAND2xp33_ASAP7_75t_R g42852 (.A(n_1732),
    .B(n_1733),
    .Y(n_3808));
 XNOR2xp5_ASAP7_75t_R g42853 (.A(n_1729),
    .B(n_1714),
    .Y(n_3741));
 AOI21xp33_ASAP7_75t_R g42854 (.A1(n_1730),
    .A2(n_1117),
    .B(n_1728),
    .Y(n_1736));
 OAI21xp33_ASAP7_75t_R g42855 (.A1(n_3515),
    .A2(n_1725),
    .B(n_1734),
    .Y(n_3770));
 AO21x1_ASAP7_75t_R g42856 (.A1(n_1706),
    .A2(n_1728),
    .B(n_1707),
    .Y(n_3818));
 INVxp33_ASAP7_75t_R g42857 (.A(n_1735),
    .Y(n_3565));
 NAND2xp33_ASAP7_75t_R g42858 (.A(n_3759),
    .B(n_1726),
    .Y(n_3766));
 NOR2xp33_ASAP7_75t_R g42859 (.A(n_3515),
    .B(n_3759),
    .Y(n_1735));
 NAND2xp33_ASAP7_75t_R g42860 (.A(n_1730),
    .B(n_1727),
    .Y(n_3727));
 NAND2xp33_ASAP7_75t_R g42861 (.A(n_3515),
    .B(n_1725),
    .Y(n_1734));
 INVxp33_ASAP7_75t_R g42862 (.A(n_1731),
    .Y(n_3742));
 NAND2xp33_ASAP7_75t_R g42863 (.A(n_1711),
    .B(n_1727),
    .Y(n_1733));
 NAND2xp33_ASAP7_75t_R g42864 (.A(n_1712),
    .B(n_1728),
    .Y(n_1732));
 OAI21xp33_ASAP7_75t_R g42865 (.A1(div_opa_ldz_r2[0]),
    .A2(n_3595),
    .B(n_1729),
    .Y(n_1731));
 XNOR2xp5_ASAP7_75t_R g42866 (.A(n_3595),
    .B(n_3717),
    .Y(n_3740));
 INVxp33_ASAP7_75t_R g42867 (.A(n_1728),
    .Y(n_1727));
 NAND2xp33_ASAP7_75t_R g42868 (.A(n_13972),
    .B(n_3595),
    .Y(n_1730));
 NAND2xp33_ASAP7_75t_R g42869 (.A(div_opa_ldz_r2[0]),
    .B(n_3595),
    .Y(n_1729));
 NOR2xp33_ASAP7_75t_R g42870 (.A(exp_r[0]),
    .B(n_3595),
    .Y(n_1728));
 INVxp33_ASAP7_75t_R g42871 (.A(n_1725),
    .Y(n_1726));
 NOR2xp33_ASAP7_75t_R g42872 (.A(n_702),
    .B(n_3595),
    .Y(n_1724));
 NAND2xp33_ASAP7_75t_R g42873 (.A(n_1704),
    .B(n_3595),
    .Y(n_3759));
 NOR2xp33_ASAP7_75t_R g42874 (.A(n_1704),
    .B(n_3595),
    .Y(n_1725));
 OAI21xp33_ASAP7_75t_R g42875 (.A1(fract_denorm[46]),
    .A2(n_1723),
    .B(n_1575),
    .Y(n_3595));
 O2A1O1Ixp33_ASAP7_75t_R g42876 (.A1(n_1722),
    .A2(fract_denorm[43]),
    .B(n_1586),
    .C(fract_denorm[45]),
    .Y(n_1723));
 O2A1O1Ixp33_ASAP7_75t_R g42877 (.A1(n_1721),
    .A2(fract_denorm[40]),
    .B(n_1578),
    .C(fract_denorm[42]),
    .Y(n_1722));
 O2A1O1Ixp33_ASAP7_75t_R g42878 (.A1(n_1719),
    .A2(fract_denorm[37]),
    .B(n_1587),
    .C(fract_denorm[39]),
    .Y(n_1721));
 AOI21xp33_ASAP7_75t_R g42879 (.A1(n_1716),
    .A2(n_13972),
    .B(n_1718),
    .Y(n_1720));
 O2A1O1Ixp33_ASAP7_75t_R g42880 (.A1(n_1713),
    .A2(fract_denorm[34]),
    .B(n_1576),
    .C(fract_denorm[36]),
    .Y(n_1719));
 NAND2xp33_ASAP7_75t_R g42881 (.A(n_1716),
    .B(n_13972),
    .Y(n_1717));
 NOR2xp33_ASAP7_75t_R g42882 (.A(n_13972),
    .B(n_1716),
    .Y(n_1718));
 XOR2xp5_ASAP7_75t_R g42883 (.A(exp_r[1]),
    .B(n_1714),
    .Y(n_1716));
 NAND2xp33_ASAP7_75t_R g42884 (.A(n_1697),
    .B(n_1710),
    .Y(n_3518));
 INVxp33_ASAP7_75t_R g42885 (.A(n_1715),
    .Y(n_3591));
 NOR2xp33_ASAP7_75t_R g42886 (.A(n_1697),
    .B(n_1710),
    .Y(n_1715));
 O2A1O1Ixp33_ASAP7_75t_R g42887 (.A1(n_1703),
    .A2(fract_denorm[31]),
    .B(n_1590),
    .C(fract_denorm[33]),
    .Y(n_1713));
 AOI21xp33_ASAP7_75t_R g42888 (.A1(n_1704),
    .A2(div_opa_ldz_r2[1]),
    .B(n_1709),
    .Y(n_1714));
 INVxp33_ASAP7_75t_R g42889 (.A(n_1711),
    .Y(n_1712));
 NOR2xp33_ASAP7_75t_R g42890 (.A(n_1705),
    .B(n_1707),
    .Y(n_1711));
 AOI21xp33_ASAP7_75t_R g42891 (.A1(n_3575),
    .A2(n_3514),
    .B(n_1131),
    .Y(n_1710));
 NAND2xp33_ASAP7_75t_R g42892 (.A(div_opa_ldz_r2[1]),
    .B(n_1704),
    .Y(n_1708));
 NOR2xp33_ASAP7_75t_R g42893 (.A(div_opa_ldz_r2[1]),
    .B(n_1704),
    .Y(n_1709));
 INVxp33_ASAP7_75t_R g42894 (.A(n_1705),
    .Y(n_1706));
 NOR2xp33_ASAP7_75t_R g42895 (.A(n_1704),
    .B(u4_sll_315_50_n_6),
    .Y(n_1707));
 NOR2xp33_ASAP7_75t_R g42896 (.A(n_3514),
    .B(n_3820),
    .Y(n_1705));
 INVxp33_ASAP7_75t_R g42897 (.A(n_1704),
    .Y(n_3514));
 O2A1O1Ixp33_ASAP7_75t_R g42898 (.A1(n_1702),
    .A2(fract_denorm[44]),
    .B(n_1612),
    .C(fract_denorm[47]),
    .Y(n_1704));
 O2A1O1Ixp33_ASAP7_75t_R g42899 (.A1(n_1701),
    .A2(fract_denorm[28]),
    .B(n_1588),
    .C(fract_denorm[30]),
    .Y(n_1703));
 AO21x1_ASAP7_75t_R g42900 (.A1(n_1593),
    .A2(n_1700),
    .B(fract_denorm[43]),
    .Y(n_1702));
 O2A1O1Ixp33_ASAP7_75t_R g42901 (.A1(n_1699),
    .A2(fract_denorm[25]),
    .B(n_1589),
    .C(fract_denorm[27]),
    .Y(n_1701));
 OAI21xp33_ASAP7_75t_R g42902 (.A1(n_1598),
    .A2(n_1698),
    .B(n_1595),
    .Y(n_1700));
 O2A1O1Ixp33_ASAP7_75t_R g42903 (.A1(n_1695),
    .A2(fract_denorm[22]),
    .B(n_1577),
    .C(fract_denorm[24]),
    .Y(n_1699));
 AOI211xp5_ASAP7_75t_R g42904 (.A1(n_1693),
    .A2(n_1599),
    .B(fract_denorm[35]),
    .C(fract_denorm[36]),
    .Y(n_1698));
 XOR2xp5_ASAP7_75t_R g42905 (.A(exp_r[2]),
    .B(n_1696),
    .Y(n_1697));
 NAND2xp33_ASAP7_75t_R g42906 (.A(n_1694),
    .B(n_1670),
    .Y(n_3589));
 OR2x2_ASAP7_75t_R g42907 (.A(n_1670),
    .B(n_1694),
    .Y(n_3520));
 O2A1O1Ixp33_ASAP7_75t_R g42908 (.A1(n_1684),
    .A2(fract_denorm[19]),
    .B(n_1591),
    .C(fract_denorm[21]),
    .Y(n_1695));
 NAND2xp33_ASAP7_75t_R g42909 (.A(n_1691),
    .B(n_1689),
    .Y(n_1696));
 A2O1A1Ixp33_ASAP7_75t_R g42910 (.A1(n_1606),
    .A2(n_1683),
    .B(u4_n_1942),
    .C(n_1604),
    .Y(n_1693));
 NAND2xp33_ASAP7_75t_R g42911 (.A(n_3823),
    .B(n_3517),
    .Y(n_1692));
 NAND2xp33_ASAP7_75t_R g42912 (.A(n_3582),
    .B(n_1688),
    .Y(n_1694));
 INVxp33_ASAP7_75t_R g42913 (.A(n_1689),
    .Y(n_1690));
 NAND2xp33_ASAP7_75t_R g42914 (.A(n_3515),
    .B(n_3563),
    .Y(n_1688));
 NAND2xp33_ASAP7_75t_R g42915 (.A(n_1130),
    .B(n_3515),
    .Y(n_1691));
 NAND2xp33_ASAP7_75t_R g42916 (.A(div_opa_ldz_r2[2]),
    .B(n_1685),
    .Y(n_1689));
 INVxp33_ASAP7_75t_R g42918 (.A(n_3823),
    .Y(n_1686));
 OR2x2_ASAP7_75t_R g42920 (.A(n_3515),
    .B(n_3824),
    .Y(n_3517));
 NAND2xp33_ASAP7_75t_R g42921 (.A(n_3515),
    .B(n_3824),
    .Y(n_3823));
 NOR2xp33_ASAP7_75t_R g42922 (.A(n_3803),
    .B(u4_f2i_zero),
    .Y(n_3597));
 OAI211xp5_ASAP7_75t_R g42924 (.A1(n_1616),
    .A2(n_1678),
    .B(n_1612),
    .C(n_1575),
    .Y(n_3515));
 O2A1O1Ixp33_ASAP7_75t_R g42925 (.A1(n_1676),
    .A2(fract_denorm[16]),
    .B(n_1585),
    .C(fract_denorm[18]),
    .Y(n_1684));
 NAND2xp33_ASAP7_75t_R g42926 (.A(n_1682),
    .B(n_1659),
    .Y(n_3588));
 A2O1A1Ixp33_ASAP7_75t_R g42927 (.A1(n_1600),
    .A2(n_1675),
    .B(u4_n_1944),
    .C(n_1605),
    .Y(n_1683));
 OR2x2_ASAP7_75t_R g42928 (.A(n_1659),
    .B(n_1682),
    .Y(n_3511));
 OAI22xp33_ASAP7_75t_R g42929 (.A1(n_1680),
    .A2(n_3755),
    .B1(n_1002),
    .B2(n_3754),
    .Y(u4_f2i_zero));
 XNOR2xp5_ASAP7_75t_R g42930 (.A(n_1666),
    .B(div_opa_ldz_r2[4]),
    .Y(n_1682));
 INVxp33_ASAP7_75t_R g42931 (.A(n_3510),
    .Y(n_1681));
 NAND2xp33_ASAP7_75t_R g42932 (.A(n_1669),
    .B(n_1671),
    .Y(n_3587));
 OAI221xp5_ASAP7_75t_R g42933 (.A1(exp_r[5]),
    .A2(n_3508),
    .B1(exp_r[6]),
    .B2(n_46),
    .C(n_1664),
    .Y(n_3586));
 NAND2xp33_ASAP7_75t_R g42934 (.A(n_1668),
    .B(n_1672),
    .Y(n_3510));
 INVxp33_ASAP7_75t_R g42935 (.A(n_3572),
    .Y(n_1680));
 AOI211xp5_ASAP7_75t_R g42936 (.A1(n_1661),
    .A2(n_1618),
    .B(n_1596),
    .C(n_1598),
    .Y(n_1678));
 NAND4xp25_ASAP7_75t_R g42937 (.A(n_3532),
    .B(opas_r2),
    .C(rmode_r3[1]),
    .D(rmode_r3[0]),
    .Y(n_3572));
 NAND2xp33_ASAP7_75t_R g42938 (.A(n_3574),
    .B(n_1674),
    .Y(n_3812));
 XNOR2xp5_ASAP7_75t_R g42939 (.A(n_1664),
    .B(exp_r[7]),
    .Y(n_1679));
 INVxp33_ASAP7_75t_R g42940 (.A(n_1677),
    .Y(n_3526));
 O2A1O1Ixp33_ASAP7_75t_R g42941 (.A1(n_1650),
    .A2(fract_denorm[13]),
    .B(n_1569),
    .C(fract_denorm[15]),
    .Y(n_1676));
 OAI31xp33_ASAP7_75t_R g42942 (.A1(fract_denorm[17]),
    .A2(n_1646),
    .A3(fract_denorm[18]),
    .B(n_1592),
    .Y(n_1675));
 NAND2xp33_ASAP7_75t_R g42943 (.A(n_3815),
    .B(n_3825),
    .Y(n_1674));
 NOR2xp33_ASAP7_75t_R g42944 (.A(exp_r[5]),
    .B(n_1664),
    .Y(n_1677));
 NOR2xp33_ASAP7_75t_R g42945 (.A(n_3594),
    .B(n_1663),
    .Y(n_3598));
 INVxp33_ASAP7_75t_R g42946 (.A(n_1673),
    .Y(n_3562));
 INVxp33_ASAP7_75t_R g42947 (.A(n_1671),
    .Y(n_1672));
 INVxp33_ASAP7_75t_R g42948 (.A(n_1668),
    .Y(n_1669));
 NOR3xp33_ASAP7_75t_R g42949 (.A(n_3532),
    .B(n_3594),
    .C(n_1002),
    .Y(n_1673));
 OAI21xp33_ASAP7_75t_R g42950 (.A1(n_1658),
    .A2(n_1119),
    .B(n_3583),
    .Y(n_1671));
 XOR2xp5_ASAP7_75t_R g42951 (.A(exp_r[3]),
    .B(n_1662),
    .Y(n_1670));
 XNOR2xp5_ASAP7_75t_R g42952 (.A(n_1070),
    .B(n_46),
    .Y(n_1667));
 XNOR2xp5_ASAP7_75t_R g42953 (.A(exp_r[4]),
    .B(n_1658),
    .Y(n_1666));
 OAI22xp33_ASAP7_75t_R g42954 (.A1(n_3508),
    .A2(n_700),
    .B1(n_46),
    .B2(exp_r[5]),
    .Y(n_1668));
 INVxp33_ASAP7_75t_R g42955 (.A(n_1665),
    .Y(n_3522));
 NOR2xp33_ASAP7_75t_R g42956 (.A(n_3508),
    .B(n_3811),
    .Y(n_1665));
 NAND2xp33_ASAP7_75t_R g42957 (.A(n_3508),
    .B(n_3811),
    .Y(n_3810));
 OR2x2_ASAP7_75t_R g42958 (.A(n_3508),
    .B(n_3816),
    .Y(n_3574));
 NAND2xp33_ASAP7_75t_R g42959 (.A(n_46),
    .B(exp_r[6]),
    .Y(n_1664));
 INVxp33_ASAP7_75t_R g42960 (.A(n_1663),
    .Y(n_3532));
 NAND2xp33_ASAP7_75t_R g42961 (.A(n_1657),
    .B(n_3826),
    .Y(n_3825));
 NAND2xp33_ASAP7_75t_R g42962 (.A(n_1658),
    .B(n_1055),
    .Y(n_3509));
 NAND2xp33_ASAP7_75t_R g42963 (.A(n_3816),
    .B(n_3508),
    .Y(n_3815));
 NOR5xp2_ASAP7_75t_R g42964 (.A(n_1641),
    .B(n_1629),
    .C(n_1631),
    .D(n_1624),
    .E(fract_denorm[24]),
    .Y(n_1663));
 OR3x1_ASAP7_75t_R g42965 (.A(n_1644),
    .B(u4_n_1938),
    .C(u4_n_1942),
    .Y(n_1661));
 NAND2xp33_ASAP7_75t_R g42966 (.A(n_1652),
    .B(n_1653),
    .Y(n_1660));
 OAI21xp33_ASAP7_75t_R g42967 (.A1(div_opa_ldz_r2[3]),
    .A2(n_3593),
    .B(n_1654),
    .Y(n_1662));
 INVxp33_ASAP7_75t_R g42968 (.A(n_1658),
    .Y(n_1657));
 INVxp33_ASAP7_75t_R g42969 (.A(n_46),
    .Y(n_3508));
 AOI31xp33_ASAP7_75t_R g42970 (.A1(n_24),
    .A2(n_1641),
    .A3(n_1002),
    .B(u4_n_1830),
    .Y(n_1655));
 NAND2xp33_ASAP7_75t_R g42971 (.A(n_3580),
    .B(n_1647),
    .Y(n_1659));
 AOI21xp33_ASAP7_75t_R g42972 (.A1(n_98),
    .A2(n_3516),
    .B(n_1648),
    .Y(n_1658));
 NOR2xp33_ASAP7_75t_R g42973 (.A(n_1643),
    .B(n_1648),
    .Y(n_46));
 INVxp33_ASAP7_75t_R g42974 (.A(n_1651),
    .Y(n_1652));
 O2A1O1Ixp33_ASAP7_75t_R g42975 (.A1(n_1639),
    .A2(fract_denorm[10]),
    .B(n_1570),
    .C(fract_denorm[12]),
    .Y(n_1650));
 NAND2xp33_ASAP7_75t_R g42976 (.A(div_opa_ldz_r2[3]),
    .B(n_3593),
    .Y(n_1654));
 NOR2xp33_ASAP7_75t_R g42977 (.A(div_opa_ldz_r2[3]),
    .B(n_3593),
    .Y(n_1649));
 NAND2xp33_ASAP7_75t_R g42978 (.A(div_opa_ldz_r2[4]),
    .B(n_1645),
    .Y(n_1653));
 NOR2xp33_ASAP7_75t_R g42979 (.A(div_opa_ldz_r2[4]),
    .B(n_1645),
    .Y(n_1651));
 NAND2xp33_ASAP7_75t_R g42980 (.A(n_3593),
    .B(n_3506),
    .Y(n_1647));
 NOR3xp33_ASAP7_75t_R g42981 (.A(n_1640),
    .B(fract_denorm[16]),
    .C(fract_denorm[15]),
    .Y(n_1646));
 NOR2xp33_ASAP7_75t_R g42982 (.A(n_98),
    .B(n_3516),
    .Y(n_1648));
 OR2x2_ASAP7_75t_R g42983 (.A(n_3593),
    .B(n_3822),
    .Y(n_3519));
 NAND2xp33_ASAP7_75t_R g42984 (.A(n_3822),
    .B(n_3593),
    .Y(n_3821));
 INVxp33_ASAP7_75t_R g42985 (.A(n_1645),
    .Y(n_3516));
 AOI31xp33_ASAP7_75t_R g42986 (.A1(n_1633),
    .A2(n_1603),
    .A3(n_1600),
    .B(n_1613),
    .Y(n_1644));
 O2A1O1Ixp33_ASAP7_75t_R g42987 (.A1(n_1634),
    .A2(n_1631),
    .B(n_1638),
    .C(n_1629),
    .Y(n_1645));
 INVxp33_ASAP7_75t_R g42988 (.A(n_1643),
    .Y(n_3523));
 NOR5xp2_ASAP7_75t_R g42990 (.A(n_1630),
    .B(n_3505),
    .C(n_1624),
    .D(n_1626),
    .E(fract_denorm[47]),
    .Y(n_1643));
 OAI32xp33_ASAP7_75t_R g42991 (.A1(n_1614),
    .A2(n_1636),
    .A3(n_1624),
    .B1(n_1637),
    .B2(n_1631),
    .Y(n_3593));
 NAND3xp33_ASAP7_75t_R g42992 (.A(n_1632),
    .B(n_1614),
    .C(n_1577),
    .Y(n_1641));
 OAI32xp33_ASAP7_75t_R g42993 (.A1(fract_denorm[9]),
    .A2(n_1628),
    .A3(fract_denorm[10]),
    .B1(n_1580),
    .B2(n_1572),
    .Y(n_1640));
 O2A1O1Ixp33_ASAP7_75t_R g42994 (.A1(n_1622),
    .A2(fract_denorm[7]),
    .B(n_1568),
    .C(fract_denorm[9]),
    .Y(n_1639));
 NAND2xp33_ASAP7_75t_R g42995 (.A(n_1614),
    .B(n_1635),
    .Y(n_1638));
 AOI21xp33_ASAP7_75t_R g42996 (.A1(n_1623),
    .A2(n_1630),
    .B(n_1629),
    .Y(n_1637));
 INVxp33_ASAP7_75t_R g42997 (.A(n_1635),
    .Y(n_1636));
 NOR2xp33_ASAP7_75t_R g42998 (.A(n_1624),
    .B(n_1630),
    .Y(n_1634));
 NOR2xp33_ASAP7_75t_R g42999 (.A(n_1621),
    .B(n_1631),
    .Y(n_1635));
 A2O1A1Ixp33_ASAP7_75t_R g43000 (.A1(n_1611),
    .A2(n_1620),
    .B(n_1610),
    .C(n_1617),
    .Y(n_1633));
 NOR3xp33_ASAP7_75t_R g43001 (.A(n_1621),
    .B(n_1627),
    .C(fract_denorm[0]),
    .Y(n_1632));
 OR2x2_ASAP7_75t_R g43002 (.A(n_1596),
    .B(n_1625),
    .Y(n_3505));
 OR2x2_ASAP7_75t_R g43003 (.A(fract_denorm[47]),
    .B(n_1625),
    .Y(n_1631));
 OAI21xp33_ASAP7_75t_R g43004 (.A1(n_1582),
    .A2(n_1619),
    .B(n_1579),
    .Y(n_1628));
 OR2x2_ASAP7_75t_R g43005 (.A(u4_n_1944),
    .B(n_1627),
    .Y(n_1630));
 OR2x2_ASAP7_75t_R g43006 (.A(n_1596),
    .B(n_1626),
    .Y(n_1629));
 NAND2xp33_ASAP7_75t_R g43007 (.A(n_1600),
    .B(n_1617),
    .Y(n_1627));
 NAND2xp33_ASAP7_75t_R g43008 (.A(n_1597),
    .B(n_1618),
    .Y(n_1626));
 INVxp33_ASAP7_75t_R g43009 (.A(n_1623),
    .Y(n_1624));
 O2A1O1Ixp33_ASAP7_75t_R g43010 (.A1(n_1594),
    .A2(fract_denorm[4]),
    .B(n_1567),
    .C(fract_denorm[6]),
    .Y(n_1622));
 NAND2xp33_ASAP7_75t_R g43011 (.A(n_1612),
    .B(n_1615),
    .Y(n_1625));
 NOR3xp33_ASAP7_75t_R g43012 (.A(n_1613),
    .B(u4_n_1938),
    .C(u4_n_1942),
    .Y(n_1623));
 NAND2xp33_ASAP7_75t_R g43013 (.A(n_1601),
    .B(n_1607),
    .Y(n_1620));
 AOI211xp5_ASAP7_75t_R g43014 (.A1(n_1581),
    .A2(n_1584),
    .B(fract_denorm[6]),
    .C(fract_denorm[5]),
    .Y(n_1619));
 NAND2xp33_ASAP7_75t_R g43015 (.A(n_1611),
    .B(n_1609),
    .Y(n_1621));
 INVxp33_ASAP7_75t_R g43016 (.A(n_1615),
    .Y(n_1616));
 NOR3xp33_ASAP7_75t_R g43017 (.A(u4_n_1934),
    .B(fract_denorm[36]),
    .C(fract_denorm[35]),
    .Y(n_1618));
 NOR4xp25_ASAP7_75t_R g43018 (.A(fract_denorm[17]),
    .B(fract_denorm[20]),
    .C(fract_denorm[19]),
    .D(fract_denorm[18]),
    .Y(n_1617));
 NOR4xp25_ASAP7_75t_R g43019 (.A(fract_denorm[44]),
    .B(fract_denorm[41]),
    .C(fract_denorm[42]),
    .D(fract_denorm[43]),
    .Y(n_1615));
 NOR2xp33_ASAP7_75t_R g43020 (.A(n_1608),
    .B(n_1601),
    .Y(n_1614));
 NAND2xp33_ASAP7_75t_R g43021 (.A(n_1605),
    .B(n_1606),
    .Y(n_1613));
 NOR2xp33_ASAP7_75t_R g43022 (.A(fract_denorm[45]),
    .B(fract_denorm[46]),
    .Y(n_1612));
 INVxp33_ASAP7_75t_R g43023 (.A(n_1609),
    .Y(n_1610));
 INVxp33_ASAP7_75t_R g43024 (.A(n_1607),
    .Y(n_1608));
 NOR4xp25_ASAP7_75t_R g43025 (.A(fract_denorm[9]),
    .B(fract_denorm[12]),
    .C(fract_denorm[11]),
    .D(fract_denorm[10]),
    .Y(n_1611));
 NOR3xp33_ASAP7_75t_R g43026 (.A(n_1580),
    .B(fract_denorm[15]),
    .C(fract_denorm[16]),
    .Y(n_1609));
 NOR3xp33_ASAP7_75t_R g43027 (.A(n_1582),
    .B(fract_denorm[5]),
    .C(fract_denorm[6]),
    .Y(n_1607));
 INVxp33_ASAP7_75t_R g43028 (.A(n_1606),
    .Y(u4_n_1948));
 INVxp33_ASAP7_75t_R g43029 (.A(n_1605),
    .Y(u4_n_1946));
 INVxp33_ASAP7_75t_R g43030 (.A(n_1604),
    .Y(u4_n_1938));
 INVxp33_ASAP7_75t_R g43031 (.A(n_1603),
    .Y(u4_n_1944));
 NOR2xp33_ASAP7_75t_R g43033 (.A(fract_denorm[27]),
    .B(fract_denorm[28]),
    .Y(n_1606));
 NOR2xp33_ASAP7_75t_R g43034 (.A(fract_denorm[25]),
    .B(fract_denorm[26]),
    .Y(n_1605));
 OR2x2_ASAP7_75t_R g43035 (.A(fract_denorm[29]),
    .B(fract_denorm[30]),
    .Y(u4_n_1942));
 NOR2xp33_ASAP7_75t_R g43036 (.A(fract_denorm[31]),
    .B(fract_denorm[32]),
    .Y(n_1604));
 NOR2xp33_ASAP7_75t_R g43037 (.A(fract_denorm[23]),
    .B(fract_denorm[24]),
    .Y(n_1603));
 INVxp33_ASAP7_75t_R g43039 (.A(n_1599),
    .Y(u4_n_1934));
 INVxp33_ASAP7_75t_R g43040 (.A(n_1597),
    .Y(n_1598));
 INVxp33_ASAP7_75t_R g43041 (.A(n_1595),
    .Y(n_1596));
 AOI21xp33_ASAP7_75t_R g43042 (.A1(n_1571),
    .A2(fract_denorm[1]),
    .B(fract_denorm[3]),
    .Y(n_1594));
 NAND2xp33_ASAP7_75t_R g43043 (.A(n_1581),
    .B(n_1583),
    .Y(n_1601));
 NOR2xp33_ASAP7_75t_R g43044 (.A(fract_denorm[41]),
    .B(fract_denorm[42]),
    .Y(n_1593));
 NOR2xp33_ASAP7_75t_R g43045 (.A(fract_denorm[20]),
    .B(fract_denorm[19]),
    .Y(n_1592));
 NOR2xp33_ASAP7_75t_R g43046 (.A(fract_denorm[22]),
    .B(fract_denorm[21]),
    .Y(n_1600));
 NOR2xp33_ASAP7_75t_R g43047 (.A(fract_denorm[33]),
    .B(fract_denorm[34]),
    .Y(n_1599));
 NOR2xp33_ASAP7_75t_R g43048 (.A(fract_denorm[37]),
    .B(fract_denorm[38]),
    .Y(n_1597));
 NOR2xp33_ASAP7_75t_R g43049 (.A(fract_denorm[39]),
    .B(fract_denorm[40]),
    .Y(n_1595));
 INVxp33_ASAP7_75t_R g43052 (.A(fract_denorm[26]),
    .Y(n_1589));
 INVxp33_ASAP7_75t_R g43055 (.A(fract_denorm[44]),
    .Y(n_1586));
 INVxp33_ASAP7_75t_R g43075 (.A(n_1583),
    .Y(n_1584));
 INVxp33_ASAP7_75t_R g43076 (.A(n_1579),
    .Y(n_1580));
 INVxp33_ASAP7_75t_R g43080 (.A(fract_denorm[47]),
    .Y(n_1575));
 NAND2xp33_ASAP7_75t_R g43081 (.A(n_1067),
    .B(n_1540),
    .Y(n_1574));
 NAND2xp33_ASAP7_75t_R g43082 (.A(n_1065),
    .B(n_1539),
    .Y(n_1573));
 NOR2xp33_ASAP7_75t_R g43083 (.A(fract_denorm[2]),
    .B(fract_denorm[1]),
    .Y(n_1583));
 OR2x2_ASAP7_75t_R g43084 (.A(fract_denorm[8]),
    .B(fract_denorm[7]),
    .Y(n_1582));
 NOR2xp33_ASAP7_75t_R g43085 (.A(fract_denorm[12]),
    .B(fract_denorm[11]),
    .Y(n_1572));
 NOR2xp33_ASAP7_75t_R g43086 (.A(fract_denorm[4]),
    .B(fract_denorm[3]),
    .Y(n_1581));
 NOR2xp33_ASAP7_75t_R g43088 (.A(fract_denorm[14]),
    .B(fract_denorm[13]),
    .Y(n_1579));
 INVxp33_ASAP7_75t_R g43099 (.A(fract_denorm[2]),
    .Y(n_1571));
 INVxp33_ASAP7_75t_R g43100 (.A(fract_denorm[11]),
    .Y(n_1570));
 NAND2xp33_ASAP7_75t_R g43104 (.A(n_1497),
    .B(n_1107),
    .Y(n_1566));
 NAND2xp33_ASAP7_75t_R g43105 (.A(n_1538),
    .B(n_1110),
    .Y(n_1565));
 NAND2xp33_ASAP7_75t_R g43106 (.A(n_1519),
    .B(n_1109),
    .Y(n_1564));
 NAND2xp33_ASAP7_75t_R g43107 (.A(n_1520),
    .B(n_1090),
    .Y(n_1563));
 NAND2xp33_ASAP7_75t_R g43108 (.A(n_1521),
    .B(n_1095),
    .Y(n_1562));
 NAND2xp33_ASAP7_75t_R g43109 (.A(n_1522),
    .B(n_1100),
    .Y(n_1561));
 NAND2xp33_ASAP7_75t_R g43110 (.A(n_1066),
    .B(n_1517),
    .Y(n_1560));
 NAND2xp33_ASAP7_75t_R g43130 (.A(n_1516),
    .B(n_1112),
    .Y(n_1559));
 NAND2xp33_ASAP7_75t_R g43131 (.A(n_1515),
    .B(n_1111),
    .Y(n_1558));
 NAND2xp33_ASAP7_75t_R g43132 (.A(n_1514),
    .B(n_1096),
    .Y(n_1557));
 NAND2xp33_ASAP7_75t_R g43133 (.A(n_1513),
    .B(n_1103),
    .Y(n_1556));
 NAND2xp33_ASAP7_75t_R g43134 (.A(n_1512),
    .B(n_1115),
    .Y(n_1555));
 NAND2xp33_ASAP7_75t_R g43135 (.A(n_1511),
    .B(n_1106),
    .Y(n_1554));
 NAND2xp33_ASAP7_75t_R g43136 (.A(n_1510),
    .B(n_1104),
    .Y(n_1553));
 NAND2xp33_ASAP7_75t_R g43137 (.A(n_1509),
    .B(n_1099),
    .Y(n_1552));
 NAND2xp33_ASAP7_75t_R g43138 (.A(n_1508),
    .B(n_1093),
    .Y(n_1551));
 NAND2xp33_ASAP7_75t_R g43139 (.A(n_1507),
    .B(n_1094),
    .Y(n_1550));
 NAND2xp33_ASAP7_75t_R g43140 (.A(n_1506),
    .B(n_1102),
    .Y(n_1549));
 NAND2xp33_ASAP7_75t_R g43141 (.A(n_1505),
    .B(n_1108),
    .Y(n_1548));
 NAND2xp33_ASAP7_75t_R g43142 (.A(n_1504),
    .B(n_1113),
    .Y(n_1547));
 NAND2xp33_ASAP7_75t_R g43143 (.A(n_1503),
    .B(n_1114),
    .Y(n_1546));
 NAND2xp33_ASAP7_75t_R g43144 (.A(n_1502),
    .B(n_1097),
    .Y(n_1545));
 NAND2xp33_ASAP7_75t_R g43145 (.A(n_1501),
    .B(n_1105),
    .Y(n_1544));
 NAND2xp33_ASAP7_75t_R g43146 (.A(n_1500),
    .B(n_1092),
    .Y(n_1543));
 NAND2xp33_ASAP7_75t_R g43147 (.A(n_1499),
    .B(n_1091),
    .Y(n_1542));
 NAND2xp33_ASAP7_75t_R g43148 (.A(n_1498),
    .B(n_1101),
    .Y(n_1541));
 AOI222xp33_ASAP7_75t_R g43152 (.A1(n_681),
    .A2(fract_i2f[43]),
    .B1(n_1059),
    .B2(quo[45]),
    .C1(n_1060),
    .C2(quo[22]),
    .Y(n_1540));
 AOI222xp33_ASAP7_75t_R g43153 (.A1(n_681),
    .A2(fract_i2f[45]),
    .B1(n_676),
    .B2(quo[47]),
    .C1(n_1060),
    .C2(quo[24]),
    .Y(n_1539));
 AOI22xp33_ASAP7_75t_R g43154 (.A1(fract_i2f[25]),
    .A2(n_682),
    .B1(prod[25]),
    .B2(n_674),
    .Y(n_1538));
 AO222x2_ASAP7_75t_R g43155 (.A1(n_681),
    .A2(fract_i2f[7]),
    .B1(n_671),
    .B2(prod[7]),
    .C1(quo[9]),
    .C2(n_1059),
    .Y(n_1537));
 AO222x2_ASAP7_75t_R g43156 (.A1(n_682),
    .A2(fract_i2f[8]),
    .B1(n_674),
    .B2(prod[8]),
    .C1(quo[10]),
    .C2(n_1059),
    .Y(n_1536));
 AO222x2_ASAP7_75t_R g43157 (.A1(n_680),
    .A2(fract_i2f[9]),
    .B1(n_671),
    .B2(prod[9]),
    .C1(quo[11]),
    .C2(n_1059),
    .Y(n_1535));
 AO222x2_ASAP7_75t_R g43158 (.A1(n_679),
    .A2(fract_i2f[10]),
    .B1(n_671),
    .B2(prod[10]),
    .C1(quo[12]),
    .C2(n_677),
    .Y(n_1534));
 AO222x2_ASAP7_75t_R g43159 (.A1(n_681),
    .A2(fract_i2f[11]),
    .B1(n_672),
    .B2(prod[11]),
    .C1(quo[13]),
    .C2(n_676),
    .Y(n_1533));
 AO222x2_ASAP7_75t_R g43160 (.A1(n_680),
    .A2(fract_i2f[12]),
    .B1(n_674),
    .B2(prod[12]),
    .C1(quo[14]),
    .C2(n_678),
    .Y(n_1532));
 AO222x2_ASAP7_75t_R g43161 (.A1(n_681),
    .A2(fract_i2f[13]),
    .B1(n_674),
    .B2(prod[13]),
    .C1(quo[15]),
    .C2(n_676),
    .Y(n_1531));
 AO222x2_ASAP7_75t_R g43162 (.A1(n_682),
    .A2(fract_i2f[14]),
    .B1(n_671),
    .B2(prod[14]),
    .C1(quo[16]),
    .C2(n_677),
    .Y(n_1530));
 AO222x2_ASAP7_75t_R g43163 (.A1(n_681),
    .A2(fract_i2f[15]),
    .B1(n_671),
    .B2(prod[15]),
    .C1(quo[17]),
    .C2(n_676),
    .Y(n_1529));
 AO222x2_ASAP7_75t_R g43164 (.A1(n_679),
    .A2(fract_i2f[16]),
    .B1(n_674),
    .B2(prod[16]),
    .C1(quo[18]),
    .C2(n_1059),
    .Y(n_1528));
 AO222x2_ASAP7_75t_R g43165 (.A1(n_680),
    .A2(fract_i2f[1]),
    .B1(n_23),
    .B2(prod[1]),
    .C1(quo[3]),
    .C2(n_676),
    .Y(n_1527));
 AO222x2_ASAP7_75t_R g43166 (.A1(n_682),
    .A2(fract_i2f[2]),
    .B1(n_23),
    .B2(prod[2]),
    .C1(quo[4]),
    .C2(n_677),
    .Y(n_1526));
 AO222x2_ASAP7_75t_R g43167 (.A1(n_682),
    .A2(fract_i2f[3]),
    .B1(n_672),
    .B2(prod[3]),
    .C1(quo[5]),
    .C2(n_678),
    .Y(n_1525));
 AO222x2_ASAP7_75t_R g43168 (.A1(n_679),
    .A2(fract_i2f[4]),
    .B1(n_23),
    .B2(prod[4]),
    .C1(quo[6]),
    .C2(n_676),
    .Y(n_1524));
 AO222x2_ASAP7_75t_R g43169 (.A1(n_680),
    .A2(fract_i2f[5]),
    .B1(n_672),
    .B2(prod[5]),
    .C1(quo[7]),
    .C2(n_677),
    .Y(n_1523));
 AOI22xp33_ASAP7_75t_R g43170 (.A1(fract_i2f[21]),
    .A2(n_682),
    .B1(prod[21]),
    .B2(n_671),
    .Y(n_1522));
 AOI22xp33_ASAP7_75t_R g43171 (.A1(fract_i2f[22]),
    .A2(n_679),
    .B1(prod[22]),
    .B2(n_23),
    .Y(n_1521));
 AOI22xp33_ASAP7_75t_R g43172 (.A1(fract_i2f[23]),
    .A2(n_680),
    .B1(prod[23]),
    .B2(n_674),
    .Y(n_1520));
 AOI22xp33_ASAP7_75t_R g43173 (.A1(fract_i2f[24]),
    .A2(n_682),
    .B1(prod[24]),
    .B2(n_672),
    .Y(n_1519));
 AO222x2_ASAP7_75t_R g43174 (.A1(n_679),
    .A2(fract_i2f[6]),
    .B1(n_672),
    .B2(prod[6]),
    .C1(quo[8]),
    .C2(n_678),
    .Y(n_1518));
 AOI22xp33_ASAP7_75t_R g43175 (.A1(fract_i2f[20]),
    .A2(n_680),
    .B1(quo[22]),
    .B2(n_677),
    .Y(n_1517));
 AOI22xp33_ASAP7_75t_R g43176 (.A1(fract_i2f[27]),
    .A2(n_681),
    .B1(prod[27]),
    .B2(n_671),
    .Y(n_1516));
 AOI22xp33_ASAP7_75t_R g43177 (.A1(fract_i2f[28]),
    .A2(n_682),
    .B1(prod[28]),
    .B2(n_23),
    .Y(n_1515));
 AOI22xp33_ASAP7_75t_R g43178 (.A1(fract_i2f[29]),
    .A2(n_682),
    .B1(prod[29]),
    .B2(n_671),
    .Y(n_1514));
 AOI22xp33_ASAP7_75t_R g43179 (.A1(fract_i2f[30]),
    .A2(n_680),
    .B1(prod[30]),
    .B2(n_672),
    .Y(n_1513));
 AOI22xp33_ASAP7_75t_R g43180 (.A1(fract_i2f[31]),
    .A2(n_681),
    .B1(prod[31]),
    .B2(n_672),
    .Y(n_1512));
 AOI22xp33_ASAP7_75t_R g43181 (.A1(fract_i2f[32]),
    .A2(n_679),
    .B1(prod[32]),
    .B2(n_672),
    .Y(n_1511));
 AOI22xp33_ASAP7_75t_R g43182 (.A1(fract_i2f[33]),
    .A2(n_681),
    .B1(prod[33]),
    .B2(n_23),
    .Y(n_1510));
 AOI22xp33_ASAP7_75t_R g43183 (.A1(fract_i2f[34]),
    .A2(n_679),
    .B1(prod[34]),
    .B2(n_672),
    .Y(n_1509));
 AOI22xp33_ASAP7_75t_R g43184 (.A1(fract_i2f[35]),
    .A2(n_681),
    .B1(prod[35]),
    .B2(n_23),
    .Y(n_1508));
 AOI22xp33_ASAP7_75t_R g43185 (.A1(fract_i2f[36]),
    .A2(n_680),
    .B1(prod[36]),
    .B2(n_23),
    .Y(n_1507));
 AOI22xp33_ASAP7_75t_R g43186 (.A1(fract_i2f[37]),
    .A2(n_679),
    .B1(prod[37]),
    .B2(n_674),
    .Y(n_1506));
 AOI22xp33_ASAP7_75t_R g43187 (.A1(fract_i2f[38]),
    .A2(n_682),
    .B1(prod[38]),
    .B2(n_23),
    .Y(n_1505));
 AOI22xp33_ASAP7_75t_R g43188 (.A1(fract_i2f[39]),
    .A2(n_679),
    .B1(prod[39]),
    .B2(n_674),
    .Y(n_1504));
 AOI22xp33_ASAP7_75t_R g43189 (.A1(fract_i2f[40]),
    .A2(n_679),
    .B1(prod[40]),
    .B2(n_23),
    .Y(n_1503));
 AOI22xp33_ASAP7_75t_R g43190 (.A1(fract_i2f[41]),
    .A2(n_680),
    .B1(prod[41]),
    .B2(n_672),
    .Y(n_1502));
 AOI22xp33_ASAP7_75t_R g43191 (.A1(fract_i2f[42]),
    .A2(n_681),
    .B1(prod[42]),
    .B2(n_671),
    .Y(n_1501));
 AOI22xp33_ASAP7_75t_R g43192 (.A1(fract_i2f[44]),
    .A2(n_680),
    .B1(prod[44]),
    .B2(n_23),
    .Y(n_1500));
 AOI22xp33_ASAP7_75t_R g43193 (.A1(fract_i2f[46]),
    .A2(n_681),
    .B1(prod[46]),
    .B2(n_674),
    .Y(n_1499));
 AOI22xp33_ASAP7_75t_R g43194 (.A1(fract_i2f[47]),
    .A2(n_679),
    .B1(prod[47]),
    .B2(n_674),
    .Y(n_1498));
 AOI22xp33_ASAP7_75t_R g43195 (.A1(fract_i2f[26]),
    .A2(n_682),
    .B1(prod[26]),
    .B2(n_672),
    .Y(n_1497));
 NOR2xp33_ASAP7_75t_R g43243 (.A(n_774),
    .B(sign),
    .Y(u4_n_1446));
 AOI221xp5_ASAP7_75t_R g43244 (.A1(n_667),
    .A2(opa_r1[7]),
    .B1(n_3833),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1496));
 AOI221xp5_ASAP7_75t_R g43245 (.A1(n_667),
    .A2(opa_r1[8]),
    .B1(n_3834),
    .B2(n_1432),
    .C(n_1443),
    .Y(n_1495));
 AOI221xp5_ASAP7_75t_R g43246 (.A1(n_1433),
    .A2(opa_r1[9]),
    .B1(n_3835),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1494));
 AOI221xp5_ASAP7_75t_R g43247 (.A1(n_667),
    .A2(opa_r1[10]),
    .B1(n_3836),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1493));
 AOI221xp5_ASAP7_75t_R g43248 (.A1(n_667),
    .A2(opa_r1[11]),
    .B1(n_3837),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1492));
 AOI221xp5_ASAP7_75t_R g43249 (.A1(n_667),
    .A2(opa_r1[12]),
    .B1(n_3648),
    .B2(n_669),
    .C(n_662),
    .Y(n_1491));
 AOI221xp5_ASAP7_75t_R g43250 (.A1(n_1433),
    .A2(opa_r1[13]),
    .B1(n_3649),
    .B2(n_1432),
    .C(n_1443),
    .Y(n_1490));
 AOI221xp5_ASAP7_75t_R g43251 (.A1(n_1433),
    .A2(opa_r1[14]),
    .B1(n_3650),
    .B2(n_1432),
    .C(n_1443),
    .Y(n_1489));
 AOI221xp5_ASAP7_75t_R g43252 (.A1(n_1433),
    .A2(opa_r1[15]),
    .B1(n_3651),
    .B2(n_1432),
    .C(n_1443),
    .Y(n_1488));
 AOI221xp5_ASAP7_75t_R g43253 (.A1(n_1433),
    .A2(opa_r1[16]),
    .B1(n_3652),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1487));
 AOI221xp5_ASAP7_75t_R g43254 (.A1(n_1433),
    .A2(opa_r1[17]),
    .B1(n_3653),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1486));
 AOI221xp5_ASAP7_75t_R g43255 (.A1(n_667),
    .A2(opa_r1[18]),
    .B1(n_3654),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1485));
 AOI221xp5_ASAP7_75t_R g43256 (.A1(n_667),
    .A2(opa_r1[19]),
    .B1(n_3655),
    .B2(n_669),
    .C(n_662),
    .Y(n_1484));
 AOI221xp5_ASAP7_75t_R g43257 (.A1(n_1433),
    .A2(opa_r1[20]),
    .B1(n_3656),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1483));
 AOI221xp5_ASAP7_75t_R g43258 (.A1(n_1433),
    .A2(opa_r1[21]),
    .B1(n_3657),
    .B2(n_669),
    .C(n_662),
    .Y(n_1482));
 AOI221xp5_ASAP7_75t_R g43259 (.A1(n_1433),
    .A2(opa_r1[22]),
    .B1(n_3658),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1481));
 AOI221xp5_ASAP7_75t_R g43260 (.A1(n_1433),
    .A2(opa_r1[23]),
    .B1(n_3659),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1480));
 AOI221xp5_ASAP7_75t_R g43261 (.A1(n_667),
    .A2(opa_r1[24]),
    .B1(n_3660),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1479));
 AOI221xp5_ASAP7_75t_R g43262 (.A1(n_667),
    .A2(opa_r1[25]),
    .B1(n_3661),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1478));
 AOI221xp5_ASAP7_75t_R g43263 (.A1(n_667),
    .A2(opa_r1[26]),
    .B1(n_3662),
    .B2(n_669),
    .C(n_1443),
    .Y(n_1477));
 AOI221xp5_ASAP7_75t_R g43264 (.A1(n_667),
    .A2(opa_r1[27]),
    .B1(n_3663),
    .B2(n_1432),
    .C(n_662),
    .Y(n_1476));
 AOI221xp5_ASAP7_75t_R g43265 (.A1(n_667),
    .A2(opa_r1[28]),
    .B1(n_3664),
    .B2(n_1432),
    .C(n_1443),
    .Y(n_1475));
 AOI221xp5_ASAP7_75t_R g43266 (.A1(n_1433),
    .A2(opa_r1[29]),
    .B1(n_3665),
    .B2(n_669),
    .C(n_662),
    .Y(n_1474));
 AOI221xp5_ASAP7_75t_R g43267 (.A1(n_1433),
    .A2(opa_r1[30]),
    .B1(n_3666),
    .B2(n_669),
    .C(n_662),
    .Y(n_1473));
 AOI221xp5_ASAP7_75t_R g43268 (.A1(n_1436),
    .A2(opa_r1[18]),
    .B1(n_1433),
    .B2(opa_r1[1]),
    .C(n_1455),
    .Y(n_1472));
 AOI221xp5_ASAP7_75t_R g43269 (.A1(n_659),
    .A2(opa_r1[21]),
    .B1(n_1433),
    .B2(opa_r1[4]),
    .C(n_1447),
    .Y(n_1471));
 AOI221xp5_ASAP7_75t_R g43270 (.A1(n_659),
    .A2(opa_r1[19]),
    .B1(n_667),
    .B2(opa_r1[2]),
    .C(n_1448),
    .Y(n_1470));
 AOI221xp5_ASAP7_75t_R g43271 (.A1(n_1436),
    .A2(opa_r1[20]),
    .B1(n_667),
    .B2(opa_r1[3]),
    .C(n_1461),
    .Y(n_1469));
 AOI221xp5_ASAP7_75t_R g43272 (.A1(n_659),
    .A2(opa_r1[22]),
    .B1(n_1433),
    .B2(opa_r1[5]),
    .C(n_1446),
    .Y(n_1468));
 AOI221xp5_ASAP7_75t_R g43273 (.A1(n_667),
    .A2(opa_r1[6]),
    .B1(n_3832),
    .B2(n_669),
    .C(n_1445),
    .Y(n_1467));
 AOI221xp5_ASAP7_75t_R g43274 (.A1(n_1436),
    .A2(opa_r1[17]),
    .B1(n_3499),
    .B2(opa_r1[0]),
    .C(n_1442),
    .Y(n_1466));
 AOI22xp33_ASAP7_75t_R g43275 (.A1(n_1435),
    .A2(n_1063),
    .B1(opa_r1[5]),
    .B2(n_659),
    .Y(n_1465));
 AOI22xp33_ASAP7_75t_R g43276 (.A1(n_1007),
    .A2(n_655),
    .B1(opa_r1[2]),
    .B2(n_659),
    .Y(n_1464));
 AOI22xp33_ASAP7_75t_R g43277 (.A1(n_1026),
    .A2(n_1435),
    .B1(opa_r1[3]),
    .B2(n_659),
    .Y(n_1463));
 AOI22xp33_ASAP7_75t_R g43278 (.A1(n_640),
    .A2(n_1435),
    .B1(opa_r1[4]),
    .B2(n_659),
    .Y(n_1462));
 AO21x1_ASAP7_75t_R g43279 (.A1(n_3829),
    .A2(n_1432),
    .B(n_1439),
    .Y(n_1461));
 AOI22xp33_ASAP7_75t_R g43280 (.A1(n_655),
    .A2(n_644),
    .B1(opa_r1[10]),
    .B2(n_659),
    .Y(n_1460));
 AOI22xp33_ASAP7_75t_R g43281 (.A1(n_1435),
    .A2(n_642),
    .B1(opa_r1[6]),
    .B2(n_659),
    .Y(n_1459));
 AOI22xp33_ASAP7_75t_R g43282 (.A1(n_1435),
    .A2(n_1089),
    .B1(opa_r1[7]),
    .B2(n_1436),
    .Y(n_1458));
 AOI22xp33_ASAP7_75t_R g43283 (.A1(n_1435),
    .A2(n_643),
    .B1(opa_r1[8]),
    .B2(n_1436),
    .Y(n_1457));
 AOI22xp33_ASAP7_75t_R g43284 (.A1(n_1435),
    .A2(n_1135),
    .B1(opa_r1[9]),
    .B2(n_1436),
    .Y(n_1456));
 AO21x1_ASAP7_75t_R g43286 (.A1(n_3827),
    .A2(n_669),
    .B(n_1441),
    .Y(n_1455));
 AOI22xp33_ASAP7_75t_R g43287 (.A1(n_1435),
    .A2(n_645),
    .B1(opa_r1[12]),
    .B2(n_1436),
    .Y(n_1454));
 AOI22xp33_ASAP7_75t_R g43288 (.A1(n_1435),
    .A2(n_1149),
    .B1(opa_r1[13]),
    .B2(n_1436),
    .Y(n_1453));
 AOI22xp33_ASAP7_75t_R g43289 (.A1(n_1435),
    .A2(n_647),
    .B1(opa_r1[14]),
    .B2(n_1436),
    .Y(n_1452));
 AOI22xp33_ASAP7_75t_R g43290 (.A1(n_1435),
    .A2(n_1160),
    .B1(opa_r1[15]),
    .B2(n_659),
    .Y(n_1451));
 AOI22xp33_ASAP7_75t_R g43291 (.A1(n_1435),
    .A2(n_648),
    .B1(opa_r1[16]),
    .B2(n_659),
    .Y(n_1450));
 AOI22xp33_ASAP7_75t_R g43292 (.A1(n_1435),
    .A2(n_1143),
    .B1(opa_r1[11]),
    .B2(n_659),
    .Y(n_1449));
 AO21x1_ASAP7_75t_R g43293 (.A1(n_3828),
    .A2(n_1432),
    .B(n_1438),
    .Y(n_1448));
 AO21x1_ASAP7_75t_R g43294 (.A1(n_1432),
    .A2(n_3830),
    .B(n_1440),
    .Y(n_1447));
 AO21x1_ASAP7_75t_R g43295 (.A1(n_669),
    .A2(n_3831),
    .B(n_1437),
    .Y(n_1446));
 OAI22xp33_ASAP7_75t_R g43296 (.A1(n_1434),
    .A2(n_1264),
    .B1(n_1077),
    .B2(n_699),
    .Y(n_1445));
 AOI22xp33_ASAP7_75t_R g43297 (.A1(n_988),
    .A2(n_1435),
    .B1(opa_r1[1]),
    .B2(n_1436),
    .Y(n_1444));
 O2A1O1Ixp33_ASAP7_75t_R g43298 (.A1(opa_r1[17]),
    .A2(n_1193),
    .B(n_1196),
    .C(n_1434),
    .Y(n_1442));
 O2A1O1Ixp33_ASAP7_75t_R g43299 (.A1(opa_r1[18]),
    .A2(n_1200),
    .B(n_1213),
    .C(n_1434),
    .Y(n_1441));
 AOI21xp33_ASAP7_75t_R g43300 (.A1(n_1261),
    .A2(n_1077),
    .B(n_1434),
    .Y(n_1443));
 O2A1O1Ixp33_ASAP7_75t_R g43301 (.A1(opa_r1[21]),
    .A2(n_1231),
    .B(n_1244),
    .C(n_1434),
    .Y(n_1440));
 O2A1O1Ixp33_ASAP7_75t_R g43302 (.A1(opa_r1[20]),
    .A2(n_1223),
    .B(n_1230),
    .C(n_1434),
    .Y(n_1439));
 O2A1O1Ixp33_ASAP7_75t_R g43303 (.A1(opa_r1[19]),
    .A2(n_1214),
    .B(n_1221),
    .C(n_1434),
    .Y(n_1438));
 O2A1O1Ixp33_ASAP7_75t_R g43304 (.A1(opa_r1[22]),
    .A2(n_1246),
    .B(n_1262),
    .C(n_1434),
    .Y(n_1437));
 INVxp33_ASAP7_75t_R g43306 (.A(n_1435),
    .Y(n_1434));
 NOR2xp33_ASAP7_75t_R g43307 (.A(n_1430),
    .B(n_3499),
    .Y(n_1436));
 NOR2xp33_ASAP7_75t_R g43308 (.A(n_1431),
    .B(n_3499),
    .Y(n_1435));
 NOR2xp33_ASAP7_75t_R g43309 (.A(n_621),
    .B(n_1430),
    .Y(n_1433));
 NOR2xp33_ASAP7_75t_R g43310 (.A(n_621),
    .B(n_1431),
    .Y(n_1432));
 INVxp33_ASAP7_75t_R g43311 (.A(n_1431),
    .Y(n_1430));
 AOI22xp33_ASAP7_75t_R g43312 (.A1(sign_fasu),
    .A2(n_801),
    .B1(sign_mul),
    .B2(fpu_op_r2[1]),
    .Y(n_1431));
 AOI22xp33_ASAP7_75t_R g43314 (.A1(u1_n_5382),
    .A2(n_9),
    .B1(opa_r[31]),
    .B2(u1_n_1066),
    .Y(n_1429));
 NAND2xp33_ASAP7_75t_R g43316 (.A(n_687),
    .B(n_1427),
    .Y(u1_n_1066));
 AOI322xp5_ASAP7_75t_R g43317 (.A1(n_1426),
    .A2(n_1406),
    .A3(n_1399),
    .B1(n_1345),
    .B2(n_1388),
    .C1(n_1421),
    .C2(n_1399),
    .Y(n_1427));
 AOI221xp5_ASAP7_75t_R g43318 (.A1(u1_n_1048),
    .A2(n_1378),
    .B1(n_1425),
    .B2(n_1415),
    .C(n_1402),
    .Y(n_1426));
 OAI221xp5_ASAP7_75t_R g43319 (.A1(u1_n_1022),
    .A2(n_1371),
    .B1(u1_n_1023),
    .B2(n_1382),
    .C(n_1424),
    .Y(n_1425));
 MAJIxp5_ASAP7_75t_R g43320 (.A(n_1423),
    .B(n_1383),
    .C(u1_n_1051),
    .Y(n_1424));
 MAJIxp5_ASAP7_75t_R g43321 (.A(n_1422),
    .B(n_1396),
    .C(u1_n_1025),
    .Y(n_1423));
 OAI322xp33_ASAP7_75t_R g43322 (.A1(n_1419),
    .A2(n_1416),
    .A3(n_1404),
    .B1(n_1416),
    .B2(n_1409),
    .C1(n_1397),
    .C2(n_1408),
    .Y(n_1422));
 OAI21xp33_ASAP7_75t_R g43323 (.A1(u1_n_1041),
    .A2(n_1341),
    .B(n_1420),
    .Y(n_1421));
 AOI322xp5_ASAP7_75t_R g43324 (.A1(n_1361),
    .A2(n_1354),
    .A3(u1_n_1015),
    .B1(n_1406),
    .B2(n_14518),
    .C1(n_1384),
    .C2(n_1400),
    .Y(n_1420));
 AOI321xp33_ASAP7_75t_R g43325 (.A1(n_1407),
    .A2(u1_n_1031),
    .A3(n_1391),
    .B1(u1_n_1030),
    .B2(n_1392),
    .C(n_13843),
    .Y(n_1419));
 A2O1A1Ixp33_ASAP7_75t_R g43328 (.A1(n_1382),
    .A2(u1_n_1023),
    .B(u1_n_1022),
    .C(n_1410),
    .Y(n_1415));
 OAI221xp5_ASAP7_75t_R g43330 (.A1(n_1394),
    .A2(u1_n_1028),
    .B1(n_1395),
    .B2(u1_n_1027),
    .C(n_1398),
    .Y(n_1416));
 AOI22xp33_ASAP7_75t_R g43331 (.A1(n_1389),
    .A2(u1_n_1032),
    .B1(u1_n_1033),
    .B2(n_1405),
    .Y(n_1412));
 OAI22xp33_ASAP7_75t_R g43332 (.A1(u1_n_1034),
    .A2(n_1403),
    .B1(n_1405),
    .B2(u1_n_1033),
    .Y(n_1411));
 OAI221xp5_ASAP7_75t_R g43333 (.A1(n_1391),
    .A2(u1_n_1031),
    .B1(n_1389),
    .B2(u1_n_1032),
    .C(n_1407),
    .Y(n_1413));
 OAI31xp33_ASAP7_75t_R g43334 (.A1(n_1377),
    .A2(u1_n_1050),
    .A3(n_1370),
    .B(u1_n_1049),
    .Y(n_1410));
 AOI22xp33_ASAP7_75t_R g43335 (.A1(u1_n_1028),
    .A2(n_1394),
    .B1(u1_n_1029),
    .B2(n_1393),
    .Y(n_1409));
 AOI22xp33_ASAP7_75t_R g43336 (.A1(n_1395),
    .A2(u1_n_1027),
    .B1(u1_n_1026),
    .B2(n_1379),
    .Y(n_1408));
 INVxp33_ASAP7_75t_R g43337 (.A(n_1405),
    .Y(u1_n_1060));
 NOR2xp33_ASAP7_75t_R g43338 (.A(n_1393),
    .B(u1_n_1029),
    .Y(n_1404));
 NAND2xp33_ASAP7_75t_R g43339 (.A(u1_n_1057),
    .B(n_1390),
    .Y(n_1407));
 OA211x2_ASAP7_75t_R g43340 (.A1(n_1366),
    .A2(u1_n_1017),
    .B(n_1384),
    .C(n_1376),
    .Y(n_1406));
 AO22x1_ASAP7_75t_R g43341 (.A1(n_689),
    .A2(n_1386),
    .B1(n_1150),
    .B2(u5_mul_69_18_n_118),
    .Y(u1_n_1034));
 AOI22xp33_ASAP7_75t_R g43342 (.A1(n_1150),
    .A2(n_1385),
    .B1(n_689),
    .B2(n_14124),
    .Y(n_1405));
 INVxp33_ASAP7_75t_R g43343 (.A(n_1403),
    .Y(u1_n_1061));
 AOI22xp33_ASAP7_75t_R g43344 (.A1(u1_n_1020),
    .A2(n_1380),
    .B1(u1_n_1021),
    .B2(n_1381),
    .Y(n_1401));
 AO32x1_ASAP7_75t_R g43345 (.A1(n_1376),
    .A2(n_1366),
    .A3(u1_n_1017),
    .B1(u1_n_1016),
    .B2(n_1353),
    .Y(n_1400));
 AOI22xp33_ASAP7_75t_R g43346 (.A1(n_1150),
    .A2(n_1386),
    .B1(n_689),
    .B2(n_3303),
    .Y(n_1403));
 OAI222xp33_ASAP7_75t_R g43347 (.A1(n_1380),
    .A2(u1_n_1020),
    .B1(n_1365),
    .B2(u1_n_1019),
    .C1(n_1352),
    .C2(u1_n_1018),
    .Y(n_1402));
 AO22x1_ASAP7_75t_R g43348 (.A1(n_689),
    .A2(n_1385),
    .B1(n_1150),
    .B2(n_3436),
    .Y(u1_n_1033));
 INVxp33_ASAP7_75t_R g43349 (.A(n_1397),
    .Y(n_1398));
 INVxp33_ASAP7_75t_R g43350 (.A(n_1396),
    .Y(u1_n_1052));
 INVxp33_ASAP7_75t_R g43351 (.A(n_1395),
    .Y(u1_n_1054));
 INVxp33_ASAP7_75t_R g43352 (.A(n_1394),
    .Y(u1_n_1055));
 INVxp33_ASAP7_75t_R g43353 (.A(n_1393),
    .Y(u1_n_1056));
 INVxp33_ASAP7_75t_R g43354 (.A(n_1392),
    .Y(u1_n_1057));
 INVxp33_ASAP7_75t_R g43355 (.A(n_1391),
    .Y(u1_n_1058));
 OA211x2_ASAP7_75t_R g43356 (.A1(n_1351),
    .A2(u1_n_1013),
    .B(n_1345),
    .C(n_1340),
    .Y(n_1399));
 NOR2xp33_ASAP7_75t_R g43357 (.A(u1_n_1026),
    .B(n_1379),
    .Y(n_1397));
 AOI22xp33_ASAP7_75t_R g43358 (.A1(n_686),
    .A2(n_1373),
    .B1(n_687),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(n_1396));
 AOI22xp33_ASAP7_75t_R g43359 (.A1(n_686),
    .A2(n_1372),
    .B1(n_688),
    .B2(n_14134),
    .Y(n_1395));
 AOI22xp33_ASAP7_75t_R g43360 (.A1(n_1375),
    .A2(n_663),
    .B1(n_14132),
    .B2(n_688),
    .Y(n_1394));
 AOI22xp33_ASAP7_75t_R g43361 (.A1(n_663),
    .A2(n_1368),
    .B1(n_688),
    .B2(n_14130),
    .Y(n_1393));
 AOI22xp33_ASAP7_75t_R g43362 (.A1(n_1150),
    .A2(n_1369),
    .B1(n_689),
    .B2(n_14128),
    .Y(n_1392));
 AOI22xp33_ASAP7_75t_R g43363 (.A1(n_1150),
    .A2(n_1374),
    .B1(n_689),
    .B2(n_14126),
    .Y(n_1391));
 INVxp33_ASAP7_75t_R g43364 (.A(n_1390),
    .Y(u1_n_1030));
 INVxp33_ASAP7_75t_R g43365 (.A(n_1389),
    .Y(u1_n_1059));
 AO32x1_ASAP7_75t_R g43366 (.A1(n_1340),
    .A2(n_1351),
    .A3(u1_n_1013),
    .B1(n_1319),
    .B2(u1_n_1012),
    .Y(n_1388));
 AO22x1_ASAP7_75t_R g43367 (.A1(n_689),
    .A2(n_1367),
    .B1(n_1150),
    .B2(n_3427),
    .Y(u1_n_1032));
 AO22x1_ASAP7_75t_R g43368 (.A1(n_689),
    .A2(n_1375),
    .B1(n_686),
    .B2(n_3409),
    .Y(u1_n_1028));
 AOI22xp33_ASAP7_75t_R g43369 (.A1(n_689),
    .A2(n_1369),
    .B1(n_1150),
    .B2(n_3440),
    .Y(n_1390));
 AO22x1_ASAP7_75t_R g43370 (.A1(n_689),
    .A2(n_1374),
    .B1(n_1150),
    .B2(n_3411),
    .Y(u1_n_1031));
 AO22x1_ASAP7_75t_R g43371 (.A1(n_688),
    .A2(n_1368),
    .B1(n_663),
    .B2(n_3395),
    .Y(u1_n_1029));
 AO22x1_ASAP7_75t_R g43372 (.A1(n_687),
    .A2(n_1373),
    .B1(n_686),
    .B2(n_3438),
    .Y(u1_n_1025));
 AOI22xp33_ASAP7_75t_R g43373 (.A1(n_1150),
    .A2(n_1367),
    .B1(n_689),
    .B2(n_14178),
    .Y(n_1389));
 AO22x1_ASAP7_75t_R g43374 (.A1(n_689),
    .A2(n_1372),
    .B1(n_663),
    .B2(n_3434),
    .Y(u1_n_1027));
 INVxp33_ASAP7_75t_R g43375 (.A(n_1383),
    .Y(u1_n_1024));
 INVxp33_ASAP7_75t_R g43376 (.A(n_1382),
    .Y(u1_n_1050));
 NAND2xp33_ASAP7_75t_R g43377 (.A(u1_n_1019),
    .B(n_1365),
    .Y(n_1387));
 OAI221xp5_ASAP7_75t_R g43378 (.A1(n_1303),
    .A2(u1_n_1593),
    .B1(n_1335),
    .B2(n_1284),
    .C(n_1363),
    .Y(n_1386));
 OAI221xp5_ASAP7_75t_R g43379 (.A1(n_1304),
    .A2(u1_n_1593),
    .B1(n_1334),
    .B2(u1_n_1594),
    .C(n_1364),
    .Y(n_1385));
 OA21x2_ASAP7_75t_R g43380 (.A1(n_1354),
    .A2(u1_n_1015),
    .B(n_1361),
    .Y(n_1384));
 AOI22xp33_ASAP7_75t_R g43381 (.A1(n_687),
    .A2(n_1362),
    .B1(n_660),
    .B2(n_3432),
    .Y(n_1383));
 AOI22xp33_ASAP7_75t_R g43382 (.A1(n_660),
    .A2(n_1360),
    .B1(n_687),
    .B2(n_14142),
    .Y(n_1382));
 INVxp33_ASAP7_75t_R g43383 (.A(n_1381),
    .Y(u1_n_1048));
 INVxp33_ASAP7_75t_R g43384 (.A(n_1380),
    .Y(u1_n_1047));
 INVxp33_ASAP7_75t_R g43385 (.A(n_1379),
    .Y(u1_n_1053));
 INVxp33_ASAP7_75t_R g43386 (.A(n_1378),
    .Y(u1_n_1021));
 INVxp33_ASAP7_75t_R g43387 (.A(n_1377),
    .Y(u1_n_1023));
 AO22x1_ASAP7_75t_R g43388 (.A1(n_686),
    .A2(n_1362),
    .B1(n_687),
    .B2(n_14140),
    .Y(u1_n_1051));
 AOI22xp33_ASAP7_75t_R g43389 (.A1(u1_n_921),
    .A2(n_1281),
    .B1(n_14146),
    .B2(n_688),
    .Y(n_1381));
 AO22x1_ASAP7_75t_R g43390 (.A1(n_1279),
    .A2(u1_n_915),
    .B1(n_663),
    .B2(n_3415),
    .Y(u1_n_1020));
 AOI22xp33_ASAP7_75t_R g43391 (.A1(u1_n_915),
    .A2(n_1281),
    .B1(n_14148),
    .B2(n_688),
    .Y(n_1380));
 AOI322xp5_ASAP7_75t_R g43392 (.A1(n_1336),
    .A2(n_94),
    .A3(n_1150),
    .B1(n_1292),
    .B2(n_1338),
    .C1(n_14136),
    .C2(n_689),
    .Y(n_1379));
 AOI22xp33_ASAP7_75t_R g43393 (.A1(n_1279),
    .A2(u1_n_921),
    .B1(n_686),
    .B2(n_3476),
    .Y(n_1378));
 AOI22xp33_ASAP7_75t_R g43394 (.A1(n_687),
    .A2(n_1360),
    .B1(n_660),
    .B2(n_3468),
    .Y(n_1377));
 INVxp33_ASAP7_75t_R g43395 (.A(n_1371),
    .Y(u1_n_1049));
 INVxp33_ASAP7_75t_R g43396 (.A(n_1370),
    .Y(u1_n_1022));
 NAND2xp33_ASAP7_75t_R g43397 (.A(u1_n_1043),
    .B(n_1350),
    .Y(n_1376));
 OAI221xp5_ASAP7_75t_R g43398 (.A1(u1_n_1592),
    .A2(n_58),
    .B1(u1_n_1593),
    .B2(n_1298),
    .C(n_1358),
    .Y(n_1375));
 OAI221xp5_ASAP7_75t_R g43399 (.A1(n_1332),
    .A2(n_1284),
    .B1(n_1305),
    .B2(u1_n_1593),
    .C(n_1356),
    .Y(n_1374));
 OAI221xp5_ASAP7_75t_R g43400 (.A1(u1_n_1592),
    .A2(n_1300),
    .B1(u1_n_1593),
    .B2(n_1299),
    .C(n_1357),
    .Y(n_1373));
 OAI221xp5_ASAP7_75t_R g43401 (.A1(n_1309),
    .A2(u1_n_4917),
    .B1(n_1325),
    .B2(n_1275),
    .C(n_1346),
    .Y(n_1372));
 AOI22xp33_ASAP7_75t_R g43402 (.A1(n_686),
    .A2(n_1342),
    .B1(n_687),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .Y(n_1371));
 OAI31xp33_ASAP7_75t_R g43403 (.A1(n_1335),
    .A2(u1_n_1594),
    .A3(n_1150),
    .B(n_1347),
    .Y(u1_n_1026));
 AOI22xp33_ASAP7_75t_R g43404 (.A1(n_687),
    .A2(n_1342),
    .B1(n_686),
    .B2(n_3466),
    .Y(n_1370));
 INVxp33_ASAP7_75t_R g43405 (.A(n_1366),
    .Y(u1_n_1044));
 INVxp33_ASAP7_75t_R g43406 (.A(n_1365),
    .Y(u1_n_1046));
 AOI22xp33_ASAP7_75t_R g43407 (.A1(u1_n_992),
    .A2(n_1293),
    .B1(n_1344),
    .B2(n_1283),
    .Y(n_1364));
 AOI332xp33_ASAP7_75t_R g43408 (.A1(n_1293),
    .A2(n_27),
    .A3(u1_n_997),
    .B1(n_1293),
    .B2(u1_n_852),
    .B3(n_1237),
    .C1(n_1338),
    .C2(n_94),
    .Y(n_1363));
 OAI221xp5_ASAP7_75t_R g43409 (.A1(n_1303),
    .A2(u1_n_1592),
    .B1(n_1322),
    .B2(n_1284),
    .C(n_1359),
    .Y(n_1369));
 OAI221xp5_ASAP7_75t_R g43410 (.A1(u1_n_4917),
    .A2(n_1299),
    .B1(u1_n_4919),
    .B2(n_1313),
    .C(n_1348),
    .Y(n_1368));
 OAI221xp5_ASAP7_75t_R g43411 (.A1(n_1330),
    .A2(n_1284),
    .B1(n_58),
    .B2(u1_n_1593),
    .C(n_1355),
    .Y(n_1367));
 AOI22xp33_ASAP7_75t_R g43412 (.A1(n_1344),
    .A2(n_1292),
    .B1(n_14154),
    .B2(n_687),
    .Y(n_1366));
 AOI22xp33_ASAP7_75t_R g43413 (.A1(u1_n_909),
    .A2(n_1281),
    .B1(n_14150),
    .B2(n_688),
    .Y(n_1365));
 AO22x1_ASAP7_75t_R g43414 (.A1(n_1279),
    .A2(u1_n_909),
    .B1(n_663),
    .B2(n_3454),
    .Y(u1_n_1019));
 AO22x1_ASAP7_75t_R g43415 (.A1(n_1295),
    .A2(n_1344),
    .B1(n_660),
    .B2(n_3456),
    .Y(u1_n_1017));
 AOI22xp33_ASAP7_75t_R g43416 (.A1(n_1294),
    .A2(n_1307),
    .B1(n_94),
    .B2(n_1327),
    .Y(n_1359));
 AOI22xp33_ASAP7_75t_R g43417 (.A1(n_1283),
    .A2(n_1297),
    .B1(n_94),
    .B2(n_1339),
    .Y(n_1358));
 NAND2xp33_ASAP7_75t_R g43418 (.A(n_1344),
    .B(n_94),
    .Y(n_1357));
 AOI22xp33_ASAP7_75t_R g43419 (.A1(n_1293),
    .A2(u1_n_980),
    .B1(n_94),
    .B2(n_1328),
    .Y(n_1356));
 AOI22xp33_ASAP7_75t_R g43420 (.A1(n_1293),
    .A2(u1_n_986),
    .B1(n_94),
    .B2(n_1329),
    .Y(n_1355));
 OAI222xp33_ASAP7_75t_R g43421 (.A1(n_1330),
    .A2(u1_n_1594),
    .B1(u1_n_1592),
    .B2(n_1298),
    .C1(u1_n_1593),
    .C2(n_1311),
    .Y(n_1362));
 NAND2xp33_ASAP7_75t_R g43422 (.A(u1_n_1041),
    .B(n_1341),
    .Y(n_1361));
 OAI222xp33_ASAP7_75t_R g43423 (.A1(u1_n_1592),
    .A2(n_1310),
    .B1(n_1332),
    .B2(u1_n_1594),
    .C1(u1_n_1593),
    .C2(n_1309),
    .Y(n_1360));
 OAI21xp33_ASAP7_75t_R g43424 (.A1(n_51),
    .A2(n_1296),
    .B(n_1343),
    .Y(u1_n_915));
 OAI222xp33_ASAP7_75t_R g43425 (.A1(n_1313),
    .A2(u1_n_5054),
    .B1(n_1299),
    .B2(n_1287),
    .C1(n_1318),
    .C2(u1_n_4993),
    .Y(u1_n_921));
 INVxp33_ASAP7_75t_R g43426 (.A(n_1354),
    .Y(u1_n_1042));
 INVxp33_ASAP7_75t_R g43427 (.A(n_1353),
    .Y(u1_n_1043));
 INVxp33_ASAP7_75t_R g43428 (.A(n_1352),
    .Y(u1_n_1045));
 INVxp33_ASAP7_75t_R g43429 (.A(n_1351),
    .Y(u1_n_1040));
 INVxp33_ASAP7_75t_R g43430 (.A(n_1350),
    .Y(u1_n_1016));
 INVxp33_ASAP7_75t_R g43431 (.A(n_1349),
    .Y(u1_n_1018));
 AOI22xp33_ASAP7_75t_R g43432 (.A1(u1_n_2218),
    .A2(n_1337),
    .B1(n_1286),
    .B2(u1_n_969),
    .Y(n_1348));
 AOI22xp33_ASAP7_75t_R g43433 (.A1(n_1338),
    .A2(n_1295),
    .B1(n_2896),
    .B2(n_1150),
    .Y(n_1347));
 AOI21xp33_ASAP7_75t_R g43434 (.A1(n_1286),
    .A2(u1_n_4761),
    .B(n_1321),
    .Y(n_1346));
 AO22x1_ASAP7_75t_R g43435 (.A1(n_1295),
    .A2(n_1333),
    .B1(n_686),
    .B2(n_3401),
    .Y(u1_n_1015));
 AOI22xp33_ASAP7_75t_R g43436 (.A1(n_1333),
    .A2(n_1292),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B2(n_688),
    .Y(n_1354));
 AOI22xp33_ASAP7_75t_R g43437 (.A1(n_1331),
    .A2(n_1292),
    .B1(n_14156),
    .B2(n_688),
    .Y(n_1353));
 AOI22xp33_ASAP7_75t_R g43438 (.A1(n_1336),
    .A2(n_1292),
    .B1(n_14152),
    .B2(n_688),
    .Y(n_1352));
 AO22x1_ASAP7_75t_R g43439 (.A1(n_1279),
    .A2(n_1337),
    .B1(n_686),
    .B2(n_3444),
    .Y(u1_n_1013));
 AOI22xp33_ASAP7_75t_R g43440 (.A1(n_1281),
    .A2(n_1337),
    .B1(n_687),
    .B2(u5_mul_69_18_n_143),
    .Y(n_1351));
 AOI22xp33_ASAP7_75t_R g43441 (.A1(n_1295),
    .A2(n_1331),
    .B1(n_663),
    .B2(n_3472),
    .Y(n_1350));
 AOI22xp33_ASAP7_75t_R g43442 (.A1(n_1295),
    .A2(n_1336),
    .B1(n_686),
    .B2(n_3452),
    .Y(n_1349));
 NAND2xp33_ASAP7_75t_R g43443 (.A(n_51),
    .B(n_1339),
    .Y(n_1343));
 NAND2xp33_ASAP7_75t_R g43444 (.A(n_1083),
    .B(u1_fractb_s[26]),
    .Y(n_1345));
 OAI22xp33_ASAP7_75t_R g43445 (.A1(n_695),
    .A2(n_1313),
    .B1(n_696),
    .B2(n_1318),
    .Y(n_1344));
 INVxp33_ASAP7_75t_R g43446 (.A(n_1341),
    .Y(u1_n_1014));
 OAI222xp33_ASAP7_75t_R g43447 (.A1(u1_n_1592),
    .A2(n_1302),
    .B1(n_1322),
    .B2(u1_n_1594),
    .C1(u1_n_1593),
    .C2(n_1312),
    .Y(n_1342));
 AOI22xp33_ASAP7_75t_R g43448 (.A1(n_1295),
    .A2(n_1323),
    .B1(n_686),
    .B2(n_3474),
    .Y(n_1341));
 OAI222xp33_ASAP7_75t_R g43449 (.A1(n_1314),
    .A2(u1_n_4993),
    .B1(n_1309),
    .B2(n_1287),
    .C1(n_1315),
    .C2(u1_n_5054),
    .Y(u1_n_909));
 AO22x1_ASAP7_75t_R g43450 (.A1(n_1292),
    .A2(n_1323),
    .B1(n_688),
    .B2(n_14160),
    .Y(u1_n_1041));
 INVxp33_ASAP7_75t_R g43451 (.A(n_1336),
    .Y(n_1335));
 OAI22xp33_ASAP7_75t_R g43452 (.A1(u1_n_840),
    .A2(n_1305),
    .B1(n_694),
    .B2(n_1310),
    .Y(u1_n_4761));
 NAND2xp33_ASAP7_75t_R g43453 (.A(u1_n_1039),
    .B(n_1320),
    .Y(n_1340));
 NAND2xp33_ASAP7_75t_R g43454 (.A(n_1275),
    .B(n_1324),
    .Y(u1_fractb_s[26]));
 OAI22xp33_ASAP7_75t_R g43455 (.A1(u1_n_840),
    .A2(n_1311),
    .B1(n_694),
    .B2(n_1317),
    .Y(n_1339));
 OAI22xp33_ASAP7_75t_R g43456 (.A1(n_695),
    .A2(n_1306),
    .B1(n_696),
    .B2(n_1302),
    .Y(n_1338));
 NOR2xp33_ASAP7_75t_R g43457 (.A(n_1287),
    .B(n_1318),
    .Y(n_1337));
 OAI22xp33_ASAP7_75t_R g43458 (.A1(n_695),
    .A2(n_1312),
    .B1(n_696),
    .B2(n_1316),
    .Y(n_1336));
 INVxp33_ASAP7_75t_R g43459 (.A(n_1326),
    .Y(n_1334));
 INVxp33_ASAP7_75t_R g43460 (.A(n_1333),
    .Y(n_1332));
 INVxp33_ASAP7_75t_R g43461 (.A(n_1331),
    .Y(n_1330));
 OAI22xp33_ASAP7_75t_R g43462 (.A1(n_695),
    .A2(n_1298),
    .B1(n_694),
    .B2(n_1311),
    .Y(n_1329));
 OAI22xp33_ASAP7_75t_R g43463 (.A1(n_695),
    .A2(n_1310),
    .B1(n_696),
    .B2(n_1309),
    .Y(n_1328));
 OAI22xp33_ASAP7_75t_R g43464 (.A1(n_695),
    .A2(n_1302),
    .B1(n_696),
    .B2(n_1312),
    .Y(n_1327));
 OAI22xp33_ASAP7_75t_R g43465 (.A1(n_1300),
    .A2(u1_n_840),
    .B1(n_1299),
    .B2(n_694),
    .Y(n_1326));
 OAI22xp33_ASAP7_75t_R g43466 (.A1(u1_n_840),
    .A2(n_1304),
    .B1(n_694),
    .B2(n_1300),
    .Y(u1_n_969));
 OAI22xp33_ASAP7_75t_R g43467 (.A1(n_695),
    .A2(n_1315),
    .B1(n_696),
    .B2(n_1314),
    .Y(n_1333));
 OAI32xp33_ASAP7_75t_R g43468 (.A1(n_1290),
    .A2(n_1248),
    .A3(n_696),
    .B1(u1_n_840),
    .B2(n_1317),
    .Y(n_1331));
 INVxp33_ASAP7_75t_R g43469 (.A(n_1324),
    .Y(n_1325));
 INVxp33_ASAP7_75t_R g43470 (.A(n_1323),
    .Y(n_1322));
 NOR2xp33_ASAP7_75t_R g43471 (.A(u1_n_4919),
    .B(n_1315),
    .Y(n_1321));
 NOR2xp33_ASAP7_75t_R g43472 (.A(n_1287),
    .B(n_1314),
    .Y(n_1324));
 NOR2xp33_ASAP7_75t_R g43473 (.A(u1_n_840),
    .B(n_1316),
    .Y(n_1323));
 INVxp33_ASAP7_75t_R g43474 (.A(n_1320),
    .Y(u1_n_1012));
 INVxp33_ASAP7_75t_R g43475 (.A(n_1319),
    .Y(u1_n_1039));
 AOI22xp33_ASAP7_75t_R g43476 (.A1(n_1295),
    .A2(n_1297),
    .B1(n_660),
    .B2(n_3386),
    .Y(n_1320));
 AOI22xp33_ASAP7_75t_R g43477 (.A1(n_1297),
    .A2(n_1292),
    .B1(n_14164),
    .B2(n_687),
    .Y(n_1319));
 AOI32xp33_ASAP7_75t_R g43478 (.A1(n_658),
    .A2(n_657),
    .A3(n_1116),
    .B1(n_1291),
    .B2(n_1236),
    .Y(n_1318));
 NOR2xp33_ASAP7_75t_R g43479 (.A(n_3496),
    .B(n_3850),
    .Y(n_3802));
 AO21x1_ASAP7_75t_R g43480 (.A1(exp_ovf_r[0]),
    .A2(n_3503),
    .B(exp_ovf_r[1]),
    .Y(n_1308));
 AOI22xp33_ASAP7_75t_R g43481 (.A1(n_1256),
    .A2(n_1291),
    .B1(n_1250),
    .B2(n_1290),
    .Y(n_1317));
 AOI22xp33_ASAP7_75t_R g43482 (.A1(n_1250),
    .A2(n_697),
    .B1(n_1247),
    .B2(n_658),
    .Y(n_1316));
 AOI22xp33_ASAP7_75t_R g43483 (.A1(n_1257),
    .A2(n_1291),
    .B1(n_1236),
    .B2(n_658),
    .Y(n_1315));
 NAND3xp33_ASAP7_75t_R g43484 (.A(n_1291),
    .B(n_657),
    .C(n_1116),
    .Y(n_1314));
 AOI22xp33_ASAP7_75t_R g43485 (.A1(n_1255),
    .A2(n_1291),
    .B1(n_1257),
    .B2(n_658),
    .Y(n_1313));
 AOI22xp33_ASAP7_75t_R g43486 (.A1(n_1254),
    .A2(n_1291),
    .B1(n_1256),
    .B2(n_658),
    .Y(n_1312));
 AOI22xp33_ASAP7_75t_R g43487 (.A1(n_1252),
    .A2(n_1291),
    .B1(n_1254),
    .B2(n_658),
    .Y(n_1311));
 AOI22xp33_ASAP7_75t_R g43488 (.A1(n_1241),
    .A2(n_1291),
    .B1(n_1251),
    .B2(n_658),
    .Y(n_1310));
 AOI22xp33_ASAP7_75t_R g43489 (.A1(n_1253),
    .A2(n_1291),
    .B1(n_1255),
    .B2(n_1290),
    .Y(n_1309));
 INVxp33_ASAP7_75t_R g43490 (.A(n_1306),
    .Y(n_1307));
 INVxp33_ASAP7_75t_R g43492 (.A(n_1298),
    .Y(u1_n_937));
 AO22x1_ASAP7_75t_R g43493 (.A1(n_1238),
    .A2(n_654),
    .B1(n_1240),
    .B2(n_658),
    .Y(u1_n_980));
 AOI22xp33_ASAP7_75t_R g43494 (.A1(n_1243),
    .A2(n_1291),
    .B1(n_1258),
    .B2(n_1290),
    .Y(n_1306));
 AOI22xp33_ASAP7_75t_R g43495 (.A1(n_1234),
    .A2(n_27),
    .B1(n_1259),
    .B2(u1_n_852),
    .Y(n_1305));
 AO22x1_ASAP7_75t_R g43496 (.A1(n_1237),
    .A2(n_654),
    .B1(n_1239),
    .B2(n_1290),
    .Y(u1_n_986));
 AOI22xp33_ASAP7_75t_R g43497 (.A1(n_1240),
    .A2(n_27),
    .B1(n_1234),
    .B2(u1_n_852),
    .Y(n_1304));
 AOI22xp33_ASAP7_75t_R g43498 (.A1(n_1239),
    .A2(n_1291),
    .B1(n_1242),
    .B2(n_1290),
    .Y(n_1303));
 AO22x1_ASAP7_75t_R g43499 (.A1(u1_n_3397),
    .A2(n_697),
    .B1(n_1238),
    .B2(u1_n_852),
    .Y(u1_n_992));
 AOI22xp33_ASAP7_75t_R g43500 (.A1(n_1260),
    .A2(n_697),
    .B1(n_1252),
    .B2(n_1290),
    .Y(n_1302));
 AOI22xp33_ASAP7_75t_R g43501 (.A1(n_1242),
    .A2(n_27),
    .B1(n_1243),
    .B2(u1_n_852),
    .Y(n_58));
 AOI22xp33_ASAP7_75t_R g43502 (.A1(n_1259),
    .A2(n_1291),
    .B1(n_1241),
    .B2(n_1290),
    .Y(n_1300));
 AOI22xp33_ASAP7_75t_R g43503 (.A1(n_1251),
    .A2(n_1291),
    .B1(n_1253),
    .B2(n_1290),
    .Y(n_1299));
 AOI22xp33_ASAP7_75t_R g43504 (.A1(n_1258),
    .A2(n_1291),
    .B1(n_1260),
    .B2(n_658),
    .Y(n_1298));
 OR2x2_ASAP7_75t_R g43505 (.A(exp_ovf_r[0]),
    .B(n_26),
    .Y(n_3496));
 INVxp33_ASAP7_75t_R g43506 (.A(n_1297),
    .Y(n_1296));
 NOR3xp33_ASAP7_75t_R g43508 (.A(u1_n_852),
    .B(n_1248),
    .C(u1_n_840),
    .Y(n_1297));
 INVxp33_ASAP7_75t_R g43509 (.A(u1_n_1593),
    .Y(n_1294));
 INVxp33_ASAP7_75t_R g43510 (.A(u1_n_1592),
    .Y(n_1293));
 NOR2xp33_ASAP7_75t_R g43512 (.A(n_1152),
    .B(n_1285),
    .Y(n_1295));
 NAND2xp33_ASAP7_75t_R g43513 (.A(n_695),
    .B(n_1286),
    .Y(u1_n_1593));
 NAND2xp33_ASAP7_75t_R g43514 (.A(n_696),
    .B(n_1286),
    .Y(u1_n_1592));
 INVxp33_ASAP7_75t_R g43516 (.A(u1_n_852),
    .Y(n_27));
 INVxp33_ASAP7_75t_R g43519 (.A(n_1291),
    .Y(u1_n_852));
 INVxp33_ASAP7_75t_R g43520 (.A(n_1290),
    .Y(n_1291));
 NAND2xp33_ASAP7_75t_R g43524 (.A(u1_n_840),
    .B(n_94),
    .Y(u1_n_4919));
 NAND2xp33_ASAP7_75t_R g43525 (.A(n_694),
    .B(n_94),
    .Y(u1_n_4917));
 NOR2xp33_ASAP7_75t_R g43526 (.A(n_1151),
    .B(n_1285),
    .Y(n_1292));
 OAI21xp33_ASAP7_75t_R g43527 (.A1(n_1204),
    .A2(n_1232),
    .B(n_1282),
    .Y(n_1290));
 INVxp33_ASAP7_75t_R g43528 (.A(exp_ovf[0]),
    .Y(n_1289));
 INVxp33_ASAP7_75t_R g43529 (.A(n_94),
    .Y(u1_n_1594));
 NAND2xp33_ASAP7_75t_R g43531 (.A(u1_n_840),
    .B(n_51),
    .Y(u1_n_5054));
 NAND2xp33_ASAP7_75t_R g43532 (.A(n_694),
    .B(u1_n_850),
    .Y(u1_n_4993));
 NOR2xp33_ASAP7_75t_R g43533 (.A(u1_n_2218),
    .B(n_51),
    .Y(n_94));
 INVxp33_ASAP7_75t_R g43534 (.A(n_1286),
    .Y(n_1285));
 INVxp33_ASAP7_75t_R g43535 (.A(n_1284),
    .Y(n_1283));
 AOI22xp33_ASAP7_75t_R g43536 (.A1(n_1276),
    .A2(u1_n_2218),
    .B1(n_1204),
    .B2(n_1232),
    .Y(n_1282));
 OAI21xp33_ASAP7_75t_R g43537 (.A1(exp_ovf_r[1]),
    .A2(n_3502),
    .B(n_1020),
    .Y(n_3529));
 NAND2xp33_ASAP7_75t_R g43538 (.A(n_694),
    .B(n_51),
    .Y(n_1287));
 NOR2xp33_ASAP7_75t_R g43539 (.A(u1_n_2218),
    .B(u1_n_850),
    .Y(n_1286));
 NAND2xp33_ASAP7_75t_R g43540 (.A(u1_n_2218),
    .B(n_51),
    .Y(n_1284));
 INVxp33_ASAP7_75t_R g43541 (.A(n_51),
    .Y(u1_n_850));
 NOR2xp33_ASAP7_75t_R g43542 (.A(n_689),
    .B(u1_n_2218),
    .Y(n_1281));
 NOR2xp33_ASAP7_75t_R g43543 (.A(n_1267),
    .B(n_1276),
    .Y(n_51));
 NOR2xp33_ASAP7_75t_R g43545 (.A(n_1150),
    .B(u1_n_2218),
    .Y(n_1279));
 INVxp33_ASAP7_75t_R g43546 (.A(exp_ovf_r[1]),
    .Y(n_26));
 INVxp33_ASAP7_75t_R g43548 (.A(u1_n_2218),
    .Y(n_1275));
 OAI211xp5_ASAP7_75t_R g43549 (.A1(n_696),
    .A2(n_1266),
    .B(n_1273),
    .C(n_1235),
    .Y(n_1276));
 NAND3xp33_ASAP7_75t_R g43550 (.A(n_1273),
    .B(n_1269),
    .C(n_1235),
    .Y(u1_n_2218));
 INVxp33_ASAP7_75t_R g43551 (.A(exp_ovf[1]),
    .Y(n_1274));
 NAND2xp33_ASAP7_75t_R g43553 (.A(u2_n_606),
    .B(u2_exp_ovf_d[1]),
    .Y(u2_n_772));
 OAI211xp5_ASAP7_75t_R g43554 (.A1(n_1170),
    .A2(n_1162),
    .B(n_1270),
    .C(n_1224),
    .Y(n_1273));
 INVxp33_ASAP7_75t_R g43555 (.A(u2_exp_ovf_d[1]),
    .Y(n_1272));
 XNOR2xp5_ASAP7_75t_R g43556 (.A(n_1271),
    .B(u2_n_710),
    .Y(u2_exp_ovf_d[1]));
 AO32x1_ASAP7_75t_R g43557 (.A1(u2_n_140),
    .A2(u2_exp_tmp1[6]),
    .A3(u2_n_606),
    .B1(n_1265),
    .B2(u2_exp_tmp1[7]),
    .Y(n_1271));
 AOI22xp33_ASAP7_75t_R g43558 (.A1(n_1268),
    .A2(n_1225),
    .B1(n_1170),
    .B2(n_1162),
    .Y(n_1270));
 XNOR2xp5_ASAP7_75t_R g43559 (.A(n_1268),
    .B(n_1229),
    .Y(n_1269));
 AOI21xp33_ASAP7_75t_R g43560 (.A1(n_1263),
    .A2(n_1209),
    .B(n_1206),
    .Y(n_1268));
 INVxp33_ASAP7_75t_R g43561 (.A(n_1266),
    .Y(n_1267));
 OR3x1_ASAP7_75t_R g43562 (.A(u2_n_140),
    .B(u2_exp_tmp1[6]),
    .C(n_13981),
    .Y(n_1265));
 XNOR2xp5_ASAP7_75t_R g43563 (.A(n_1263),
    .B(n_1216),
    .Y(n_1266));
 XNOR2xp5_ASAP7_75t_R g43564 (.A(n_1261),
    .B(n_1077),
    .Y(n_1264));
 OAI21xp33_ASAP7_75t_R g43565 (.A1(n_13981),
    .A2(n_1228),
    .B(u2_n_1831),
    .Y(u2_n_140));
 OAI21xp33_ASAP7_75t_R g43566 (.A1(n_1210),
    .A2(n_1249),
    .B(n_1201),
    .Y(n_1263));
 INVxp33_ASAP7_75t_R g43570 (.A(n_695),
    .Y(n_696));
 INVxp33_ASAP7_75t_R g43580 (.A(u1_n_840),
    .Y(n_694));
 HB1xp67_ASAP7_75t_R g43583 (.A(n_695),
    .Y(u1_n_840));
 XOR2xp5_ASAP7_75t_R g43586 (.A(n_1233),
    .B(n_1053),
    .Y(u2_exp_tmp1[7]));
 XNOR2xp5_ASAP7_75t_R g43587 (.A(n_1217),
    .B(n_1249),
    .Y(n_695));
 NAND2xp33_ASAP7_75t_R g43588 (.A(opa_r1[22]),
    .B(n_1246),
    .Y(n_1262));
 NAND2xp33_ASAP7_75t_R g43589 (.A(u2_n_1384),
    .B(u2_n_1399),
    .Y(u2_n_1831));
 NOR2xp33_ASAP7_75t_R g43590 (.A(opa_r1[22]),
    .B(n_1245),
    .Y(n_1261));
 INVxp33_ASAP7_75t_R g43591 (.A(n_1247),
    .Y(n_1248));
 INVxp33_ASAP7_75t_R g43592 (.A(n_1245),
    .Y(n_1246));
 NAND2xp33_ASAP7_75t_R g43593 (.A(opa_r1[21]),
    .B(n_1231),
    .Y(n_1244));
 OAI22xp33_ASAP7_75t_R g43594 (.A1(n_1218),
    .A2(n_1181),
    .B1(n_693),
    .B2(n_1185),
    .Y(n_1260));
 NAND2xp33_ASAP7_75t_R g43595 (.A(u2_n_1487),
    .B(u2_n_606),
    .Y(u2_n_1399));
 OAI22xp33_ASAP7_75t_R g43596 (.A1(n_1182),
    .A2(u1_n_853),
    .B1(n_1183),
    .B2(n_657),
    .Y(n_1259));
 OAI22xp33_ASAP7_75t_R g43597 (.A1(n_1218),
    .A2(n_1183),
    .B1(n_693),
    .B2(n_1184),
    .Y(n_1258));
 OAI22xp33_ASAP7_75t_R g43598 (.A1(n_1190),
    .A2(n_1218),
    .B1(n_1191),
    .B2(n_693),
    .Y(n_1257));
 OAI22xp33_ASAP7_75t_R g43599 (.A1(n_1189),
    .A2(n_1218),
    .B1(n_1190),
    .B2(n_693),
    .Y(n_1256));
 OAI22xp33_ASAP7_75t_R g43600 (.A1(n_1218),
    .A2(n_1188),
    .B1(n_693),
    .B2(n_1189),
    .Y(n_1255));
 OAI22xp33_ASAP7_75t_R g43601 (.A1(n_1218),
    .A2(n_1187),
    .B1(n_693),
    .B2(n_1188),
    .Y(n_1254));
 OAI22xp33_ASAP7_75t_R g43602 (.A1(n_1218),
    .A2(n_1186),
    .B1(n_693),
    .B2(n_1187),
    .Y(n_1253));
 OAI22xp33_ASAP7_75t_R g43603 (.A1(n_1218),
    .A2(n_1177),
    .B1(n_693),
    .B2(n_1186),
    .Y(n_1252));
 OAI22xp33_ASAP7_75t_R g43604 (.A1(n_1218),
    .A2(n_1185),
    .B1(n_693),
    .B2(n_1177),
    .Y(n_1251));
 OAI22xp33_ASAP7_75t_R g43605 (.A1(n_1218),
    .A2(n_1191),
    .B1(n_693),
    .B2(n_1192),
    .Y(n_1250));
 AOI21xp33_ASAP7_75t_R g43606 (.A1(n_1220),
    .A2(n_1203),
    .B(n_1226),
    .Y(n_1249));
 OAI21xp33_ASAP7_75t_R g43607 (.A1(n_1218),
    .A2(n_1163),
    .B(n_1144),
    .Y(n_1247));
 NAND2xp33_ASAP7_75t_R g43608 (.A(n_724),
    .B(n_1231),
    .Y(n_1245));
 OAI22xp33_ASAP7_75t_R g43609 (.A1(n_1218),
    .A2(n_1180),
    .B1(n_693),
    .B2(n_1182),
    .Y(n_1243));
 OAI22xp33_ASAP7_75t_R g43610 (.A1(n_1178),
    .A2(u1_n_853),
    .B1(n_1179),
    .B2(n_657),
    .Y(n_1242));
 OAI22xp33_ASAP7_75t_R g43611 (.A1(n_1218),
    .A2(n_1184),
    .B1(n_693),
    .B2(n_1181),
    .Y(n_1241));
 OAI22xp33_ASAP7_75t_R g43612 (.A1(u1_n_853),
    .A2(n_1169),
    .B1(n_657),
    .B2(n_1178),
    .Y(n_1240));
 OAI22xp33_ASAP7_75t_R g43613 (.A1(n_1172),
    .A2(u1_n_853),
    .B1(n_1169),
    .B2(n_657),
    .Y(n_1239));
 OAI22xp33_ASAP7_75t_R g43614 (.A1(u1_n_853),
    .A2(n_1171),
    .B1(n_657),
    .B2(n_1172),
    .Y(n_1238));
 OAI22xp33_ASAP7_75t_R g43615 (.A1(u1_n_853),
    .A2(n_1167),
    .B1(n_657),
    .B2(n_1171),
    .Y(n_1237));
 OAI22xp33_ASAP7_75t_R g43616 (.A1(u1_n_853),
    .A2(n_1166),
    .B1(n_657),
    .B2(n_1167),
    .Y(u1_n_3397));
 OAI22xp33_ASAP7_75t_R g43617 (.A1(n_1176),
    .A2(u1_n_853),
    .B1(n_1166),
    .B2(n_657),
    .Y(u1_n_997));
 OAI22xp33_ASAP7_75t_R g43618 (.A1(n_1218),
    .A2(n_1192),
    .B1(n_693),
    .B2(n_1163),
    .Y(n_1236));
 OAI31xp33_ASAP7_75t_R g43620 (.A1(n_1205),
    .A2(n_1173),
    .A3(u1_exp_large[6]),
    .B(n_1227),
    .Y(n_1235));
 XOR2xp5_ASAP7_75t_R g43621 (.A(n_1219),
    .B(opa_r[30]),
    .Y(n_1233));
 OAI22xp33_ASAP7_75t_R g43622 (.A1(u1_n_853),
    .A2(n_1179),
    .B1(n_657),
    .B2(n_1180),
    .Y(n_1234));
 XOR2xp5_ASAP7_75t_R g43623 (.A(n_1215),
    .B(opa_r[29]),
    .Y(u2_exp_tmp1[6]));
 MAJIxp5_ASAP7_75t_R g43624 (.A(n_1219),
    .B(n_62),
    .C(n_1053),
    .Y(u2_n_710));
 NAND2xp33_ASAP7_75t_R g43625 (.A(opa_r1[20]),
    .B(n_1223),
    .Y(n_1230));
 AOI21xp33_ASAP7_75t_R g43626 (.A1(n_1207),
    .A2(n_1164),
    .B(n_1226),
    .Y(n_1232));
 NAND2xp33_ASAP7_75t_R g43627 (.A(n_1224),
    .B(n_1225),
    .Y(n_1229));
 NOR2xp33_ASAP7_75t_R g43628 (.A(opa_r1[20]),
    .B(n_1222),
    .Y(n_1231));
 NOR2xp33_ASAP7_75t_R g43629 (.A(u2_exp_tmp1[4]),
    .B(u2_exp_tmp1[5]),
    .Y(n_1228));
 NAND2xp33_ASAP7_75t_R g43630 (.A(n_683),
    .B(u2_exp_tmp1[5]),
    .Y(u2_n_1792));
 AO32x1_ASAP7_75t_R g43631 (.A1(n_1205),
    .A2(u1_exp_large[6]),
    .A3(n_1173),
    .B1(n_1001),
    .B2(u1_exp_large[7]),
    .Y(n_1227));
 NAND5xp2_ASAP7_75t_R g43632 (.A(n_3581),
    .B(n_3583),
    .C(n_700),
    .D(n_24),
    .E(n_792),
    .Y(n_3592));
 NAND2xp33_ASAP7_75t_R g43633 (.A(u2_exp_tmp1[4]),
    .B(u2_exp_tmp1[5]),
    .Y(u2_n_1487));
 INVxp33_ASAP7_75t_R g43634 (.A(n_1222),
    .Y(n_1223));
 NAND2xp33_ASAP7_75t_R g43635 (.A(opa_r1[19]),
    .B(n_1214),
    .Y(n_1221));
 NAND2xp33_ASAP7_75t_R g43636 (.A(n_1164),
    .B(n_1207),
    .Y(n_1220));
 NOR2xp33_ASAP7_75t_R g43637 (.A(n_1164),
    .B(n_1207),
    .Y(n_1226));
 NAND2xp33_ASAP7_75t_R g43638 (.A(u1_exp_large[4]),
    .B(n_1212),
    .Y(n_1225));
 NAND2xp33_ASAP7_75t_R g43639 (.A(n_1168),
    .B(n_1211),
    .Y(n_1224));
 NAND2xp33_ASAP7_75t_R g43640 (.A(n_721),
    .B(n_1214),
    .Y(n_1222));
 OAI211xp5_ASAP7_75t_R g43665 (.A1(u2_n_1448),
    .A2(n_1194),
    .B(u2_n_1777),
    .C(u2_n_1475),
    .Y(u2_n_1384));
 AOI21xp33_ASAP7_75t_R g43666 (.A1(u1_exp_large[2]),
    .A2(n_1175),
    .B(n_1210),
    .Y(n_1217));
 NOR2xp33_ASAP7_75t_R g43667 (.A(n_1208),
    .B(n_1206),
    .Y(n_1216));
 XOR2xp5_ASAP7_75t_R g43668 (.A(n_1197),
    .B(n_1047),
    .Y(n_1215));
 MAJIxp5_ASAP7_75t_R g43669 (.A(n_1198),
    .B(opa_r[29]),
    .C(n_1048),
    .Y(n_1219));
 XOR2xp5_ASAP7_75t_R g43670 (.A(n_1195),
    .B(opa_r[28]),
    .Y(u2_exp_tmp1[5]));
 OAI21xp33_ASAP7_75t_R g43671 (.A1(n_1116),
    .A2(n_1202),
    .B(n_1144),
    .Y(n_1218));
 NAND2xp33_ASAP7_75t_R g43672 (.A(opa_r1[18]),
    .B(n_1200),
    .Y(n_1213));
 NAND2xp33_ASAP7_75t_R g43673 (.A(u2_exp_tmp1[4]),
    .B(n_683),
    .Y(u2_n_1444));
 NOR2xp33_ASAP7_75t_R g43674 (.A(opa_r1[18]),
    .B(n_1199),
    .Y(n_1214));
 INVxp33_ASAP7_75t_R g43675 (.A(n_1211),
    .Y(n_1212));
 INVxp33_ASAP7_75t_R g43676 (.A(n_1208),
    .Y(n_1209));
 AOI21xp33_ASAP7_75t_R g43677 (.A1(n_1159),
    .A2(n_1116),
    .B(n_1125),
    .Y(n_1211));
 AOI21xp33_ASAP7_75t_R g43678 (.A1(n_1175),
    .A2(u1_fracta_s[26]),
    .B(u1_exp_large[2]),
    .Y(n_1210));
 AOI21xp33_ASAP7_75t_R g43679 (.A1(n_1174),
    .A2(u1_fracta_s[26]),
    .B(u1_exp_large[3]),
    .Y(n_1208));
 AOI21xp33_ASAP7_75t_R g43680 (.A1(n_1161),
    .A2(n_1116),
    .B(n_1125),
    .Y(n_1207));
 INVxp33_ASAP7_75t_R g43681 (.A(n_1204),
    .Y(n_1203));
 NAND2xp33_ASAP7_75t_R g43682 (.A(n_1137),
    .B(n_1165),
    .Y(n_1202));
 AND2x2_ASAP7_75t_R g43683 (.A(u1_exp_large[3]),
    .B(n_1174),
    .Y(n_1206));
 OR2x2_ASAP7_75t_R g43684 (.A(n_1170),
    .B(u1_exp_large[5]),
    .Y(n_1205));
 NAND2xp33_ASAP7_75t_R g43685 (.A(u1_exp_large[2]),
    .B(n_1175),
    .Y(n_1201));
 NOR2xp33_ASAP7_75t_R g43686 (.A(n_1128),
    .B(u1_exp_large[0]),
    .Y(n_1204));
 INVxp33_ASAP7_75t_R g43687 (.A(n_1199),
    .Y(n_1200));
 INVxp33_ASAP7_75t_R g43688 (.A(n_1197),
    .Y(n_1198));
 NAND2xp33_ASAP7_75t_R g43689 (.A(opa_r1[17]),
    .B(n_1193),
    .Y(n_1196));
 XOR2xp5_ASAP7_75t_R g43691 (.A(n_1156),
    .B(n_1044),
    .Y(n_1195));
 NAND2xp33_ASAP7_75t_R g43692 (.A(n_799),
    .B(n_1193),
    .Y(n_1199));
 MAJIxp5_ASAP7_75t_R g43693 (.A(n_1157),
    .B(opa_r[28]),
    .C(n_1045),
    .Y(n_1197));
 XOR2xp5_ASAP7_75t_R g43694 (.A(n_646),
    .B(opa_r[27]),
    .Y(u2_exp_tmp1[4]));
 INVxp33_ASAP7_75t_R g43695 (.A(n_1194),
    .Y(u2_n_1489));
 INVxp33_ASAP7_75t_R g43696 (.A(n_1192),
    .Y(u1_n_867));
 INVxp33_ASAP7_75t_R g43697 (.A(n_1191),
    .Y(u1_n_873));
 INVxp33_ASAP7_75t_R g43698 (.A(n_1190),
    .Y(u1_n_880));
 INVxp33_ASAP7_75t_R g43699 (.A(n_1189),
    .Y(u1_n_886));
 INVxp33_ASAP7_75t_R g43703 (.A(n_1185),
    .Y(u1_n_917));
 INVxp33_ASAP7_75t_R g43706 (.A(n_1182),
    .Y(u1_n_941));
 INVxp33_ASAP7_75t_R g43707 (.A(n_1181),
    .Y(u1_n_923));
 INVxp33_ASAP7_75t_R g43708 (.A(n_1180),
    .Y(u1_n_947));
 NAND2xp33_ASAP7_75t_R g43712 (.A(n_3718),
    .B(n_3507),
    .Y(n_3581));
 NAND2xp33_ASAP7_75t_R g43713 (.A(n_656),
    .B(n_14295),
    .Y(u2_n_1777));
 NOR2xp33_ASAP7_75t_R g43714 (.A(n_656),
    .B(n_14295),
    .Y(n_1194));
 NOR2xp33_ASAP7_75t_R g43715 (.A(opa_r1[16]),
    .B(n_1158),
    .Y(n_1193));
 AOI22xp33_ASAP7_75t_R g43716 (.A1(n_691),
    .A2(u5_mul_69_18_n_143),
    .B1(n_670),
    .B2(n_3444),
    .Y(n_1192));
 AOI22xp33_ASAP7_75t_R g43717 (.A1(n_691),
    .A2(n_14160),
    .B1(n_690),
    .B2(n_3474),
    .Y(n_1191));
 AOI22xp33_ASAP7_75t_R g43718 (.A1(n_691),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B1(n_670),
    .B2(n_3401),
    .Y(n_1190));
 AOI22xp33_ASAP7_75t_R g43719 (.A1(n_691),
    .A2(n_14156),
    .B1(n_670),
    .B2(n_3472),
    .Y(n_1189));
 AOI22xp33_ASAP7_75t_R g43720 (.A1(n_691),
    .A2(n_14154),
    .B1(n_670),
    .B2(n_3456),
    .Y(n_1188));
 AOI22xp33_ASAP7_75t_R g43721 (.A1(n_691),
    .A2(n_14152),
    .B1(n_670),
    .B2(n_3452),
    .Y(n_1187));
 AOI22xp33_ASAP7_75t_R g43722 (.A1(n_691),
    .A2(n_14150),
    .B1(n_690),
    .B2(n_3454),
    .Y(n_1186));
 AOI22xp33_ASAP7_75t_R g43723 (.A1(n_691),
    .A2(n_14146),
    .B1(n_690),
    .B2(n_3476),
    .Y(n_1185));
 AOI22xp33_ASAP7_75t_R g43724 (.A1(n_691),
    .A2(n_14142),
    .B1(n_690),
    .B2(n_3468),
    .Y(n_1184));
 AOI22xp33_ASAP7_75t_R g43725 (.A1(n_691),
    .A2(n_14140),
    .B1(n_690),
    .B2(n_3432),
    .Y(n_1183));
 AOI22xp33_ASAP7_75t_R g43726 (.A1(n_691),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B1(n_670),
    .B2(n_3438),
    .Y(n_1182));
 AOI22xp33_ASAP7_75t_R g43727 (.A1(n_691),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .B1(n_670),
    .B2(n_3466),
    .Y(n_1181));
 AOI22xp33_ASAP7_75t_R g43728 (.A1(n_691),
    .A2(n_14136),
    .B1(n_690),
    .B2(n_2896),
    .Y(n_1180));
 AOI22xp33_ASAP7_75t_R g43729 (.A1(n_1152),
    .A2(n_14134),
    .B1(n_1151),
    .B2(n_3434),
    .Y(n_1179));
 AOI22xp33_ASAP7_75t_R g43730 (.A1(n_1152),
    .A2(n_14132),
    .B1(n_1151),
    .B2(n_3409),
    .Y(n_1178));
 AOI22xp33_ASAP7_75t_R g43731 (.A1(n_691),
    .A2(n_14148),
    .B1(n_690),
    .B2(n_3415),
    .Y(n_1177));
 INVxp33_ASAP7_75t_R g43732 (.A(n_1176),
    .Y(u1_n_996));
 INVxp33_ASAP7_75t_R g43733 (.A(n_1172),
    .Y(u1_n_972));
 INVxp33_ASAP7_75t_R g43734 (.A(n_1171),
    .Y(u1_n_978));
 INVxp33_ASAP7_75t_R g43735 (.A(n_1169),
    .Y(u1_n_966));
 INVxp33_ASAP7_75t_R g43736 (.A(n_1168),
    .Y(u1_exp_large[4]));
 INVxp33_ASAP7_75t_R g43737 (.A(n_1167),
    .Y(u1_n_984));
 INVxp33_ASAP7_75t_R g43738 (.A(n_1166),
    .Y(u1_n_990));
 INVxp33_ASAP7_75t_R g43739 (.A(n_1165),
    .Y(u1_exp_large[0]));
 INVxp33_ASAP7_75t_R g43740 (.A(n_1164),
    .Y(u1_exp_large[1]));
 INVxp33_ASAP7_75t_R g43742 (.A(n_1162),
    .Y(u1_exp_large[5]));
 OAI22xp33_ASAP7_75t_R g43743 (.A1(opb_r[24]),
    .A2(n_692),
    .B1(opa_r[24]),
    .B2(n_1153),
    .Y(n_1161));
 XNOR2xp5_ASAP7_75t_R g43744 (.A(n_1155),
    .B(opa_r1[15]),
    .Y(n_1160));
 OAI22xp33_ASAP7_75t_R g43745 (.A1(n_690),
    .A2(opb_r[27]),
    .B1(n_1153),
    .B2(opa_r[27]),
    .Y(n_1159));
 AOI22xp33_ASAP7_75t_R g43746 (.A1(n_1152),
    .A2(n_3303),
    .B1(n_1151),
    .B2(u5_mul_69_18_n_118),
    .Y(n_1176));
 AOI22xp33_ASAP7_75t_R g43747 (.A1(opb_r[25]),
    .A2(n_1153),
    .B1(opa_r[25]),
    .B2(n_690),
    .Y(n_1175));
 AOI22xp33_ASAP7_75t_R g43748 (.A1(n_1153),
    .A2(opb_r[26]),
    .B1(n_690),
    .B2(opa_r[26]),
    .Y(n_1174));
 AOI22xp33_ASAP7_75t_R g43749 (.A1(n_1153),
    .A2(opb_r[29]),
    .B1(n_692),
    .B2(opa_r[29]),
    .Y(n_1173));
 AOI22xp33_ASAP7_75t_R g43750 (.A1(n_1152),
    .A2(n_14128),
    .B1(n_1151),
    .B2(n_3440),
    .Y(n_1172));
 OAI22xp33_ASAP7_75t_R g43751 (.A1(n_42),
    .A2(n_690),
    .B1(n_714),
    .B2(n_1153),
    .Y(u1_exp_large[6]));
 AOI22xp33_ASAP7_75t_R g43752 (.A1(n_1152),
    .A2(n_14126),
    .B1(n_1151),
    .B2(n_3411),
    .Y(n_1171));
 AOI22xp33_ASAP7_75t_R g43753 (.A1(n_1153),
    .A2(opb_r[28]),
    .B1(n_690),
    .B2(opa_r[28]),
    .Y(n_1170));
 AOI22xp33_ASAP7_75t_R g43754 (.A1(n_1152),
    .A2(n_14130),
    .B1(n_1151),
    .B2(n_3395),
    .Y(n_1169));
 AOI22xp33_ASAP7_75t_R g43755 (.A1(opa_r[27]),
    .A2(n_1153),
    .B1(opb_r[27]),
    .B2(n_692),
    .Y(n_1168));
 AOI22xp33_ASAP7_75t_R g43756 (.A1(n_1152),
    .A2(n_14178),
    .B1(n_1151),
    .B2(n_3427),
    .Y(n_1167));
 OAI22xp33_ASAP7_75t_R g43757 (.A1(n_41),
    .A2(n_692),
    .B1(n_795),
    .B2(n_1153),
    .Y(u1_exp_large[3]));
 AOI22xp33_ASAP7_75t_R g43758 (.A1(n_1152),
    .A2(n_14124),
    .B1(n_1151),
    .B2(n_3436),
    .Y(n_1166));
 OAI22xp33_ASAP7_75t_R g43759 (.A1(n_44),
    .A2(n_692),
    .B1(n_713),
    .B2(n_1153),
    .Y(u1_exp_large[2]));
 AOI22xp33_ASAP7_75t_R g43760 (.A1(opa_r[23]),
    .A2(n_1153),
    .B1(opb_r[23]),
    .B2(n_692),
    .Y(n_1165));
 AOI22xp33_ASAP7_75t_R g43761 (.A1(opa_r[24]),
    .A2(n_1153),
    .B1(opb_r[24]),
    .B2(n_692),
    .Y(n_1164));
 AOI22xp33_ASAP7_75t_R g43762 (.A1(n_691),
    .A2(n_14164),
    .B1(n_670),
    .B2(n_3386),
    .Y(n_1163));
 AOI22xp33_ASAP7_75t_R g43763 (.A1(opa_r[28]),
    .A2(n_1153),
    .B1(opb_r[28]),
    .B2(n_692),
    .Y(n_1162));
 NAND2xp33_ASAP7_75t_R g43765 (.A(u2_n_1392),
    .B(u2_n_1494),
    .Y(u2_n_1448));
 NAND2xp33_ASAP7_75t_R g43766 (.A(n_3580),
    .B(n_1154),
    .Y(n_3718));
 NAND2xp33_ASAP7_75t_R g43767 (.A(n_719),
    .B(n_1155),
    .Y(n_1158));
 INVxp33_ASAP7_75t_R g43768 (.A(n_1156),
    .Y(n_1157));
 MAJIxp5_ASAP7_75t_R g43772 (.A(n_1147),
    .B(opa_r[27]),
    .C(n_1049),
    .Y(n_1156));
 NAND2xp33_ASAP7_75t_R g43773 (.A(n_3569),
    .B(n_3506),
    .Y(n_1154));
 OR2x2_ASAP7_75t_R g43774 (.A(n_656),
    .B(u2_exp_tmp1[2]),
    .Y(u2_n_1494));
 NOR2xp33_ASAP7_75t_R g43775 (.A(opa_r1[14]),
    .B(n_1148),
    .Y(n_1155));
 INVxp33_ASAP7_75t_R g43788 (.A(n_1151),
    .Y(n_1152));
 INVxp33_ASAP7_75t_R g43836 (.A(n_1151),
    .Y(n_1150));
 HB1xp67_ASAP7_75t_R g43837 (.A(n_670),
    .Y(n_1151));
 INVxp33_ASAP7_75t_R g43854 (.A(n_1153),
    .Y(n_692));
 XNOR2xp5_ASAP7_75t_R g43856 (.A(n_1145),
    .B(opa_r1[13]),
    .Y(n_1149));
 NAND2xp33_ASAP7_75t_R g43857 (.A(n_656),
    .B(u2_exp_tmp1[2]),
    .Y(u2_n_1475));
 AOI21xp33_ASAP7_75t_R g43858 (.A1(n_62),
    .A2(opb_r[30]),
    .B(n_1146),
    .Y(n_1153));
 AO21x1_ASAP7_75t_R g43862 (.A1(n_3563),
    .A2(n_3719),
    .B(n_1139),
    .Y(n_3569));
 NAND2xp33_ASAP7_75t_R g43863 (.A(n_723),
    .B(n_1145),
    .Y(n_1148));
 OAI332xp33_ASAP7_75t_R g43865 (.A1(n_1123),
    .A2(n_1000),
    .A3(n_879),
    .B1(n_878),
    .B2(opa_r[29]),
    .B3(n_714),
    .C1(n_1000),
    .C2(n_1032),
    .Y(n_1146));
 MAJx2_ASAP7_75t_R g43866 (.A(u2_exp_tmp1[1]),
    .B(n_656),
    .C(u2_exp_tmp1[0]),
    .Y(u2_n_1392));
 OAI32xp33_ASAP7_75t_R g43867 (.A1(n_1133),
    .A2(n_1134),
    .A3(n_44),
    .B1(opa_r[25]),
    .B2(n_1140),
    .Y(u2_exp_tmp1[2]));
 MAJIxp5_ASAP7_75t_R g43868 (.A(n_1141),
    .B(n_41),
    .C(n_1052),
    .Y(n_1147));
 NAND2xp33_ASAP7_75t_R g43869 (.A(n_683),
    .B(u2_exp_tmp1[1]),
    .Y(u2_n_1756));
 NOR2xp33_ASAP7_75t_R g43870 (.A(opa_r1[12]),
    .B(n_1142),
    .Y(n_1145));
 OR2x2_ASAP7_75t_R g43871 (.A(n_683),
    .B(u2_exp_tmp1[1]),
    .Y(u2_n_1398));
 XNOR2xp5_ASAP7_75t_R g43872 (.A(n_1138),
    .B(opa_r1[11]),
    .Y(n_1143));
 NAND3xp33_ASAP7_75t_R g43873 (.A(n_1136),
    .B(n_1116),
    .C(u1_n_8071),
    .Y(n_1144));
 AO21x1_ASAP7_75t_R g43875 (.A1(n_3575),
    .A2(n_3720),
    .B(n_1131),
    .Y(n_3719));
 NAND2xp33_ASAP7_75t_R g43876 (.A(n_720),
    .B(n_1138),
    .Y(n_1142));
 XOR2xp5_ASAP7_75t_R g43877 (.A(n_1122),
    .B(n_1046),
    .Y(u2_exp_tmp1[1]));
 XNOR2xp5_ASAP7_75t_R g43879 (.A(n_1126),
    .B(n_1050),
    .Y(n_1140));
 MAJIxp5_ASAP7_75t_R g43880 (.A(n_1127),
    .B(opa_r[25]),
    .C(n_1051),
    .Y(n_1141));
 INVxp33_ASAP7_75t_R g43881 (.A(n_3582),
    .Y(n_1139));
 NAND2xp33_ASAP7_75t_R g43882 (.A(div_opa_ldz_r2[2]),
    .B(n_706),
    .Y(n_3563));
 NAND2xp33_ASAP7_75t_R g43883 (.A(exp_r[2]),
    .B(n_1130),
    .Y(n_3582));
 NAND2xp33_ASAP7_75t_R g43884 (.A(n_1129),
    .B(exp_r[3]),
    .Y(n_3580));
 NAND2xp33_ASAP7_75t_R g43885 (.A(div_opa_ldz_r2[3]),
    .B(n_43),
    .Y(n_3506));
 NOR2xp33_ASAP7_75t_R g43886 (.A(opa_r1[10]),
    .B(n_1132),
    .Y(n_1138));
 INVxp33_ASAP7_75t_R g43887 (.A(n_1136),
    .Y(n_1137));
 XNOR2xp5_ASAP7_75t_R g43888 (.A(n_1118),
    .B(opa_r1[9]),
    .Y(n_1135));
 NOR2xp33_ASAP7_75t_R g43889 (.A(n_1051),
    .B(n_1126),
    .Y(n_1134));
 NOR2xp33_ASAP7_75t_R g43890 (.A(n_1050),
    .B(n_1127),
    .Y(n_1133));
 NOR2xp33_ASAP7_75t_R g43891 (.A(n_1128),
    .B(n_1125),
    .Y(n_1136));
 OR5x1_ASAP7_75t_R g43892 (.A(n_1124),
    .B(u4_n_1798),
    .C(u4_n_1805),
    .D(u4_n_1796),
    .E(u4_n_1803),
    .Y(n_3530));
 NAND2xp33_ASAP7_75t_R g43893 (.A(n_3720),
    .B(n_3576),
    .Y(n_3717));
 INVxp33_ASAP7_75t_R g43895 (.A(n_1131),
    .Y(n_3584));
 INVxp33_ASAP7_75t_R g43896 (.A(div_opa_ldz_r2[2]),
    .Y(n_1130));
 INVxp33_ASAP7_75t_R g43897 (.A(div_opa_ldz_r2[3]),
    .Y(n_1129));
 NAND2xp33_ASAP7_75t_R g43898 (.A(exp_r[0]),
    .B(n_1117),
    .Y(n_3576));
 NAND2xp33_ASAP7_75t_R g43900 (.A(n_722),
    .B(n_1118),
    .Y(n_1132));
 NAND2xp33_ASAP7_75t_R g43901 (.A(div_opa_ldz_r2[1]),
    .B(n_716),
    .Y(n_3575));
 NOR2xp33_ASAP7_75t_R g43902 (.A(div_opa_ldz_r2[1]),
    .B(n_716),
    .Y(n_1131));
 INVxp33_ASAP7_75t_R g43905 (.A(n_1127),
    .Y(n_1126));
 OR4x1_ASAP7_75t_R g43906 (.A(u4_n_1794),
    .B(u4_n_1795),
    .C(n_1010),
    .D(n_1068),
    .Y(n_1124));
 OAI21xp33_ASAP7_75t_R g43908 (.A1(opb_r[27]),
    .A2(n_45),
    .B(n_1088),
    .Y(n_1123));
 NOR3xp33_ASAP7_75t_R g43909 (.A(u1_n_68),
    .B(opb_r[23]),
    .C(opa_r[23]),
    .Y(n_1128));
 XOR2xp5_ASAP7_75t_R g43910 (.A(n_1078),
    .B(opa_r[24]),
    .Y(n_1122));
 MAJIxp5_ASAP7_75t_R g43911 (.A(n_1078),
    .B(n_71),
    .C(n_1046),
    .Y(n_1127));
 AND2x2_ASAP7_75t_R g43912 (.A(u1_fracta_s[26]),
    .B(u1_n_68),
    .Y(n_1125));
 NAND2xp33_ASAP7_75t_R g43913 (.A(div_opa_ldz_r2[0]),
    .B(u4_sll_315_50_n_29),
    .Y(n_3720));
 INVxp33_ASAP7_75t_R g43914 (.A(div_opa_ldz_r1[3]),
    .Y(n_1121));
 INVxp33_ASAP7_75t_R g43915 (.A(div_opa_ldz_r1[2]),
    .Y(n_1120));
 INVxp33_ASAP7_75t_R g43916 (.A(n_3507),
    .Y(n_1119));
 INVxp33_ASAP7_75t_R g43917 (.A(div_opa_ldz_r2[0]),
    .Y(n_1117));
 INVxp33_ASAP7_75t_R g43918 (.A(u1_n_68),
    .Y(n_1116));
 AOI222xp33_ASAP7_75t_R g43919 (.A1(n_676),
    .A2(quo[33]),
    .B1(n_652),
    .B2(fract_out_q[11]),
    .C1(n_1060),
    .C2(quo[10]),
    .Y(n_1115));
 AOI222xp33_ASAP7_75t_R g43922 (.A1(n_1059),
    .A2(quo[42]),
    .B1(n_653),
    .B2(fract_out_q[20]),
    .C1(n_665),
    .C2(quo[19]),
    .Y(n_1114));
 AOI222xp33_ASAP7_75t_R g43923 (.A1(n_677),
    .A2(quo[41]),
    .B1(n_653),
    .B2(fract_out_q[19]),
    .C1(n_665),
    .C2(quo[18]),
    .Y(n_1113));
 AOI222xp33_ASAP7_75t_R g43924 (.A1(n_678),
    .A2(quo[29]),
    .B1(n_652),
    .B2(fract_out_q[7]),
    .C1(n_665),
    .C2(quo[6]),
    .Y(n_1112));
 AOI222xp33_ASAP7_75t_R g43925 (.A1(n_1059),
    .A2(quo[30]),
    .B1(n_652),
    .B2(fract_out_q[8]),
    .C1(n_1060),
    .C2(quo[7]),
    .Y(n_1111));
 AOI222xp33_ASAP7_75t_R g43926 (.A1(n_677),
    .A2(quo[27]),
    .B1(n_653),
    .B2(fract_out_q[5]),
    .C1(n_1060),
    .C2(quo[4]),
    .Y(n_1110));
 AOI222xp33_ASAP7_75t_R g43927 (.A1(n_1060),
    .A2(quo[3]),
    .B1(n_678),
    .B2(quo[26]),
    .C1(n_652),
    .C2(fract_out_q[4]),
    .Y(n_1109));
 AOI222xp33_ASAP7_75t_R g43928 (.A1(n_678),
    .A2(quo[40]),
    .B1(n_652),
    .B2(fract_out_q[18]),
    .C1(n_1060),
    .C2(quo[17]),
    .Y(n_1108));
 AOI222xp33_ASAP7_75t_R g43929 (.A1(n_1059),
    .A2(quo[28]),
    .B1(n_653),
    .B2(fract_out_q[6]),
    .C1(n_665),
    .C2(quo[5]),
    .Y(n_1107));
 OAI31xp33_ASAP7_75t_R g43930 (.A1(n_3500),
    .A2(n_3715),
    .A3(n_1057),
    .B(n_24),
    .Y(n_3755));
 NAND2xp33_ASAP7_75t_R g43931 (.A(div_opa_ldz_r2[4]),
    .B(n_790),
    .Y(n_3507));
 NOR2xp33_ASAP7_75t_R g43932 (.A(opa_r1[8]),
    .B(n_1081),
    .Y(n_1118));
 NAND2xp33_ASAP7_75t_R g43933 (.A(n_1080),
    .B(exp_r[4]),
    .Y(n_3583));
 NAND2xp33_ASAP7_75t_R g43934 (.A(n_1084),
    .B(n_1082),
    .Y(u1_fracta_s[26]));
 NAND2xp33_ASAP7_75t_R g43937 (.A(n_1085),
    .B(n_1083),
    .Y(u1_n_68));
 AOI222xp33_ASAP7_75t_R g43938 (.A1(n_676),
    .A2(quo[34]),
    .B1(n_652),
    .B2(fract_out_q[12]),
    .C1(n_1060),
    .C2(quo[11]),
    .Y(n_1106));
 AOI222xp33_ASAP7_75t_R g43939 (.A1(n_678),
    .A2(quo[44]),
    .B1(n_652),
    .B2(fract_out_q[22]),
    .C1(n_1060),
    .C2(quo[21]),
    .Y(n_1105));
 AOI222xp33_ASAP7_75t_R g43940 (.A1(n_677),
    .A2(quo[35]),
    .B1(n_653),
    .B2(fract_out_q[13]),
    .C1(n_1060),
    .C2(quo[12]),
    .Y(n_1104));
 AOI222xp33_ASAP7_75t_R g43941 (.A1(n_676),
    .A2(quo[32]),
    .B1(n_653),
    .B2(fract_out_q[10]),
    .C1(n_1060),
    .C2(quo[9]),
    .Y(n_1103));
 AOI222xp33_ASAP7_75t_R g43942 (.A1(n_678),
    .A2(quo[39]),
    .B1(n_653),
    .B2(fract_out_q[17]),
    .C1(n_1060),
    .C2(quo[16]),
    .Y(n_1102));
 AOI222xp33_ASAP7_75t_R g43943 (.A1(n_676),
    .A2(quo[49]),
    .B1(n_652),
    .B2(fract_out_q[27]),
    .C1(n_665),
    .C2(quo[26]),
    .Y(n_1101));
 AOI222xp33_ASAP7_75t_R g43944 (.A1(n_1060),
    .A2(quo[0]),
    .B1(n_1059),
    .B2(quo[23]),
    .C1(n_653),
    .C2(fract_out_q[1]),
    .Y(n_1100));
 AOI222xp33_ASAP7_75t_R g43945 (.A1(n_678),
    .A2(quo[36]),
    .B1(n_652),
    .B2(fract_out_q[14]),
    .C1(n_1060),
    .C2(quo[13]),
    .Y(n_1099));
 AO222x2_ASAP7_75t_R g43946 (.A1(n_679),
    .A2(fract_i2f[0]),
    .B1(n_671),
    .B2(prod[0]),
    .C1(quo[2]),
    .C2(n_678),
    .Y(n_1098));
 AOI222xp33_ASAP7_75t_R g43947 (.A1(n_1059),
    .A2(quo[43]),
    .B1(n_653),
    .B2(fract_out_q[21]),
    .C1(n_665),
    .C2(quo[20]),
    .Y(n_1097));
 AOI222xp33_ASAP7_75t_R g43948 (.A1(n_677),
    .A2(quo[31]),
    .B1(n_653),
    .B2(fract_out_q[9]),
    .C1(n_665),
    .C2(quo[8]),
    .Y(n_1096));
 AOI222xp33_ASAP7_75t_R g43949 (.A1(n_665),
    .A2(quo[1]),
    .B1(n_678),
    .B2(quo[24]),
    .C1(n_653),
    .C2(fract_out_q[2]),
    .Y(n_1095));
 AOI222xp33_ASAP7_75t_R g43950 (.A1(n_1059),
    .A2(quo[38]),
    .B1(n_652),
    .B2(fract_out_q[16]),
    .C1(n_665),
    .C2(quo[15]),
    .Y(n_1094));
 AOI222xp33_ASAP7_75t_R g43951 (.A1(n_677),
    .A2(quo[37]),
    .B1(n_652),
    .B2(fract_out_q[15]),
    .C1(n_665),
    .C2(quo[14]),
    .Y(n_1093));
 AOI222xp33_ASAP7_75t_R g43952 (.A1(n_1059),
    .A2(quo[46]),
    .B1(n_653),
    .B2(fract_out_q[24]),
    .C1(n_665),
    .C2(quo[23]),
    .Y(n_1092));
 AOI222xp33_ASAP7_75t_R g43953 (.A1(n_676),
    .A2(quo[48]),
    .B1(n_653),
    .B2(fract_out_q[26]),
    .C1(n_665),
    .C2(quo[25]),
    .Y(n_1091));
 AOI222xp33_ASAP7_75t_R g43954 (.A1(n_665),
    .A2(quo[2]),
    .B1(n_678),
    .B2(quo[25]),
    .C1(n_652),
    .C2(fract_out_q[3]),
    .Y(n_1090));
 XNOR2xp5_ASAP7_75t_R g43955 (.A(n_1073),
    .B(opa_r1[7]),
    .Y(n_1089));
 MAJIxp5_ASAP7_75t_R g43956 (.A(n_1064),
    .B(n_795),
    .C(opa_r[26]),
    .Y(n_1088));
 INVxp33_ASAP7_75t_R g43957 (.A(div_opa_ldz_r1[0]),
    .Y(n_1087));
 INVxp33_ASAP7_75t_R g43958 (.A(div_opa_ldz_r1[1]),
    .Y(n_1086));
 INVxp33_ASAP7_75t_R g43959 (.A(n_1084),
    .Y(n_1085));
 INVxp33_ASAP7_75t_R g43960 (.A(n_1082),
    .Y(n_1083));
 INVxp33_ASAP7_75t_R g43962 (.A(div_opa_ldz_r2[4]),
    .Y(n_1080));
 NAND4xp25_ASAP7_75t_R g43965 (.A(n_1027),
    .B(n_3844),
    .C(n_2950),
    .D(n_3053),
    .Y(n_1079));
 NOR5xp2_ASAP7_75t_R g43966 (.A(n_1006),
    .B(opa_r[23]),
    .C(opa_r[30]),
    .D(opa_r[25]),
    .E(opa_r[26]),
    .Y(n_1084));
 NOR5xp2_ASAP7_75t_R g43967 (.A(n_1008),
    .B(opb_r[23]),
    .C(opb_r[24]),
    .D(opb_r[26]),
    .E(opb_r[25]),
    .Y(n_1082));
 NAND2xp33_ASAP7_75t_R g43968 (.A(n_800),
    .B(n_1073),
    .Y(n_1081));
 INVxp33_ASAP7_75t_R g43970 (.A(n_1076),
    .Y(n_3772));
 AND5x1_ASAP7_75t_R g43971 (.A(n_1005),
    .B(n_14294),
    .C(n_14293),
    .D(n_3053),
    .E(n_3052),
    .Y(n_1075));
 MAJIxp5_ASAP7_75t_R g43973 (.A(n_1054),
    .B(opa_r[23]),
    .C(n_656),
    .Y(n_1078));
 XOR2xp5_ASAP7_75t_R g43974 (.A(n_1042),
    .B(n_1054),
    .Y(u2_exp_tmp1[0]));
 OAI21xp33_ASAP7_75t_R g43975 (.A1(n_792),
    .A2(n_1056),
    .B(n_1034),
    .Y(n_3811));
 NOR5xp2_ASAP7_75t_R g43976 (.A(n_1004),
    .B(opa_r1[28]),
    .C(opa_r1[27]),
    .D(opa_r1[29]),
    .E(opa_r1[30]),
    .Y(n_1077));
 XNOR2xp5_ASAP7_75t_R g43977 (.A(n_3504),
    .B(n_24),
    .Y(n_1076));
 INVxp33_ASAP7_75t_R g43978 (.A(div_opa_ldz_r1[4]),
    .Y(n_1074));
 NAND5xp2_ASAP7_75t_R g43979 (.A(n_1015),
    .B(n_1016),
    .C(n_3846),
    .D(n_14293),
    .E(n_3034),
    .Y(n_1072));
 NAND4xp25_ASAP7_75t_R g43980 (.A(n_1009),
    .B(n_1016),
    .C(n_3543),
    .D(n_3052),
    .Y(n_1071));
 NOR2xp33_ASAP7_75t_R g43982 (.A(n_1019),
    .B(n_3801),
    .Y(n_3596));
 AOI21xp33_ASAP7_75t_R g43983 (.A1(n_1034),
    .A2(exp_r[7]),
    .B(n_36),
    .Y(n_1070));
 OAI311xp33_ASAP7_75t_R g43984 (.A1(n_991),
    .A2(n_13946),
    .A3(exp_r[6]),
    .B1(exp_r[7]),
    .C1(n_997),
    .Y(n_3754));
 OR2x2_ASAP7_75t_R g43985 (.A(n_24),
    .B(n_3504),
    .Y(n_3573));
 NOR2xp33_ASAP7_75t_R g43986 (.A(opa_r1[6]),
    .B(n_1061),
    .Y(n_1073));
 OAI21xp33_ASAP7_75t_R g43987 (.A1(n_13946),
    .A2(n_1035),
    .B(n_3564),
    .Y(n_3816));
 OR5x1_ASAP7_75t_R g43989 (.A(u4_n_1812),
    .B(u4_n_1801),
    .C(u4_n_1809),
    .D(n_987),
    .E(n_1011),
    .Y(n_1068));
 AOI22xp33_ASAP7_75t_R g43990 (.A1(prod[43]),
    .A2(n_671),
    .B1(fract_out_q[23]),
    .B2(n_653),
    .Y(n_1067));
 AOI22xp33_ASAP7_75t_R g43991 (.A1(prod[20]),
    .A2(n_672),
    .B1(fract_out_q[0]),
    .B2(n_652),
    .Y(n_1066));
 AOI22xp33_ASAP7_75t_R g43992 (.A1(prod[45]),
    .A2(n_23),
    .B1(fract_out_q[25]),
    .B2(n_652),
    .Y(n_1065));
 MAJIxp5_ASAP7_75t_R g43993 (.A(n_1025),
    .B(opb_r[25]),
    .C(n_44),
    .Y(n_1064));
 XNOR2xp5_ASAP7_75t_R g43994 (.A(n_1039),
    .B(opa_r1[5]),
    .Y(n_1063));
 XNOR2xp5_ASAP7_75t_R g43995 (.A(n_1037),
    .B(n_700),
    .Y(n_3753));
 XNOR2xp5_ASAP7_75t_R g43996 (.A(n_1038),
    .B(n_792),
    .Y(n_3773));
 XNOR2xp5_ASAP7_75t_R g43997 (.A(n_1036),
    .B(n_700),
    .Y(n_3775));
 INVxp33_ASAP7_75t_R g43998 (.A(n_36),
    .Y(n_3502));
 AND4x1_ASAP7_75t_R g44001 (.A(n_986),
    .B(n_3844),
    .C(n_3849),
    .D(n_2950),
    .Y(n_1058));
 NOR2xp33_ASAP7_75t_R g44002 (.A(n_67),
    .B(n_13972),
    .Y(n_1057));
 NOR2xp33_ASAP7_75t_R g44003 (.A(n_13946),
    .B(n_1035),
    .Y(n_1056));
 OR2x2_ASAP7_75t_R g44004 (.A(n_24),
    .B(n_1034),
    .Y(n_3503));
 NOR2xp33_ASAP7_75t_R g44005 (.A(n_682),
    .B(n_1029),
    .Y(n_3599));
 NAND2xp33_ASAP7_75t_R g44006 (.A(exp_r[5]),
    .B(n_1035),
    .Y(n_3564));
 NOR2xp33_ASAP7_75t_R g44007 (.A(exp_r[7]),
    .B(n_1034),
    .Y(n_36));
 NAND2xp33_ASAP7_75t_R g44008 (.A(n_798),
    .B(n_1039),
    .Y(n_1061));
 NAND2xp33_ASAP7_75t_R g44009 (.A(n_3850),
    .B(u4_n_1362),
    .Y(n_3801));
 NAND2xp33_ASAP7_75t_R g44010 (.A(exp_r[6]),
    .B(n_1038),
    .Y(n_3504));
 NOR2xp33_ASAP7_75t_R g44011 (.A(opb_dn),
    .B(n_13919),
    .Y(n_1060));
 AND2x2_ASAP7_75t_R g44012 (.A(opb_dn),
    .B(n_22),
    .Y(n_1059));
 INVxp33_ASAP7_75t_R g44013 (.A(n_3826),
    .Y(n_1055));
 INVxp33_ASAP7_75t_R g44015 (.A(n_1051),
    .Y(n_1050));
 INVxp33_ASAP7_75t_R g44017 (.A(n_1047),
    .Y(n_1048));
 INVxp33_ASAP7_75t_R g44018 (.A(n_1044),
    .Y(n_1045));
 AOI21xp33_ASAP7_75t_R g44020 (.A1(n_1021),
    .A2(n_790),
    .B(n_1037),
    .Y(n_3752));
 OAI22xp33_ASAP7_75t_R g44022 (.A1(opa_r[23]),
    .A2(u2_n_606),
    .B1(n_54),
    .B2(n_656),
    .Y(n_1042));
 OAI21xp33_ASAP7_75t_R g44023 (.A1(n_790),
    .A2(n_1018),
    .B(n_1035),
    .Y(n_3826));
 OAI22xp33_ASAP7_75t_R g44024 (.A1(opb_r[23]),
    .A2(u2_n_606),
    .B1(n_796),
    .B2(n_656),
    .Y(n_1054));
 AOI21xp33_ASAP7_75t_R g44025 (.A1(u2_n_606),
    .A2(opb_r[30]),
    .B(n_1040),
    .Y(n_1053));
 AOI22xp33_ASAP7_75t_R g44026 (.A1(n_795),
    .A2(n_656),
    .B1(opb_r[26]),
    .B2(n_13981),
    .Y(n_1052));
 OAI22xp33_ASAP7_75t_R g44027 (.A1(opb_r[25]),
    .A2(u2_n_606),
    .B1(n_713),
    .B2(n_656),
    .Y(n_1051));
 OAI22xp33_ASAP7_75t_R g44028 (.A1(opb_r[27]),
    .A2(u2_n_606),
    .B1(n_717),
    .B2(n_656),
    .Y(n_1049));
 AOI22xp33_ASAP7_75t_R g44029 (.A1(n_714),
    .A2(n_656),
    .B1(opb_r[29]),
    .B2(n_13981),
    .Y(n_1047));
 AOI22xp33_ASAP7_75t_R g44030 (.A1(n_715),
    .A2(n_656),
    .B1(opb_r[24]),
    .B2(u2_n_606),
    .Y(n_1046));
 AOI22xp33_ASAP7_75t_R g44031 (.A1(n_712),
    .A2(n_656),
    .B1(opb_r[28]),
    .B2(n_13981),
    .Y(n_1044));
 INVxp33_ASAP7_75t_R g44033 (.A(n_67),
    .Y(n_3756));
 NAND2xp33_ASAP7_75t_R g44034 (.A(opa_r1[0]),
    .B(n_621),
    .Y(n_1033));
 NOR2xp33_ASAP7_75t_R g44035 (.A(rmode_r3[0]),
    .B(rmode_r3[1]),
    .Y(n_67));
 NOR2xp33_ASAP7_75t_R g44036 (.A(opb_r[30]),
    .B(u2_n_606),
    .Y(n_1040));
 NOR2xp33_ASAP7_75t_R g44037 (.A(opa_r1[4]),
    .B(n_1023),
    .Y(n_1039));
 NOR2xp33_ASAP7_75t_R g44038 (.A(n_3774),
    .B(n_1022),
    .Y(n_1038));
 NOR2xp33_ASAP7_75t_R g44039 (.A(n_790),
    .B(n_1021),
    .Y(n_1037));
 NOR2xp33_ASAP7_75t_R g44040 (.A(n_790),
    .B(n_1022),
    .Y(n_1036));
 NAND2xp33_ASAP7_75t_R g44041 (.A(n_790),
    .B(n_1018),
    .Y(n_1035));
 NAND2xp33_ASAP7_75t_R g44042 (.A(n_998),
    .B(n_1018),
    .Y(n_1034));
 INVxp33_ASAP7_75t_R g44043 (.A(n_1028),
    .Y(n_1032));
 INVxp33_ASAP7_75t_R g44046 (.A(u4_n_1362),
    .Y(n_1029));
 OAI32xp33_ASAP7_75t_R g44053 (.A1(n_879),
    .A2(n_717),
    .A3(opa_r[27]),
    .B1(n_712),
    .B2(opa_r[28]),
    .Y(n_1028));
 AND3x1_ASAP7_75t_R g44054 (.A(n_1015),
    .B(n_999),
    .C(n_3020),
    .Y(n_1027));
 OA21x2_ASAP7_75t_R g44055 (.A1(exp_r[3]),
    .A2(n_995),
    .B(n_1021),
    .Y(n_3751));
 XNOR2xp5_ASAP7_75t_R g44056 (.A(n_14564),
    .B(opa_r1[3]),
    .Y(n_1026));
 AOI32xp33_ASAP7_75t_R g44057 (.A1(n_872),
    .A2(n_796),
    .A3(opa_r[23]),
    .B1(n_715),
    .B2(opa_r[24]),
    .Y(n_1025));
 AO21x1_ASAP7_75t_R g44058 (.A1(exp_r[3]),
    .A2(n_992),
    .B(n_1018),
    .Y(n_3822));
 XNOR2xp5_ASAP7_75t_R g44059 (.A(n_3769),
    .B(exp_r[3]),
    .Y(n_3768));
 NAND3xp33_ASAP7_75t_R g44060 (.A(n_47),
    .B(fpu_op_r3[1]),
    .C(fpu_op_r3[0]),
    .Y(u4_n_1362));
 INVxp33_ASAP7_75t_R g44062 (.A(n_1024),
    .Y(n_3527));
 INVxp33_ASAP7_75t_R g44064 (.A(n_1020),
    .Y(u4_op_dn));
 NAND2xp33_ASAP7_75t_R g44066 (.A(n_998),
    .B(n_24),
    .Y(n_3501));
 NAND2xp33_ASAP7_75t_R g44067 (.A(rmode_r2[1]),
    .B(rmode_r2[0]),
    .Y(n_1017));
 NOR2xp33_ASAP7_75t_R g44069 (.A(opa_dn),
    .B(n_989),
    .Y(n_1024));
 NAND2xp33_ASAP7_75t_R g44070 (.A(opa_dn),
    .B(opb_dn),
    .Y(n_3528));
 OR2x2_ASAP7_75t_R g44071 (.A(fpu_op_r3[0]),
    .B(n_3497),
    .Y(n_3594));
 NAND2xp33_ASAP7_75t_R g44073 (.A(n_797),
    .B(n_14564),
    .Y(n_1023));
 NAND2xp33_ASAP7_75t_R g44074 (.A(n_991),
    .B(exp_r[0]),
    .Y(n_1022));
 NAND2xp33_ASAP7_75t_R g44075 (.A(exp_r[3]),
    .B(n_995),
    .Y(n_1021));
 NOR2xp33_ASAP7_75t_R g44076 (.A(opa_dn),
    .B(opb_dn),
    .Y(n_1020));
 NAND2xp33_ASAP7_75t_R g44077 (.A(fpu_op_r3[0]),
    .B(n_682),
    .Y(n_3803));
 NOR2xp33_ASAP7_75t_R g44078 (.A(exp_r[3]),
    .B(n_992),
    .Y(n_1018));
 NAND2xp33_ASAP7_75t_R g44080 (.A(n_3497),
    .B(fpu_op_r3[2]),
    .Y(n_1602));
 INVxp33_ASAP7_75t_R g44081 (.A(n_1014),
    .Y(n_3771));
 INVxp33_ASAP7_75t_R g44086 (.A(n_13981),
    .Y(n_683));
 INVxp33_ASAP7_75t_R g44089 (.A(n_656),
    .Y(u2_n_606));
 OR5x1_ASAP7_75t_R g44099 (.A(u4_n_1814),
    .B(u4_n_1813),
    .C(u4_n_1816),
    .D(u4_n_1811),
    .E(u4_n_1800),
    .Y(n_1011));
 OR5x1_ASAP7_75t_R g44100 (.A(u4_n_1810),
    .B(u4_n_1799),
    .C(u4_n_1806),
    .D(u4_n_1797),
    .E(u4_n_1804),
    .Y(n_1010));
 AOI211xp5_ASAP7_75t_R g44101 (.A1(u4_n_1847),
    .A2(u4_n_1848),
    .B(u4_n_1850),
    .C(u4_n_1849),
    .Y(u4_round2a_BAR));
 AND3x1_ASAP7_75t_R g44102 (.A(n_999),
    .B(n_3847),
    .C(n_2935),
    .Y(n_1009));
 OR4x1_ASAP7_75t_R g44103 (.A(opb_r[27]),
    .B(opb_r[28]),
    .C(opb_r[29]),
    .D(opb_r[30]),
    .Y(n_1008));
 XNOR2xp5_ASAP7_75t_R g44104 (.A(n_14033),
    .B(opa_r1[2]),
    .Y(n_1007));
 OR4x1_ASAP7_75t_R g44105 (.A(opa_r[24]),
    .B(opa_r[27]),
    .C(opa_r[29]),
    .D(opa_r[28]),
    .Y(n_1006));
 AND4x1_ASAP7_75t_R g44106 (.A(n_3541),
    .B(n_3543),
    .C(n_3055),
    .D(n_3045),
    .Y(n_1005));
 OR4x1_ASAP7_75t_R g44107 (.A(opa_r1[23]),
    .B(opa_r1[24]),
    .C(opa_r1[26]),
    .D(opa_r1[25]),
    .Y(n_1004));
 NAND2xp33_ASAP7_75t_R g44108 (.A(u1_exp_large[7]),
    .B(n_1001),
    .Y(u1_n_5489));
 AND4x1_ASAP7_75t_R g44109 (.A(n_3845),
    .B(n_2950),
    .C(n_3055),
    .D(n_3840),
    .Y(n_1016));
 AND4x1_ASAP7_75t_R g44110 (.A(n_3849),
    .B(n_3045),
    .C(n_3052),
    .D(n_802),
    .Y(n_1015));
 NAND2xp33_ASAP7_75t_R g44111 (.A(n_994),
    .B(n_992),
    .Y(n_3824));
 OAI21xp33_ASAP7_75t_R g44112 (.A1(exp_r[2]),
    .A2(n_876),
    .B(n_3769),
    .Y(n_1014));
 NAND3xp33_ASAP7_75t_R g44113 (.A(n_801),
    .B(fpu_op_r2[2]),
    .C(fpu_op_r2[0]),
    .Y(n_3499));
 AND3x1_ASAP7_75t_R g44114 (.A(fpu_op_r1[0]),
    .B(n_56),
    .C(fpu_op_r1[1]),
    .Y(n_656));
 INVxp33_ASAP7_75t_R g44115 (.A(rmode_r2[1]),
    .Y(n_1003));
 INVxp33_ASAP7_75t_R g44116 (.A(opas_r2),
    .Y(n_1002));
 INVxp33_ASAP7_75t_R g44177 (.A(n_998),
    .Y(n_997));
 INVxp33_ASAP7_75t_R g44178 (.A(rmode_r2[0]),
    .Y(n_996));
 INVxp33_ASAP7_75t_R g44179 (.A(n_995),
    .Y(n_994));
 INVxp33_ASAP7_75t_R g44180 (.A(n_991),
    .Y(n_3715));
 INVxp33_ASAP7_75t_R g44183 (.A(opb_dn),
    .Y(n_989));
 XOR2xp5_ASAP7_75t_R g44193 (.A(opa_r1[0]),
    .B(opa_r1[1]),
    .Y(n_988));
 OR4x1_ASAP7_75t_R g44199 (.A(u4_n_1808),
    .B(u4_n_1807),
    .C(u4_n_1802),
    .D(u4_n_1815),
    .Y(n_987));
 AND3x1_ASAP7_75t_R g44201 (.A(n_3848),
    .B(n_3070),
    .C(n_3845),
    .Y(n_986));
 OR2x2_ASAP7_75t_R g44202 (.A(n_62),
    .B(n_878),
    .Y(n_1001));
 AO21x1_ASAP7_75t_R g44234 (.A1(opa_r[29]),
    .A2(n_714),
    .B(n_878),
    .Y(n_1000));
 AND3x1_ASAP7_75t_R g44236 (.A(n_3070),
    .B(n_14294),
    .C(n_2928),
    .Y(n_999));
 OR2x2_ASAP7_75t_R g44238 (.A(n_792),
    .B(n_3774),
    .Y(n_3500));
 NOR3xp33_ASAP7_75t_R g44239 (.A(n_13946),
    .B(exp_r[4]),
    .C(exp_r[6]),
    .Y(n_998));
 NOR2xp33_ASAP7_75t_R g44241 (.A(n_706),
    .B(n_877),
    .Y(n_995));
 NAND2xp33_ASAP7_75t_R g44243 (.A(n_706),
    .B(n_877),
    .Y(n_992));
 NAND2xp33_ASAP7_75t_R g44244 (.A(exp_r[2]),
    .B(n_876),
    .Y(n_3769));
 NOR2xp33_ASAP7_75t_R g44245 (.A(n_43),
    .B(n_3716),
    .Y(n_991));
 OR2x2_ASAP7_75t_R g44246 (.A(n_876),
    .B(n_877),
    .Y(n_3820));
 NOR2xp33_ASAP7_75t_R g44249 (.A(fpu_op_r3[1]),
    .B(n_47),
    .Y(n_682));
 INVxp33_ASAP7_75t_R g44250 (.A(u6_quo1[36]),
    .Y(n_985));
 INVxp33_ASAP7_75t_R g44251 (.A(u6_quo1[24]),
    .Y(n_984));
 INVxp33_ASAP7_75t_R g44252 (.A(u5_prod1[39]),
    .Y(n_983));
 INVxp33_ASAP7_75t_R g44253 (.A(u6_quo1[16]),
    .Y(n_982));
 INVxp33_ASAP7_75t_R g44254 (.A(u6_quo1[42]),
    .Y(n_981));
 INVxp33_ASAP7_75t_R g44255 (.A(u5_prod1[23]),
    .Y(n_980));
 INVxp33_ASAP7_75t_R g44256 (.A(u5_prod1[37]),
    .Y(n_979));
 INVxp33_ASAP7_75t_R g44257 (.A(u5_prod1[5]),
    .Y(n_978));
 INVxp33_ASAP7_75t_R g44258 (.A(u6_quo1[3]),
    .Y(n_977));
 INVxp33_ASAP7_75t_R g44259 (.A(u6_quo1[12]),
    .Y(n_976));
 INVxp33_ASAP7_75t_R g44260 (.A(u6_quo1[33]),
    .Y(n_975));
 INVxp33_ASAP7_75t_R g44261 (.A(u6_quo1[40]),
    .Y(n_974));
 INVxp33_ASAP7_75t_R g44262 (.A(u5_prod1[17]),
    .Y(n_973));
 INVxp33_ASAP7_75t_R g44263 (.A(u6_quo1[6]),
    .Y(n_972));
 INVxp33_ASAP7_75t_R g44264 (.A(u6_quo1[11]),
    .Y(n_971));
 INVxp33_ASAP7_75t_R g44265 (.A(u5_prod1[20]),
    .Y(n_970));
 INVxp33_ASAP7_75t_R g44266 (.A(u6_quo1[47]),
    .Y(n_969));
 INVxp33_ASAP7_75t_R g44267 (.A(u5_prod1[44]),
    .Y(n_968));
 INVxp33_ASAP7_75t_R g44268 (.A(u6_quo1[15]),
    .Y(n_967));
 INVxp33_ASAP7_75t_R g44269 (.A(u5_prod1[2]),
    .Y(n_966));
 INVxp33_ASAP7_75t_R g44270 (.A(u5_prod1[35]),
    .Y(n_965));
 INVxp33_ASAP7_75t_R g44271 (.A(u6_quo1[25]),
    .Y(n_964));
 INVxp33_ASAP7_75t_R g44272 (.A(u6_quo1[30]),
    .Y(n_963));
 INVxp33_ASAP7_75t_R g44273 (.A(u6_quo1[27]),
    .Y(n_962));
 INVxp33_ASAP7_75t_R g44274 (.A(u6_quo1[29]),
    .Y(n_961));
 INVxp33_ASAP7_75t_R g44275 (.A(u6_quo1[5]),
    .Y(n_960));
 INVxp33_ASAP7_75t_R g44276 (.A(u6_quo1[48]),
    .Y(n_959));
 INVxp33_ASAP7_75t_R g44277 (.A(u6_quo1[34]),
    .Y(n_958));
 INVxp33_ASAP7_75t_R g44278 (.A(u5_prod1[47]),
    .Y(n_957));
 INVxp33_ASAP7_75t_R g44279 (.A(u6_quo1[19]),
    .Y(n_956));
 INVxp33_ASAP7_75t_R g44280 (.A(u6_quo1[35]),
    .Y(n_955));
 INVxp33_ASAP7_75t_R g44281 (.A(u5_prod1[22]),
    .Y(n_954));
 INVxp33_ASAP7_75t_R g44282 (.A(u6_quo1[22]),
    .Y(n_953));
 INVxp33_ASAP7_75t_R g44283 (.A(u5_prod1[15]),
    .Y(n_952));
 INVxp33_ASAP7_75t_R g44284 (.A(u6_quo1[4]),
    .Y(n_951));
 INVxp33_ASAP7_75t_R g44285 (.A(u6_quo1[44]),
    .Y(n_950));
 INVxp33_ASAP7_75t_R g44286 (.A(u5_prod1[4]),
    .Y(n_949));
 INVxp33_ASAP7_75t_R g44287 (.A(u6_quo1[9]),
    .Y(n_948));
 INVxp33_ASAP7_75t_R g44288 (.A(u6_quo1[49]),
    .Y(n_947));
 INVxp33_ASAP7_75t_R g44289 (.A(u6_quo1[46]),
    .Y(n_946));
 INVxp33_ASAP7_75t_R g44290 (.A(u5_prod1[0]),
    .Y(n_945));
 INVxp33_ASAP7_75t_R g44291 (.A(u6_quo1[17]),
    .Y(n_944));
 INVxp33_ASAP7_75t_R g44292 (.A(u5_prod1[40]),
    .Y(n_943));
 INVxp33_ASAP7_75t_R g44293 (.A(rmode_r1[1]),
    .Y(n_942));
 INVxp33_ASAP7_75t_R g44294 (.A(u5_prod1[33]),
    .Y(n_941));
 INVxp33_ASAP7_75t_R g44295 (.A(rmode_r1[0]),
    .Y(n_940));
 INVxp33_ASAP7_75t_R g44297 (.A(u5_prod1[46]),
    .Y(n_938));
 INVxp33_ASAP7_75t_R g44298 (.A(u5_prod1[45]),
    .Y(n_937));
 INVxp33_ASAP7_75t_R g44299 (.A(u6_quo1[41]),
    .Y(n_936));
 INVxp33_ASAP7_75t_R g44300 (.A(u5_prod1[11]),
    .Y(n_935));
 INVxp33_ASAP7_75t_R g44301 (.A(u5_prod1[27]),
    .Y(n_934));
 INVxp33_ASAP7_75t_R g44302 (.A(u5_prod1[12]),
    .Y(n_933));
 INVxp33_ASAP7_75t_R g44303 (.A(u5_prod1[24]),
    .Y(n_932));
 INVxp33_ASAP7_75t_R g44304 (.A(u5_prod1[43]),
    .Y(n_931));
 INVxp33_ASAP7_75t_R g44305 (.A(u5_prod1[31]),
    .Y(n_930));
 INVxp33_ASAP7_75t_R g44306 (.A(u6_quo1[14]),
    .Y(n_929));
 INVxp33_ASAP7_75t_R g44307 (.A(u5_prod1[7]),
    .Y(n_928));
 INVxp33_ASAP7_75t_R g44308 (.A(u5_prod1[28]),
    .Y(n_927));
 INVxp33_ASAP7_75t_R g44309 (.A(fpu_op_r1[2]),
    .Y(n_56));
 INVxp33_ASAP7_75t_R g44310 (.A(fpu_op_r3[1]),
    .Y(n_925));
 INVxp33_ASAP7_75t_R g44311 (.A(fpu_op_r3[2]),
    .Y(n_47));
 INVxp33_ASAP7_75t_R g44385 (.A(u6_quo1[43]),
    .Y(n_923));
 INVxp33_ASAP7_75t_R g44386 (.A(u5_prod1[1]),
    .Y(n_922));
 INVxp33_ASAP7_75t_R g44387 (.A(u6_quo1[31]),
    .Y(n_921));
 INVxp33_ASAP7_75t_R g44388 (.A(u6_quo1[39]),
    .Y(n_920));
 INVxp33_ASAP7_75t_R g44389 (.A(u5_prod1[29]),
    .Y(n_919));
 INVxp33_ASAP7_75t_R g44390 (.A(u5_prod1[38]),
    .Y(n_918));
 INVxp33_ASAP7_75t_R g44391 (.A(u6_quo1[38]),
    .Y(n_917));
 INVxp33_ASAP7_75t_R g44392 (.A(u5_prod1[8]),
    .Y(n_916));
 INVxp33_ASAP7_75t_R g44393 (.A(u5_prod1[21]),
    .Y(n_915));
 INVxp33_ASAP7_75t_R g44394 (.A(u5_prod1[30]),
    .Y(n_914));
 INVxp33_ASAP7_75t_R g44395 (.A(u5_prod1[36]),
    .Y(n_913));
 INVxp33_ASAP7_75t_R g44396 (.A(u5_prod1[42]),
    .Y(n_912));
 INVxp33_ASAP7_75t_R g44397 (.A(u5_prod1[26]),
    .Y(n_911));
 INVxp33_ASAP7_75t_R g44398 (.A(u6_quo1[37]),
    .Y(n_910));
 INVxp33_ASAP7_75t_R g44399 (.A(u6_quo1[20]),
    .Y(n_909));
 INVxp33_ASAP7_75t_R g44400 (.A(u6_quo1[23]),
    .Y(n_908));
 INVxp33_ASAP7_75t_R g44401 (.A(u6_quo1[45]),
    .Y(n_907));
 INVxp33_ASAP7_75t_R g44402 (.A(u5_prod1[41]),
    .Y(n_906));
 INVxp33_ASAP7_75t_R g44403 (.A(u6_quo1[32]),
    .Y(n_905));
 INVxp33_ASAP7_75t_R g44404 (.A(u6_quo1[28]),
    .Y(n_904));
 INVxp33_ASAP7_75t_R g44405 (.A(u5_prod1[16]),
    .Y(n_903));
 INVxp33_ASAP7_75t_R g44406 (.A(u5_prod1[10]),
    .Y(n_902));
 INVxp33_ASAP7_75t_R g44407 (.A(u6_quo1[26]),
    .Y(n_901));
 INVxp33_ASAP7_75t_R g44408 (.A(u6_quo1[8]),
    .Y(n_900));
 INVxp33_ASAP7_75t_R g44410 (.A(u6_quo1[2]),
    .Y(n_898));
 INVxp33_ASAP7_75t_R g44411 (.A(u6_quo1[21]),
    .Y(n_897));
 INVxp33_ASAP7_75t_R g44412 (.A(u5_prod1[3]),
    .Y(n_896));
 INVxp33_ASAP7_75t_R g44413 (.A(u6_quo1[18]),
    .Y(n_895));
 INVxp33_ASAP7_75t_R g44414 (.A(u5_prod1[9]),
    .Y(n_894));
 INVxp33_ASAP7_75t_R g44415 (.A(u6_quo1[7]),
    .Y(n_893));
 INVxp33_ASAP7_75t_R g44416 (.A(u5_prod1[32]),
    .Y(n_892));
 INVxp33_ASAP7_75t_R g44417 (.A(u6_quo1[10]),
    .Y(n_891));
 INVxp33_ASAP7_75t_R g44418 (.A(u5_prod1[19]),
    .Y(n_890));
 INVxp33_ASAP7_75t_R g44419 (.A(u5_prod1[25]),
    .Y(n_889));
 INVxp33_ASAP7_75t_R g44420 (.A(u5_prod1[6]),
    .Y(n_888));
 INVxp33_ASAP7_75t_R g44421 (.A(u5_prod1[18]),
    .Y(n_887));
 INVxp33_ASAP7_75t_R g44422 (.A(u6_quo1[13]),
    .Y(n_886));
 INVxp33_ASAP7_75t_R g44423 (.A(u5_prod1[34]),
    .Y(n_885));
 INVxp33_ASAP7_75t_R g44424 (.A(opas_r1),
    .Y(n_884));
 INVxp33_ASAP7_75t_R g44425 (.A(u5_prod1[14]),
    .Y(n_883));
 INVxp33_ASAP7_75t_R g44426 (.A(u5_prod1[13]),
    .Y(n_882));
 INVxp33_ASAP7_75t_R g44427 (.A(u0_expb_00),
    .Y(n_881));
 INVxp33_ASAP7_75t_R g44428 (.A(u0_expa_00),
    .Y(n_880));
 INVxp33_ASAP7_75t_R g44429 (.A(fpu_op_r2[0]),
    .Y(n_875));
 NAND2xp33_ASAP7_75t_R g44445 (.A(opb_r[24]),
    .B(n_71),
    .Y(n_872));
 NAND2xp33_ASAP7_75t_R g44493 (.A(n_62),
    .B(n_718),
    .Y(u1_exp_large[7]));
 NOR2xp33_ASAP7_75t_R g44494 (.A(opb_r[28]),
    .B(n_49),
    .Y(n_879));
 NAND2xp33_ASAP7_75t_R g44495 (.A(opa_r[23]),
    .B(opb_r[23]),
    .Y(u1_n_8071));
 NAND2xp33_ASAP7_75t_R g44496 (.A(exp_r[1]),
    .B(exp_r[2]),
    .Y(n_3716));
 NAND2xp33_ASAP7_75t_R g44498 (.A(exp_r[4]),
    .B(exp_r[5]),
    .Y(n_3774));
 NOR2xp33_ASAP7_75t_R g44499 (.A(opb_r[30]),
    .B(n_62),
    .Y(n_878));
 NOR2xp33_ASAP7_75t_R g44500 (.A(exp_r[0]),
    .B(exp_r[1]),
    .Y(n_877));
 NOR2xp33_ASAP7_75t_R g44501 (.A(n_716),
    .B(u4_sll_315_50_n_29),
    .Y(n_876));
 INVxp33_ASAP7_75t_R g44505 (.A(u6_n_123),
    .Y(n_870));
 INVxp33_ASAP7_75t_R g44509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3619),
    .Y(n_866));
 INVxp33_ASAP7_75t_R g44519 (.A(u6_n_91),
    .Y(n_856));
 INVxp33_ASAP7_75t_R g44522 (.A(u6_n_99),
    .Y(n_853));
 INVxp33_ASAP7_75t_R g44523 (.A(u6_n_113),
    .Y(n_852));
 INVxp33_ASAP7_75t_R g44524 (.A(u6_n_95),
    .Y(n_851));
 INVxp33_ASAP7_75t_R g44526 (.A(u6_n_104),
    .Y(n_849));
 INVxp33_ASAP7_75t_R g44527 (.A(u6_n_108),
    .Y(n_848));
 INVxp33_ASAP7_75t_R g44528 (.A(u6_n_119),
    .Y(n_847));
 INVxp33_ASAP7_75t_R g44531 (.A(u6_n_83),
    .Y(n_844));
 INVxp33_ASAP7_75t_R g44536 (.A(u6_n_79),
    .Y(n_839));
 INVxp33_ASAP7_75t_R g44537 (.A(u6_n_112),
    .Y(n_838));
 INVxp33_ASAP7_75t_R g44541 (.A(fpu_op[1]),
    .Y(n_834));
 INVxp33_ASAP7_75t_R g44542 (.A(u6_n_111),
    .Y(n_833));
 INVxp33_ASAP7_75t_R g44545 (.A(u6_n_96),
    .Y(n_830));
 INVxp33_ASAP7_75t_R g44553 (.A(fpu_op[2]),
    .Y(n_822));
 INVxp33_ASAP7_75t_R g44558 (.A(u6_n_109),
    .Y(n_817));
 INVxp33_ASAP7_75t_R g44565 (.A(u6_n_116),
    .Y(n_810));
 INVxp33_ASAP7_75t_R g44566 (.A(u6_n_117),
    .Y(n_809));
 INVxp33_ASAP7_75t_R g44570 (.A(u6_n_84),
    .Y(n_805));
 INVxp33_ASAP7_75t_R g44574 (.A(fpu_op_r2[1]),
    .Y(n_801));
 INVxp33_ASAP7_75t_R g44575 (.A(opa_r1[7]),
    .Y(n_800));
 INVxp33_ASAP7_75t_R g44576 (.A(opa_r1[17]),
    .Y(n_799));
 INVxp33_ASAP7_75t_R g44577 (.A(opa_r1[5]),
    .Y(n_798));
 INVxp33_ASAP7_75t_R g44578 (.A(opa_r1[3]),
    .Y(n_797));
 INVxp33_ASAP7_75t_R g44579 (.A(opb_r[23]),
    .Y(n_796));
 INVxp33_ASAP7_75t_R g44580 (.A(opb_r[26]),
    .Y(n_795));
 INVxp33_ASAP7_75t_R g44581 (.A(opa_r[24]),
    .Y(n_71));
 INVxp33_ASAP7_75t_R g44582 (.A(opa_r[25]),
    .Y(n_44));
 INVxp33_ASAP7_75t_R g44583 (.A(exp_r[6]),
    .Y(n_792));
 INVxp33_ASAP7_75t_R g44584 (.A(opa_r[30]),
    .Y(n_62));
 INVxp33_ASAP7_75t_R g44585 (.A(exp_r[4]),
    .Y(n_790));
 INVxp33_ASAP7_75t_R g44586 (.A(exp_r[7]),
    .Y(n_24));
 INVxp33_ASAP7_75t_R g44601 (.A(u4_n_1852),
    .Y(n_774));
 INVxp33_ASAP7_75t_R g44604 (.A(u6_n_118),
    .Y(n_771));
 INVxp33_ASAP7_75t_R g44606 (.A(u6_n_101),
    .Y(n_769));
 INVxp33_ASAP7_75t_R g44612 (.A(u6_n_124),
    .Y(n_763));
 INVxp33_ASAP7_75t_R g44614 (.A(u6_n_120),
    .Y(n_761));
 INVxp33_ASAP7_75t_R g44624 (.A(fractb[0]),
    .Y(n_751));
 INVxp33_ASAP7_75t_R g44629 (.A(rmode[0]),
    .Y(n_746));
 INVxp33_ASAP7_75t_R g44632 (.A(rmode[1]),
    .Y(n_743));
 INVxp33_ASAP7_75t_R g44633 (.A(u5_n_2),
    .Y(n_742));
 INVxp33_ASAP7_75t_R g44635 (.A(u6_n_89),
    .Y(n_740));
 INVxp33_ASAP7_75t_R g44638 (.A(u6_n_87),
    .Y(n_737));
 INVxp33_ASAP7_75t_R g44642 (.A(u6_n_82),
    .Y(n_733));
 INVxp33_ASAP7_75t_R g44648 (.A(fpu_op_r2[2]),
    .Y(n_727));
 INVxp33_ASAP7_75t_R g44649 (.A(fpu_op_r1[0]),
    .Y(n_726));
 INVxp33_ASAP7_75t_R g44651 (.A(opa_r1[21]),
    .Y(n_724));
 INVxp33_ASAP7_75t_R g44652 (.A(opa_r1[13]),
    .Y(n_723));
 INVxp33_ASAP7_75t_R g44653 (.A(opa_r1[9]),
    .Y(n_722));
 INVxp33_ASAP7_75t_R g44654 (.A(opa_r1[19]),
    .Y(n_721));
 INVxp33_ASAP7_75t_R g44655 (.A(opa_r1[11]),
    .Y(n_720));
 INVxp33_ASAP7_75t_R g44656 (.A(opa_r1[15]),
    .Y(n_719));
 INVxp33_ASAP7_75t_R g44657 (.A(opb_r[30]),
    .Y(n_718));
 INVxp33_ASAP7_75t_R g44658 (.A(opb_r[27]),
    .Y(n_717));
 INVxp33_ASAP7_75t_R g44660 (.A(opb_r[24]),
    .Y(n_715));
 INVxp33_ASAP7_75t_R g44661 (.A(opb_r[29]),
    .Y(n_714));
 INVxp33_ASAP7_75t_R g44662 (.A(opb_r[25]),
    .Y(n_713));
 INVxp33_ASAP7_75t_R g44663 (.A(opb_r[28]),
    .Y(n_712));
 INVxp33_ASAP7_75t_R g44667 (.A(opa_r[26]),
    .Y(n_41));
 INVxp33_ASAP7_75t_R g44669 (.A(exp_r[2]),
    .Y(n_706));
 INVxp33_ASAP7_75t_R g44670 (.A(exp_r[3]),
    .Y(n_43));
 INVxp33_ASAP7_75t_R g44671 (.A(exp_r[0]),
    .Y(n_3819));
 INVxp33_ASAP7_75t_R g44674 (.A(n_13972),
    .Y(n_702));
 INVxp33_ASAP7_75t_R g44676 (.A(exp_r[5]),
    .Y(n_700));
 AO222x2_ASAP7_75t_R g44844 (.A1(n_680),
    .A2(fract_i2f[18]),
    .B1(n_677),
    .B2(quo[20]),
    .C1(n_674),
    .C2(prod[18]),
    .Y(n_650));
 AO222x2_ASAP7_75t_R g44845 (.A1(n_679),
    .A2(fract_i2f[19]),
    .B1(n_676),
    .B2(quo[21]),
    .C1(n_674),
    .C2(prod[19]),
    .Y(n_649));
 OR3x1_ASAP7_75t_R g44846 (.A(n_925),
    .B(fpu_op_r3[2]),
    .C(fpu_op_r3[0]),
    .Y(n_3850));
 OR2x2_ASAP7_75t_R g44847 (.A(fpu_op_r3[1]),
    .B(fpu_op_r3[2]),
    .Y(n_3498));
 XOR2xp5_ASAP7_75t_R g44848 (.A(n_1158),
    .B(opa_r1[16]),
    .Y(n_648));
 XOR2xp5_ASAP7_75t_R g44849 (.A(n_1148),
    .B(opa_r1[14]),
    .Y(n_647));
 XOR2xp5_ASAP7_75t_R g44850 (.A(n_1147),
    .B(n_1049),
    .Y(n_646));
 XOR2xp5_ASAP7_75t_R g44851 (.A(n_1142),
    .B(opa_r1[12]),
    .Y(n_645));
 XOR2xp5_ASAP7_75t_R g44852 (.A(n_1132),
    .B(opa_r1[10]),
    .Y(n_644));
 XOR2xp5_ASAP7_75t_R g44853 (.A(n_1081),
    .B(opa_r1[8]),
    .Y(n_643));
 XOR2xp5_ASAP7_75t_R g44854 (.A(n_1061),
    .B(opa_r1[6]),
    .Y(n_642));
 XOR2xp5_ASAP7_75t_R g44856 (.A(n_1023),
    .B(opa_r1[4]),
    .Y(n_640));
 NAND2xp33_ASAP7_75t_R g52051__1705 (.A(n_3555),
    .B(n_2875),
    .Y(u4_n_1454));
 INVxp33_ASAP7_75t_R g52052 (.A(u4_n_1442),
    .Y(n_2875));
 NAND2xp33_ASAP7_75t_R g52053__5122 (.A(n_2874),
    .B(n_3558),
    .Y(u4_n_1442));
 INVxp33_ASAP7_75t_R g52054 (.A(n_2874),
    .Y(n_3559));
 AOI22xp33_ASAP7_75t_R g52055__8246 (.A1(n_2455),
    .A2(n_2873),
    .B1(n_2456),
    .B2(u4_n_1248),
    .Y(n_2874));
 OR5x1_ASAP7_75t_R g52056__7098 (.A(n_2871),
    .B(n_2870),
    .C(u4_fract_trunc[16]),
    .D(u4_fract_trunc[18]),
    .E(u4_fract_trunc[17]),
    .Y(n_2873));
 NAND5xp2_ASAP7_75t_R g52057__6131 (.A(n_2872),
    .B(n_2860),
    .C(n_2849),
    .D(n_2850),
    .E(n_2855),
    .Y(u4_n_1248));
 NOR4xp25_ASAP7_75t_R g52058__1881 (.A(n_2870),
    .B(n_2835),
    .C(n_2065),
    .D(n_2171),
    .Y(n_2872));
 AO21x1_ASAP7_75t_R g52059__5115 (.A1(n_1844),
    .A2(u4_fract_trunc[24]),
    .B(n_2869),
    .Y(n_2871));
 OAI221xp5_ASAP7_75t_R g52060__7482 (.A1(n_2660),
    .A2(n_2563),
    .B1(n_2547),
    .B2(n_2324),
    .C(n_2868),
    .Y(n_2870));
 OR3x1_ASAP7_75t_R g52061__4733 (.A(n_2866),
    .B(u4_fract_trunc[20]),
    .C(u4_fract_trunc[21]),
    .Y(n_2869));
 AOI211xp5_ASAP7_75t_R g52062__6161 (.A1(n_2556),
    .A2(n_2092),
    .B(n_2867),
    .C(n_2510),
    .Y(n_2868));
 NAND5xp2_ASAP7_75t_R g52063__9315 (.A(n_2864),
    .B(n_2856),
    .C(n_2781),
    .D(n_2792),
    .E(n_2542),
    .Y(n_2867));
 NAND3xp33_ASAP7_75t_R g52064__9945 (.A(n_2860),
    .B(n_2859),
    .C(n_2865),
    .Y(n_2866));
 NAND5xp2_ASAP7_75t_R g52065__2883 (.A(n_2863),
    .B(u4_fract_out[6]),
    .C(u4_fract_out[5]),
    .D(u4_fract_out[4]),
    .E(u4_g),
    .Y(u4_n_1439));
 NOR5xp2_ASAP7_75t_R g52066__2346 (.A(n_2861),
    .B(u4_fract_trunc[15]),
    .C(u4_fract_trunc[14]),
    .D(u4_fract_trunc[19]),
    .E(n_2835),
    .Y(n_2865));
 AOI211xp5_ASAP7_75t_R g52067__1666 (.A1(n_2556),
    .A2(fract_denorm[8]),
    .B(n_2862),
    .C(n_2540),
    .Y(n_2864));
 AND5x1_ASAP7_75t_R g52068__7410 (.A(u4_fract_out[3]),
    .B(u4_fract_out[2]),
    .C(u4_fract_out[1]),
    .D(n_2064),
    .E(n_2168),
    .Y(n_2863));
 OAI221xp5_ASAP7_75t_R g52069__6417 (.A1(n_2661),
    .A2(n_2563),
    .B1(n_2553),
    .B2(n_2365),
    .C(n_2857),
    .Y(n_2862));
 NAND4xp25_ASAP7_75t_R g52070__5477 (.A(n_2848),
    .B(n_2855),
    .C(n_2849),
    .D(n_2850),
    .Y(n_2861));
 OAI221xp5_ASAP7_75t_R g52071__2398 (.A1(n_2555),
    .A2(n_2313),
    .B1(n_2547),
    .B2(n_2303),
    .C(n_2858),
    .Y(u4_fract_trunc[15]));
 OAI211xp5_ASAP7_75t_R g52072__5107 (.A1(n_2565),
    .A2(n_2682),
    .B(n_2838),
    .C(n_2791),
    .Y(u4_fract_out[15]));
 OAI211xp5_ASAP7_75t_R g52073__6260 (.A1(n_2565),
    .A2(n_2683),
    .B(n_2843),
    .C(n_2784),
    .Y(u4_fract_out[16]));
 AO221x1_ASAP7_75t_R g52074__4319 (.A1(n_2687),
    .A2(n_2564),
    .B1(n_2793),
    .B2(n_2524),
    .C(n_2851),
    .Y(u4_fract_out[21]));
 AOI221xp5_ASAP7_75t_R g52075__8428 (.A1(n_2503),
    .A2(n_2416),
    .B1(n_2556),
    .B2(n_2317),
    .C(n_2853),
    .Y(n_2860));
 OAI221xp5_ASAP7_75t_R g52076__5526 (.A1(n_2553),
    .A2(n_2324),
    .B1(n_2533),
    .B2(n_2295),
    .C(n_2852),
    .Y(u4_fract_trunc[14]));
 INVxp33_ASAP7_75t_R g52077 (.A(n_2859),
    .Y(u4_fract_trunc[13]));
 AOI221xp5_ASAP7_75t_R g52078__6783 (.A1(n_2549),
    .A2(n_2341),
    .B1(n_2503),
    .B2(n_2436),
    .C(n_2836),
    .Y(n_2858));
 AOI211xp5_ASAP7_75t_R g52079__3680 (.A1(n_1835),
    .A2(n_2441),
    .B(n_2840),
    .C(n_2658),
    .Y(n_2857));
 AOI211xp5_ASAP7_75t_R g52080__1617 (.A1(n_2556),
    .A2(n_2353),
    .B(n_2846),
    .C(n_2601),
    .Y(n_2856));
 OAI321xp33_ASAP7_75t_R g52081__2802 (.A1(n_2686),
    .A2(n_2560),
    .A3(n_2501),
    .B1(n_2552),
    .B2(n_2796),
    .C(n_2847),
    .Y(u4_fract_out[19]));
 OAI321xp33_ASAP7_75t_R g52082__1705 (.A1(n_2719),
    .A2(n_2560),
    .A3(n_2501),
    .B1(n_2526),
    .B2(n_2787),
    .C(n_2841),
    .Y(u4_fract_out[20]));
 AOI221xp5_ASAP7_75t_R g52083__5122 (.A1(n_2556),
    .A2(n_2335),
    .B1(n_2549),
    .B2(n_2318),
    .C(n_2854),
    .Y(n_2859));
 OAI21xp33_ASAP7_75t_R g52084__8246 (.A1(n_2300),
    .A2(n_2536),
    .B(n_2839),
    .Y(n_2854));
 OAI221xp5_ASAP7_75t_R g52085__7098 (.A1(n_2685),
    .A2(n_2565),
    .B1(n_2808),
    .B2(n_2526),
    .C(n_2842),
    .Y(u4_fract_out[22]));
 OAI211xp5_ASAP7_75t_R g52086__6131 (.A1(n_2526),
    .A2(n_2810),
    .B(n_2803),
    .C(n_2813),
    .Y(u4_fract_out[17]));
 OAI221xp5_ASAP7_75t_R g52087__1881 (.A1(n_2809),
    .A2(n_2525),
    .B1(n_2766),
    .B2(n_2526),
    .C(n_2575),
    .Y(u4_fract_out[2]));
 AOI221xp5_ASAP7_75t_R g52088__5115 (.A1(n_2503),
    .A2(n_2410),
    .B1(n_2532),
    .B2(n_2390),
    .C(n_2845),
    .Y(n_2855));
 OAI31xp33_ASAP7_75t_R g52089__7482 (.A1(n_2483),
    .A2(fract_denorm[35]),
    .A3(fract_denorm[36]),
    .B(u4_fract_trunc[24]),
    .Y(n_3558));
 OAI221xp5_ASAP7_75t_R g52090__4733 (.A1(n_2550),
    .A2(n_2305),
    .B1(n_2536),
    .B2(n_2301),
    .C(n_2833),
    .Y(n_2853));
 AOI211xp5_ASAP7_75t_R g52091__6161 (.A1(n_2503),
    .A2(n_2435),
    .B(n_2823),
    .C(n_2602),
    .Y(n_2852));
 OAI221xp5_ASAP7_75t_R g52092__9315 (.A1(n_2685),
    .A2(n_2563),
    .B1(n_2766),
    .B2(n_2552),
    .C(n_2844),
    .Y(u4_fract_out[18]));
 OAI222xp33_ASAP7_75t_R g52093__9945 (.A1(n_2799),
    .A2(n_2552),
    .B1(n_2807),
    .B2(n_2526),
    .C1(n_2567),
    .C2(n_2295),
    .Y(n_2851));
 OAI221xp5_ASAP7_75t_R g52094__2883 (.A1(n_2517),
    .A2(n_2412),
    .B1(n_2535),
    .B2(n_2392),
    .C(n_2837),
    .Y(u4_fract_out[1]));
 OAI221xp5_ASAP7_75t_R g52095__2346 (.A1(n_2807),
    .A2(n_2525),
    .B1(n_2799),
    .B2(n_2526),
    .C(n_2579),
    .Y(u4_fract_out[5]));
 OAI221xp5_ASAP7_75t_R g52096__1666 (.A1(n_2808),
    .A2(n_2525),
    .B1(n_2797),
    .B2(n_2526),
    .C(n_2574),
    .Y(u4_fract_out[6]));
 OAI221xp5_ASAP7_75t_R g52097__7410 (.A1(n_2758),
    .A2(n_2597),
    .B1(n_2517),
    .B2(n_2404),
    .C(n_2825),
    .Y(u4_fract_out[12]));
 NOR2xp33_ASAP7_75t_R g52098__6417 (.A(u4_fract_trunc[22]),
    .B(u4_fract_trunc[23]),
    .Y(n_2848));
 OAI221xp5_ASAP7_75t_R g52099__5477 (.A1(n_2726),
    .A2(n_1830),
    .B1(n_2661),
    .B2(n_2598),
    .C(n_2828),
    .Y(u4_fract_out[9]));
 AOI221xp5_ASAP7_75t_R g52100__2398 (.A1(n_2733),
    .A2(n_2544),
    .B1(n_2789),
    .B2(n_2527),
    .C(n_2742),
    .Y(n_2847));
 OAI221xp5_ASAP7_75t_R g52101__5107 (.A1(n_2737),
    .A2(n_2560),
    .B1(n_2517),
    .B2(n_2409),
    .C(n_2830),
    .Y(u4_fract_out[7]));
 OAI221xp5_ASAP7_75t_R g52102__6260 (.A1(n_2502),
    .A2(n_2414),
    .B1(n_2555),
    .B2(n_2355),
    .C(n_2826),
    .Y(n_2846));
 OAI221xp5_ASAP7_75t_R g52103__4319 (.A1(n_2740),
    .A2(n_2543),
    .B1(n_2655),
    .B2(n_2597),
    .C(n_2827),
    .Y(u4_fract_out[8]));
 AOI221xp5_ASAP7_75t_R g52104__8428 (.A1(n_2532),
    .A2(n_2393),
    .B1(n_1835),
    .B2(n_2386),
    .C(n_2829),
    .Y(n_2850));
 OAI221xp5_ASAP7_75t_R g52105__5526 (.A1(n_2765),
    .A2(n_2526),
    .B1(n_2785),
    .B2(n_2525),
    .C(n_2577),
    .Y(u4_g));
 AOI211xp5_ASAP7_75t_R g52106__6783 (.A1(n_1835),
    .A2(n_2387),
    .B(n_2834),
    .C(n_2585),
    .Y(n_2849));
 OAI221xp5_ASAP7_75t_R g52107__3680 (.A1(n_2516),
    .A2(n_2422),
    .B1(n_2535),
    .B2(n_2391),
    .C(n_2832),
    .Y(u4_fract_trunc[24]));
 OAI221xp5_ASAP7_75t_R g52108__1617 (.A1(n_2550),
    .A2(n_2308),
    .B1(n_2555),
    .B2(n_2311),
    .C(n_2801),
    .Y(n_2845));
 OA21x2_ASAP7_75t_R g52109__2802 (.A1(n_2526),
    .A2(n_2809),
    .B(n_2816),
    .Y(n_2844));
 OA222x2_ASAP7_75t_R g52110__1705 (.A1(n_2719),
    .A2(n_2563),
    .B1(n_2765),
    .B2(n_2552),
    .C1(n_2785),
    .C2(n_2526),
    .Y(n_2843));
 AOI221xp5_ASAP7_75t_R g52111__5122 (.A1(n_2795),
    .A2(n_2524),
    .B1(n_2554),
    .B2(n_2253),
    .C(n_2822),
    .Y(n_2842));
 AOI221xp5_ASAP7_75t_R g52112__8246 (.A1(n_2738),
    .A2(n_2544),
    .B1(n_2798),
    .B2(n_2551),
    .C(n_2750),
    .Y(n_2841));
 OR3x1_ASAP7_75t_R g52113__7098 (.A(n_2821),
    .B(n_2604),
    .C(n_2512),
    .Y(n_2840));
 AOI221xp5_ASAP7_75t_R g52114__6131 (.A1(n_2798),
    .A2(n_2524),
    .B1(n_2548),
    .B2(n_2309),
    .C(n_2606),
    .Y(n_2839));
 AOI221xp5_ASAP7_75t_R g52115__1881 (.A1(n_2767),
    .A2(n_2551),
    .B1(n_2786),
    .B2(n_2527),
    .C(n_2721),
    .Y(n_2838));
 AOI22xp33_ASAP7_75t_R g52116__5115 (.A1(n_2527),
    .A2(n_2768),
    .B1(n_2524),
    .B2(n_2811),
    .Y(n_2837));
 OAI222xp33_ASAP7_75t_R g52117__7482 (.A1(n_2536),
    .A2(n_2254),
    .B1(n_2797),
    .B2(n_2525),
    .C1(n_2553),
    .C2(n_2342),
    .Y(n_2836));
 OAI221xp5_ASAP7_75t_R g52118__4733 (.A1(n_2790),
    .A2(n_2525),
    .B1(n_2796),
    .B2(n_2526),
    .C(n_2578),
    .Y(u4_fract_out[3]));
 OAI221xp5_ASAP7_75t_R g52119__6161 (.A1(n_2517),
    .A2(n_2434),
    .B1(n_2538),
    .B2(n_2300),
    .C(n_2824),
    .Y(u4_fract_out[4]));
 OAI221xp5_ASAP7_75t_R g52120__9315 (.A1(n_2778),
    .A2(n_2526),
    .B1(n_2517),
    .B2(n_2428),
    .C(n_2800),
    .Y(u4_fract_out[10]));
 OAI221xp5_ASAP7_75t_R g52121__9945 (.A1(n_2739),
    .A2(n_2543),
    .B1(n_2517),
    .B2(n_2399),
    .C(n_2819),
    .Y(u4_fract_out[11]));
 OAI221xp5_ASAP7_75t_R g52122__2883 (.A1(n_2757),
    .A2(n_2597),
    .B1(n_2771),
    .B2(n_2526),
    .C(n_2818),
    .Y(u4_fract_out[14]));
 OAI221xp5_ASAP7_75t_R g52123__2346 (.A1(n_2769),
    .A2(n_2526),
    .B1(n_2516),
    .B2(n_2401),
    .C(n_2820),
    .Y(u4_fract_out[13]));
 OAI221xp5_ASAP7_75t_R g52124__1666 (.A1(n_2766),
    .A2(n_2525),
    .B1(n_2502),
    .B2(n_2432),
    .C(n_2603),
    .Y(n_2834));
 OAI221xp5_ASAP7_75t_R g52125__7410 (.A1(n_2780),
    .A2(n_2525),
    .B1(n_2610),
    .B2(n_2570),
    .C(n_2571),
    .Y(u4_fract_trunc[16]));
 OAI221xp5_ASAP7_75t_R g52126__6417 (.A1(n_2533),
    .A2(n_2391),
    .B1(n_2550),
    .B2(n_2315),
    .C(n_2817),
    .Y(n_2835));
 OAI221xp5_ASAP7_75t_R g52127__5477 (.A1(n_2516),
    .A2(n_2417),
    .B1(n_2502),
    .B2(n_2431),
    .C(n_2804),
    .Y(u4_fract_trunc[17]));
 OAI221xp5_ASAP7_75t_R g52128__2398 (.A1(n_2757),
    .A2(n_2568),
    .B1(n_2771),
    .B2(n_2525),
    .C(n_2572),
    .Y(u4_fract_trunc[23]));
 OAI221xp5_ASAP7_75t_R g52129__5107 (.A1(n_2516),
    .A2(n_2421),
    .B1(n_2502),
    .B2(n_2428),
    .C(n_2812),
    .Y(u4_fract_trunc[19]));
 OAI221xp5_ASAP7_75t_R g52130__6260 (.A1(n_2516),
    .A2(n_2413),
    .B1(n_2502),
    .B2(n_2401),
    .C(n_2815),
    .Y(u4_fract_trunc[22]));
 OAI221xp5_ASAP7_75t_R g52131__4319 (.A1(n_2516),
    .A2(n_2418),
    .B1(n_2502),
    .B2(n_2399),
    .C(n_2814),
    .Y(u4_fract_trunc[20]));
 INVxp33_ASAP7_75t_R g52132 (.A(n_2831),
    .Y(n_2833));
 AOI22xp33_ASAP7_75t_R g52133__8428 (.A1(n_2527),
    .A2(n_2767),
    .B1(n_2524),
    .B2(n_2786),
    .Y(n_2832));
 OAI22xp33_ASAP7_75t_R g52134__5526 (.A1(n_2525),
    .A2(n_2796),
    .B1(n_2315),
    .B2(n_2547),
    .Y(n_2831));
 AOI21xp33_ASAP7_75t_R g52135__6783 (.A1(n_2741),
    .A2(n_2544),
    .B(n_2802),
    .Y(n_2830));
 OAI221xp5_ASAP7_75t_R g52136__3680 (.A1(n_2547),
    .A2(n_2302),
    .B1(n_2550),
    .B2(n_2336),
    .C(n_2805),
    .Y(n_2829));
 AOI222xp33_ASAP7_75t_R g52137__1617 (.A1(n_2736),
    .A2(n_1830),
    .B1(n_2774),
    .B2(n_2527),
    .C1(n_1834),
    .C2(n_2430),
    .Y(n_2828));
 AOI221xp5_ASAP7_75t_R g52138__2802 (.A1(n_2779),
    .A2(n_2527),
    .B1(n_2732),
    .B2(n_2561),
    .C(n_2558),
    .Y(n_2827));
 AOI221xp5_ASAP7_75t_R g52139__1705 (.A1(n_2505),
    .A2(n_2405),
    .B1(n_2548),
    .B2(n_2312),
    .C(n_2782),
    .Y(n_2826));
 AOI222xp33_ASAP7_75t_R g52140__5122 (.A1(n_2738),
    .A2(n_2561),
    .B1(n_2735),
    .B2(n_2544),
    .C1(n_2775),
    .C2(n_2527),
    .Y(n_2825));
 AOI22xp33_ASAP7_75t_R g52141__8246 (.A1(n_2524),
    .A2(n_2788),
    .B1(n_2527),
    .B2(n_2798),
    .Y(n_2824));
 OAI22xp33_ASAP7_75t_R g52142__7098 (.A1(n_2525),
    .A2(n_2799),
    .B1(n_2319),
    .B2(n_2550),
    .Y(n_2823));
 OAI221xp5_ASAP7_75t_R g52143__6131 (.A1(n_2773),
    .A2(n_2525),
    .B1(n_2661),
    .B2(n_2570),
    .C(n_2573),
    .Y(u4_fract_trunc[18]));
 OAI221xp5_ASAP7_75t_R g52144__1881 (.A1(n_2758),
    .A2(n_2568),
    .B1(n_2776),
    .B2(n_2525),
    .C(n_2576),
    .Y(u4_fract_trunc[21]));
 NOR2xp33_ASAP7_75t_R g52145__5115 (.A(n_2552),
    .B(n_2797),
    .Y(n_2822));
 A2O1A1Ixp33_ASAP7_75t_R g52146__7482 (.A1(n_2399),
    .A2(n_2431),
    .B(n_2504),
    .C(n_2794),
    .Y(n_2821));
 AOI222xp33_ASAP7_75t_R g52147__4733 (.A1(n_2736),
    .A2(n_1829),
    .B1(n_2724),
    .B2(n_2501),
    .C1(n_2760),
    .C2(n_2596),
    .Y(n_2820));
 AOI222xp33_ASAP7_75t_R g52148__6161 (.A1(n_2733),
    .A2(n_2561),
    .B1(n_2759),
    .B2(n_2596),
    .C1(n_2777),
    .C2(n_2527),
    .Y(n_2819));
 AOI222xp33_ASAP7_75t_R g52149__9315 (.A1(n_2734),
    .A2(n_1829),
    .B1(n_2725),
    .B2(n_2501),
    .C1(n_1835),
    .C2(n_2402),
    .Y(n_2818));
 AOI221xp5_ASAP7_75t_R g52150__9945 (.A1(n_2767),
    .A2(n_2524),
    .B1(n_2548),
    .B2(n_2317),
    .C(n_2514),
    .Y(n_2817));
 AOI222xp33_ASAP7_75t_R g52151__2883 (.A1(n_2730),
    .A2(n_2544),
    .B1(n_2679),
    .B2(n_2564),
    .C1(n_2566),
    .C2(n_2389),
    .Y(n_2816));
 AOI22xp33_ASAP7_75t_R g52152__2346 (.A1(n_2569),
    .A2(n_2760),
    .B1(n_2524),
    .B2(n_2770),
    .Y(n_2815));
 AOI22xp33_ASAP7_75t_R g52153__1666 (.A1(n_2569),
    .A2(n_2759),
    .B1(n_2524),
    .B2(n_2777),
    .Y(n_2814));
 AOI22xp33_ASAP7_75t_R g52154__7410 (.A1(n_2551),
    .A2(n_2768),
    .B1(n_2562),
    .B2(n_2687),
    .Y(n_2813));
 INVxp33_ASAP7_75t_R g52155 (.A(n_2806),
    .Y(n_2812));
 INVxp33_ASAP7_75t_R g52156 (.A(n_2810),
    .Y(n_2811));
 OAI22xp33_ASAP7_75t_R g52157__6417 (.A1(n_2525),
    .A2(n_2778),
    .B1(n_2570),
    .B2(n_2660),
    .Y(n_2806));
 AOI22xp33_ASAP7_75t_R g52158__5477 (.A1(n_2524),
    .A2(n_2768),
    .B1(n_2411),
    .B2(n_2503),
    .Y(n_2805));
 AOI22xp33_ASAP7_75t_R g52159__2398 (.A1(n_2524),
    .A2(n_2779),
    .B1(n_2569),
    .B2(n_2654),
    .Y(n_2804));
 AOI222xp33_ASAP7_75t_R g52160__5107 (.A1(n_2727),
    .A2(n_2544),
    .B1(n_2566),
    .B2(n_2393),
    .C1(n_2681),
    .C2(n_2564),
    .Y(n_2803));
 OAI22xp33_ASAP7_75t_R g52161__6260 (.A1(n_2526),
    .A2(n_2780),
    .B1(n_2598),
    .B2(n_2610),
    .Y(n_2802));
 AOI22xp33_ASAP7_75t_R g52162__4319 (.A1(n_2524),
    .A2(n_2764),
    .B1(n_2335),
    .B2(n_2548),
    .Y(n_2801));
 AOI221xp5_ASAP7_75t_R g52163__8428 (.A1(n_2731),
    .A2(n_1831),
    .B1(n_2734),
    .B2(n_1830),
    .C(n_2723),
    .Y(n_2800));
 AOI222xp33_ASAP7_75t_R g52164__5526 (.A1(n_2673),
    .A2(n_2521),
    .B1(n_2744),
    .B2(n_2493),
    .C1(n_2663),
    .C2(n_2519),
    .Y(n_2810));
 AOI222xp33_ASAP7_75t_R g52165__6783 (.A1(n_2747),
    .A2(n_2493),
    .B1(n_2696),
    .B2(n_2521),
    .C1(n_2695),
    .C2(n_2519),
    .Y(n_2809));
 AOI222xp33_ASAP7_75t_R g52166__3680 (.A1(n_2748),
    .A2(n_2493),
    .B1(n_2695),
    .B2(n_2521),
    .C1(n_2671),
    .C2(n_2519),
    .Y(n_2808));
 AOI222xp33_ASAP7_75t_R g52167__1617 (.A1(n_2746),
    .A2(n_2493),
    .B1(n_2663),
    .B2(n_2521),
    .C1(n_2665),
    .C2(n_2519),
    .Y(n_2807));
 A2O1A1Ixp33_ASAP7_75t_R g52168__2802 (.A1(n_2634),
    .A2(n_2648),
    .B(n_2529),
    .C(n_2762),
    .Y(n_2795));
 OAI21xp33_ASAP7_75t_R g52169__1705 (.A1(n_2654),
    .A2(n_2759),
    .B(n_2561),
    .Y(n_2794));
 A2O1A1Ixp33_ASAP7_75t_R g52170__5122 (.A1(n_2626),
    .A2(n_2647),
    .B(n_2529),
    .C(n_2763),
    .Y(n_2793));
 AOI22xp33_ASAP7_75t_R g52171__8246 (.A1(n_2561),
    .A2(n_2760),
    .B1(n_2400),
    .B2(n_2505),
    .Y(n_2792));
 AOI222xp33_ASAP7_75t_R g52172__7098 (.A1(n_2673),
    .A2(n_2528),
    .B1(n_2697),
    .B2(n_2530),
    .C1(n_2760),
    .C2(n_2494),
    .Y(n_2799));
 OAI222xp33_ASAP7_75t_R g52173__6131 (.A1(n_2689),
    .A2(n_2529),
    .B1(n_2758),
    .B2(n_2493),
    .C1(n_2691),
    .C2(n_2531),
    .Y(n_2798));
 AOI221xp5_ASAP7_75t_R g52174__1881 (.A1(n_2696),
    .A2(n_2528),
    .B1(n_2698),
    .B2(n_2530),
    .C(n_2772),
    .Y(n_2797));
 AOI21xp33_ASAP7_75t_R g52175__5115 (.A1(n_2759),
    .A2(n_2494),
    .B(n_2753),
    .Y(n_2796));
 INVxp33_ASAP7_75t_R g52176 (.A(n_2783),
    .Y(n_2791));
 INVxp33_ASAP7_75t_R g52177 (.A(n_2789),
    .Y(n_2790));
 INVxp33_ASAP7_75t_R g52178 (.A(n_2787),
    .Y(n_2788));
 AOI22xp33_ASAP7_75t_R g52179__7482 (.A1(n_2544),
    .A2(n_2732),
    .B1(n_2390),
    .B2(n_2566),
    .Y(n_2784));
 OAI22xp33_ASAP7_75t_R g52180__4733 (.A1(n_2737),
    .A2(n_2543),
    .B1(n_2567),
    .B2(n_2391),
    .Y(n_2783));
 OAI221xp5_ASAP7_75t_R g52181__6161 (.A1(n_2758),
    .A2(n_2560),
    .B1(n_2553),
    .B2(n_2091),
    .C(n_2584),
    .Y(n_2782));
 AOI22xp33_ASAP7_75t_R g52182__9315 (.A1(n_2561),
    .A2(n_2756),
    .B1(fract_denorm[8]),
    .B2(n_2554),
    .Y(n_2781));
 OAI222xp33_ASAP7_75t_R g52183__9945 (.A1(n_2705),
    .A2(n_2518),
    .B1(n_2739),
    .B2(n_2494),
    .C1(n_2700),
    .C2(n_2520),
    .Y(n_2789));
 AOI222xp33_ASAP7_75t_R g52184__2883 (.A1(n_2703),
    .A2(n_2519),
    .B1(n_2666),
    .B2(n_2521),
    .C1(n_2735),
    .C2(n_2493),
    .Y(n_2787));
 AO21x1_ASAP7_75t_R g52185__2346 (.A1(n_2493),
    .A2(n_2741),
    .B(n_2755),
    .Y(n_2786));
 OA222x2_ASAP7_75t_R g52186__1666 (.A1(n_2740),
    .A2(n_2494),
    .B1(n_2667),
    .B2(n_2518),
    .C1(n_2689),
    .C2(n_2520),
    .Y(n_2785));
 INVxp33_ASAP7_75t_R g52187 (.A(n_2775),
    .Y(n_2776));
 INVxp33_ASAP7_75t_R g52188 (.A(n_2773),
    .Y(n_2774));
 NOR2xp33_ASAP7_75t_R g52189__7410 (.A(n_2493),
    .B(n_2757),
    .Y(n_2772));
 AOI221xp5_ASAP7_75t_R g52190__6417 (.A1(n_2701),
    .A2(n_2519),
    .B1(n_2692),
    .B2(n_2530),
    .C(n_2754),
    .Y(n_2780));
 OAI221xp5_ASAP7_75t_R g52191__5477 (.A1(n_2667),
    .A2(n_2529),
    .B1(n_2707),
    .B2(n_2520),
    .C(n_2761),
    .Y(n_2779));
 AOI221xp5_ASAP7_75t_R g52192__2398 (.A1(n_2698),
    .A2(n_2519),
    .B1(n_2696),
    .B2(n_2530),
    .C(n_2752),
    .Y(n_2778));
 OAI221xp5_ASAP7_75t_R g52193__5107 (.A1(n_2705),
    .A2(n_2529),
    .B1(n_2702),
    .B2(n_2520),
    .C(n_2743),
    .Y(n_2777));
 OAI221xp5_ASAP7_75t_R g52194__6260 (.A1(n_2689),
    .A2(n_2518),
    .B1(n_2667),
    .B2(n_2531),
    .C(n_2745),
    .Y(n_2775));
 AOI221xp5_ASAP7_75t_R g52195__4319 (.A1(n_2697),
    .A2(n_2519),
    .B1(n_2673),
    .B2(n_2530),
    .C(n_2751),
    .Y(n_2773));
 INVxp33_ASAP7_75t_R g52196 (.A(n_2769),
    .Y(n_2770));
 INVxp33_ASAP7_75t_R g52197 (.A(n_2764),
    .Y(n_2765));
 OAI221xp5_ASAP7_75t_R g52198__8428 (.A1(n_2681),
    .A2(n_1829),
    .B1(n_2708),
    .B2(n_2501),
    .C(n_2494),
    .Y(n_2763));
 OAI221xp5_ASAP7_75t_R g52199__5526 (.A1(n_2679),
    .A2(n_1829),
    .B1(n_2674),
    .B2(n_2501),
    .C(n_2494),
    .Y(n_2762));
 AOI221xp5_ASAP7_75t_R g52200__6783 (.A1(n_2671),
    .A2(n_2528),
    .B1(n_2698),
    .B2(n_2521),
    .C(n_2729),
    .Y(n_2771));
 AOI221xp5_ASAP7_75t_R g52201__3680 (.A1(n_2665),
    .A2(n_2528),
    .B1(n_2697),
    .B2(n_2521),
    .C(n_2728),
    .Y(n_2769));
 OAI221xp5_ASAP7_75t_R g52202__1617 (.A1(n_2661),
    .A2(n_2518),
    .B1(n_2710),
    .B2(n_2531),
    .C(n_2722),
    .Y(n_2768));
 OAI222xp33_ASAP7_75t_R g52203__2802 (.A1(n_2702),
    .A2(n_2529),
    .B1(n_2676),
    .B2(n_2531),
    .C1(n_2610),
    .C2(n_2518),
    .Y(n_2767));
 AOI221xp5_ASAP7_75t_R g52204__1705 (.A1(n_2698),
    .A2(n_2528),
    .B1(n_2704),
    .B2(n_2530),
    .C(n_2720),
    .Y(n_2766));
 OAI222xp33_ASAP7_75t_R g52205__5122 (.A1(n_2707),
    .A2(n_2531),
    .B1(n_2691),
    .B2(n_2529),
    .C1(n_2655),
    .C2(n_2493),
    .Y(n_2764));
 INVxp33_ASAP7_75t_R g52206 (.A(n_2749),
    .Y(n_2761));
 INVxp33_ASAP7_75t_R g52207 (.A(n_2757),
    .Y(n_2756));
 OAI22xp33_ASAP7_75t_R g52208__8246 (.A1(n_2518),
    .A2(n_2700),
    .B1(n_2520),
    .B2(n_2693),
    .Y(n_2755));
 OAI22xp33_ASAP7_75t_R g52209__7098 (.A1(n_2529),
    .A2(n_2700),
    .B1(n_2520),
    .B2(n_2676),
    .Y(n_2754));
 OAI22xp33_ASAP7_75t_R g52210__6131 (.A1(n_2529),
    .A2(n_2693),
    .B1(n_2531),
    .B2(n_2702),
    .Y(n_2753));
 AO22x1_ASAP7_75t_R g52211__1881 (.A1(n_2528),
    .A2(n_2695),
    .B1(n_2521),
    .B2(n_2704),
    .Y(n_2752));
 OAI22xp33_ASAP7_75t_R g52212__5115 (.A1(n_2529),
    .A2(n_2662),
    .B1(n_2520),
    .B2(n_2710),
    .Y(n_2751));
 OAI22xp33_ASAP7_75t_R g52213__7482 (.A1(n_2657),
    .A2(n_2563),
    .B1(n_2553),
    .B2(n_2300),
    .Y(n_2750));
 OAI22xp33_ASAP7_75t_R g52214__4733 (.A1(n_2518),
    .A2(n_2691),
    .B1(n_2531),
    .B2(n_2689),
    .Y(n_2749));
 OAI22xp33_ASAP7_75t_R g52215__6161 (.A1(n_1831),
    .A2(n_2694),
    .B1(n_1830),
    .B2(n_2711),
    .Y(n_2748));
 OAI22xp33_ASAP7_75t_R g52216__9315 (.A1(n_2711),
    .A2(n_1833),
    .B1(n_2670),
    .B2(n_1830),
    .Y(n_2747));
 OAI22xp33_ASAP7_75t_R g52217__9945 (.A1(n_1831),
    .A2(n_2669),
    .B1(n_1830),
    .B2(n_2677),
    .Y(n_2746));
 AOI22xp33_ASAP7_75t_R g52218__2883 (.A1(n_2528),
    .A2(n_2703),
    .B1(n_2521),
    .B2(n_2690),
    .Y(n_2745));
 OAI22xp33_ASAP7_75t_R g52219__2346 (.A1(n_1832),
    .A2(n_2664),
    .B1(n_1833),
    .B2(n_2677),
    .Y(n_2744));
 AOI22xp33_ASAP7_75t_R g52220__1666 (.A1(n_2519),
    .A2(n_2692),
    .B1(n_2530),
    .B2(n_2699),
    .Y(n_2743));
 OAI22xp33_ASAP7_75t_R g52221__7410 (.A1(n_2563),
    .A2(n_2656),
    .B1(n_2301),
    .B2(n_2553),
    .Y(n_2742));
 OAI22xp33_ASAP7_75t_R g52222__6417 (.A1(n_1833),
    .A2(n_2710),
    .B1(n_1832),
    .B2(n_2661),
    .Y(n_2760));
 OAI22xp33_ASAP7_75t_R g52223__5477 (.A1(n_1831),
    .A2(n_2676),
    .B1(n_1832),
    .B2(n_2610),
    .Y(n_2759));
 AOI22xp33_ASAP7_75t_R g52224__2398 (.A1(n_1832),
    .A2(n_2706),
    .B1(n_1833),
    .B2(n_2611),
    .Y(n_2758));
 AOI22xp33_ASAP7_75t_R g52225__5107 (.A1(n_1830),
    .A2(n_2704),
    .B1(n_1833),
    .B2(n_2659),
    .Y(n_2757));
 OAI22xp33_ASAP7_75t_R g52226__6260 (.A1(n_2560),
    .A2(n_2694),
    .B1(n_2543),
    .B2(n_2670),
    .Y(n_2731));
 OAI22xp33_ASAP7_75t_R g52227__4319 (.A1(n_1829),
    .A2(n_2675),
    .B1(n_2501),
    .B2(n_2694),
    .Y(n_2730));
 AO22x1_ASAP7_75t_R g52228__8428 (.A1(n_2519),
    .A2(n_2696),
    .B1(n_2530),
    .B2(n_2695),
    .Y(n_2729));
 OAI22xp33_ASAP7_75t_R g52229__5526 (.A1(n_2518),
    .A2(n_2672),
    .B1(n_2531),
    .B2(n_2662),
    .Y(n_2728));
 OAI22xp33_ASAP7_75t_R g52230__6783 (.A1(n_1829),
    .A2(n_2709),
    .B1(n_2501),
    .B2(n_2669),
    .Y(n_2727));
 AOI22xp33_ASAP7_75t_R g52231__3680 (.A1(n_2668),
    .A2(n_2561),
    .B1(n_2544),
    .B2(n_2665),
    .Y(n_2726));
 OAI22xp33_ASAP7_75t_R g52232__1617 (.A1(n_2560),
    .A2(n_2678),
    .B1(n_2543),
    .B2(n_2694),
    .Y(n_2725));
 OAI22xp33_ASAP7_75t_R g52233__2802 (.A1(n_2560),
    .A2(n_2680),
    .B1(n_2543),
    .B2(n_2669),
    .Y(n_2724));
 OAI22xp33_ASAP7_75t_R g52234__1705 (.A1(n_1829),
    .A2(n_2715),
    .B1(n_1830),
    .B2(n_2705),
    .Y(n_2741));
 AOI22xp33_ASAP7_75t_R g52235__5122 (.A1(n_1832),
    .A2(n_2714),
    .B1(n_1833),
    .B2(n_2703),
    .Y(n_2740));
 AOI22xp33_ASAP7_75t_R g52236__8246 (.A1(n_1832),
    .A2(n_2712),
    .B1(n_1833),
    .B2(n_2716),
    .Y(n_2739));
 OAI22xp33_ASAP7_75t_R g52237__7098 (.A1(n_1829),
    .A2(n_2683),
    .B1(n_2501),
    .B2(n_2684),
    .Y(n_2738));
 AOI22xp33_ASAP7_75t_R g52238__6131 (.A1(n_2718),
    .A2(n_1830),
    .B1(n_2712),
    .B2(n_1831),
    .Y(n_2737));
 OAI22xp33_ASAP7_75t_R g52239__1881 (.A1(n_2560),
    .A2(n_2709),
    .B1(n_2677),
    .B2(n_2543),
    .Y(n_2736));
 OAI22xp33_ASAP7_75t_R g52240__5115 (.A1(n_1831),
    .A2(n_2688),
    .B1(n_1832),
    .B2(n_2713),
    .Y(n_2735));
 OAI22xp33_ASAP7_75t_R g52241__7482 (.A1(n_2560),
    .A2(n_2675),
    .B1(n_2543),
    .B2(n_2711),
    .Y(n_2734));
 OAI22xp33_ASAP7_75t_R g52242__4733 (.A1(n_1829),
    .A2(n_2682),
    .B1(n_1830),
    .B2(n_2717),
    .Y(n_2733));
 OAI22xp33_ASAP7_75t_R g52243__6161 (.A1(n_1829),
    .A2(n_2684),
    .B1(n_1830),
    .B2(n_2688),
    .Y(n_2732));
 NOR2xp33_ASAP7_75t_R g52244__9315 (.A(n_2598),
    .B(n_2660),
    .Y(n_2723));
 NAND2xp33_ASAP7_75t_R g52245__9945 (.A(n_2528),
    .B(n_2697),
    .Y(n_2722));
 NOR2xp33_ASAP7_75t_R g52246__2883 (.A(n_2563),
    .B(n_2686),
    .Y(n_2721));
 NOR2xp33_ASAP7_75t_R g52247__2346 (.A(n_2518),
    .B(n_2660),
    .Y(n_2720));
 INVxp33_ASAP7_75t_R g52248 (.A(n_2717),
    .Y(n_2718));
 INVxp33_ASAP7_75t_R g52249 (.A(n_2715),
    .Y(n_2716));
 INVxp33_ASAP7_75t_R g52250 (.A(n_2713),
    .Y(n_2714));
 INVxp33_ASAP7_75t_R g52251 (.A(n_2709),
    .Y(n_2708));
 INVxp33_ASAP7_75t_R g52252 (.A(n_2707),
    .Y(n_2706));
 INVxp33_ASAP7_75t_R g52253 (.A(n_2702),
    .Y(n_2701));
 INVxp33_ASAP7_75t_R g52254 (.A(n_2700),
    .Y(n_2699));
 INVxp33_ASAP7_75t_R g52255 (.A(n_2693),
    .Y(n_2692));
 INVxp33_ASAP7_75t_R g52256 (.A(n_2691),
    .Y(n_2690));
 AOI221xp5_ASAP7_75t_R g52257__1666 (.A1(n_1821),
    .A2(fract_denorm[39]),
    .B1(n_2594),
    .B2(fract_denorm[38]),
    .C(n_2621),
    .Y(n_2719));
 AOI221xp5_ASAP7_75t_R g52258__7410 (.A1(n_1822),
    .A2(fract_denorm[30]),
    .B1(n_2594),
    .B2(fract_denorm[29]),
    .C(n_2636),
    .Y(n_2717));
 AOI221xp5_ASAP7_75t_R g52259__6417 (.A1(n_1821),
    .A2(fract_denorm[22]),
    .B1(n_1823),
    .B2(fract_denorm[21]),
    .C(n_2639),
    .Y(n_2715));
 AOI221xp5_ASAP7_75t_R g52260__5477 (.A1(n_1841),
    .A2(fract_denorm[24]),
    .B1(n_1823),
    .B2(fract_denorm[22]),
    .C(n_2615),
    .Y(n_2713));
 OAI221xp5_ASAP7_75t_R g52261__2398 (.A1(n_2586),
    .A2(n_1911),
    .B1(n_2589),
    .B2(n_1860),
    .C(n_2652),
    .Y(n_2712));
 AOI221xp5_ASAP7_75t_R g52262__5107 (.A1(n_1842),
    .A2(fract_denorm[25]),
    .B1(n_2595),
    .B2(fract_denorm[24]),
    .C(n_2628),
    .Y(n_2711));
 AOI221xp5_ASAP7_75t_R g52263__6260 (.A1(n_1842),
    .A2(fract_denorm[4]),
    .B1(n_1841),
    .B2(fract_denorm[5]),
    .C(n_2623),
    .Y(n_2710));
 AOI221xp5_ASAP7_75t_R g52264__4319 (.A1(n_1822),
    .A2(fract_denorm[32]),
    .B1(n_2594),
    .B2(fract_denorm[31]),
    .C(n_2625),
    .Y(n_2709));
 AOI221xp5_ASAP7_75t_R g52265__8428 (.A1(n_1842),
    .A2(fract_denorm[3]),
    .B1(n_2595),
    .B2(fract_denorm[2]),
    .C(n_2620),
    .Y(n_2707));
 AOI221xp5_ASAP7_75t_R g52266__5526 (.A1(n_1821),
    .A2(fract_denorm[18]),
    .B1(n_1823),
    .B2(fract_denorm[17]),
    .C(n_2637),
    .Y(n_2705));
 OAI221xp5_ASAP7_75t_R g52267__6783 (.A1(n_2592),
    .A2(n_1567),
    .B1(n_2590),
    .B2(n_1925),
    .C(n_2631),
    .Y(n_2704));
 OAI221xp5_ASAP7_75t_R g52268__3680 (.A1(n_2592),
    .A2(n_1855),
    .B1(n_2591),
    .B2(n_1591),
    .C(n_2612),
    .Y(n_2703));
 AOI221xp5_ASAP7_75t_R g52269__1617 (.A1(n_1822),
    .A2(fract_denorm[6]),
    .B1(n_1823),
    .B2(fract_denorm[5]),
    .C(n_2641),
    .Y(n_2702));
 AOI221xp5_ASAP7_75t_R g52270__2802 (.A1(n_1822),
    .A2(fract_denorm[14]),
    .B1(n_2595),
    .B2(fract_denorm[13]),
    .C(n_2638),
    .Y(n_2700));
 OAI221xp5_ASAP7_75t_R g52271__1705 (.A1(n_2592),
    .A2(n_1917),
    .B1(n_1843),
    .B2(n_1568),
    .C(n_2630),
    .Y(n_2698));
 OAI221xp5_ASAP7_75t_R g52272__5122 (.A1(n_2586),
    .A2(n_1913),
    .B1(n_2590),
    .B2(n_1917),
    .C(n_2650),
    .Y(n_2697));
 OAI221xp5_ASAP7_75t_R g52273__8246 (.A1(n_2587),
    .A2(n_1849),
    .B1(n_2590),
    .B2(n_1569),
    .C(n_2651),
    .Y(n_2696));
 OAI221xp5_ASAP7_75t_R g52274__7098 (.A1(n_2587),
    .A2(n_1855),
    .B1(n_2590),
    .B2(n_1853),
    .C(n_2645),
    .Y(n_2695));
 AOI221xp5_ASAP7_75t_R g52275__6131 (.A1(n_1821),
    .A2(fract_denorm[29]),
    .B1(n_2594),
    .B2(fract_denorm[28]),
    .C(n_2627),
    .Y(n_2694));
 AOI221xp5_ASAP7_75t_R g52276__1881 (.A1(n_1822),
    .A2(fract_denorm[10]),
    .B1(n_2595),
    .B2(fract_denorm[9]),
    .C(n_2640),
    .Y(n_2693));
 AOI221xp5_ASAP7_75t_R g52277__5115 (.A1(n_1842),
    .A2(fract_denorm[7]),
    .B1(n_1823),
    .B2(fract_denorm[6]),
    .C(n_2619),
    .Y(n_2691));
 AOI221xp5_ASAP7_75t_R g52278__7482 (.A1(n_1842),
    .A2(fract_denorm[11]),
    .B1(n_1823),
    .B2(fract_denorm[10]),
    .C(n_2618),
    .Y(n_2689));
 INVxp33_ASAP7_75t_R g52279 (.A(n_2680),
    .Y(n_2681));
 INVxp33_ASAP7_75t_R g52280 (.A(n_2678),
    .Y(n_2679));
 INVxp33_ASAP7_75t_R g52281 (.A(n_2675),
    .Y(n_2674));
 INVxp33_ASAP7_75t_R g52282 (.A(n_2673),
    .Y(n_2672));
 INVxp33_ASAP7_75t_R g52283 (.A(n_2671),
    .Y(n_2670));
 INVxp33_ASAP7_75t_R g52284 (.A(n_2668),
    .Y(n_2669));
 INVxp33_ASAP7_75t_R g52285 (.A(n_2666),
    .Y(n_2667));
 INVxp33_ASAP7_75t_R g52286 (.A(n_2665),
    .Y(n_2664));
 INVxp33_ASAP7_75t_R g52287 (.A(n_2663),
    .Y(n_2662));
 INVxp33_ASAP7_75t_R g52288 (.A(n_2659),
    .Y(n_2660));
 OAI22xp33_ASAP7_75t_R g52289__4733 (.A1(n_2563),
    .A2(n_2610),
    .B1(n_2409),
    .B2(n_2504),
    .Y(n_2658));
 AOI221xp5_ASAP7_75t_R g52290__6161 (.A1(n_1839),
    .A2(fract_denorm[44]),
    .B1(n_1836),
    .B2(fract_denorm[45]),
    .C(n_2608),
    .Y(n_2657));
 AOI221xp5_ASAP7_75t_R g52291__9315 (.A1(n_1836),
    .A2(fract_denorm[44]),
    .B1(n_1839),
    .B2(fract_denorm[43]),
    .C(n_2607),
    .Y(n_2656));
 AOI221xp5_ASAP7_75t_R g52292__9945 (.A1(n_1822),
    .A2(fract_denorm[27]),
    .B1(n_2595),
    .B2(fract_denorm[26]),
    .C(n_2614),
    .Y(n_2688));
 OAI21xp33_ASAP7_75t_R g52293__2883 (.A1(n_2545),
    .A2(n_2580),
    .B(n_2644),
    .Y(n_2687));
 AOI221xp5_ASAP7_75t_R g52294__2346 (.A1(n_1822),
    .A2(fract_denorm[38]),
    .B1(n_2594),
    .B2(fract_denorm[37]),
    .C(n_2642),
    .Y(n_2686));
 AOI221xp5_ASAP7_75t_R g52295__1666 (.A1(n_1821),
    .A2(fract_denorm[41]),
    .B1(n_2594),
    .B2(fract_denorm[40]),
    .C(n_2609),
    .Y(n_2685));
 AOI221xp5_ASAP7_75t_R g52296__7410 (.A1(n_1821),
    .A2(fract_denorm[31]),
    .B1(n_2594),
    .B2(fract_denorm[30]),
    .C(n_2617),
    .Y(n_2684));
 AOI221xp5_ASAP7_75t_R g52297__6417 (.A1(n_1821),
    .A2(fract_denorm[35]),
    .B1(n_2594),
    .B2(fract_denorm[34]),
    .C(n_2616),
    .Y(n_2683));
 AOI221xp5_ASAP7_75t_R g52298__5477 (.A1(n_1822),
    .A2(fract_denorm[34]),
    .B1(n_2594),
    .B2(fract_denorm[33]),
    .C(n_2635),
    .Y(n_2682));
 AOI221xp5_ASAP7_75t_R g52299__2398 (.A1(n_1822),
    .A2(fract_denorm[36]),
    .B1(n_2594),
    .B2(fract_denorm[35]),
    .C(n_2624),
    .Y(n_2680));
 AOI221xp5_ASAP7_75t_R g52300__5107 (.A1(n_1821),
    .A2(fract_denorm[37]),
    .B1(n_2594),
    .B2(fract_denorm[36]),
    .C(n_2622),
    .Y(n_2678));
 AOI221xp5_ASAP7_75t_R g52301__6260 (.A1(n_2595),
    .A2(fract_denorm[23]),
    .B1(n_1842),
    .B2(fract_denorm[24]),
    .C(n_2605),
    .Y(n_2677));
 AOI221xp5_ASAP7_75t_R g52302__4319 (.A1(n_1840),
    .A2(fract_denorm[3]),
    .B1(n_1837),
    .B2(fract_denorm[4]),
    .C(n_2600),
    .Y(n_2676));
 AOI221xp5_ASAP7_75t_R g52303__8428 (.A1(n_1821),
    .A2(fract_denorm[33]),
    .B1(n_2594),
    .B2(fract_denorm[32]),
    .C(n_2653),
    .Y(n_2675));
 OAI221xp5_ASAP7_75t_R g52304__5526 (.A1(n_2587),
    .A2(n_1569),
    .B1(n_2591),
    .B2(n_1915),
    .C(n_2649),
    .Y(n_2673));
 OAI221xp5_ASAP7_75t_R g52305__6783 (.A1(n_2590),
    .A2(n_1846),
    .B1(n_1843),
    .B2(n_1591),
    .C(n_2629),
    .Y(n_2671));
 OAI221xp5_ASAP7_75t_R g52306__3680 (.A1(n_2592),
    .A2(n_1911),
    .B1(n_2593),
    .B2(n_1860),
    .C(n_2633),
    .Y(n_2668));
 OAI221xp5_ASAP7_75t_R g52307__1617 (.A1(n_2592),
    .A2(n_1849),
    .B1(n_1843),
    .B2(n_1569),
    .C(n_2613),
    .Y(n_2666));
 OAI221xp5_ASAP7_75t_R g52308__2802 (.A1(n_2588),
    .A2(n_1846),
    .B1(n_2592),
    .B2(n_1591),
    .C(n_2646),
    .Y(n_2665));
 OAI221xp5_ASAP7_75t_R g52309__1705 (.A1(n_2587),
    .A2(n_1853),
    .B1(n_2590),
    .B2(n_1585),
    .C(n_2643),
    .Y(n_2663));
 AOI222xp33_ASAP7_75t_R g52310__5122 (.A1(n_1838),
    .A2(fract_denorm[2]),
    .B1(n_1842),
    .B2(fract_denorm[0]),
    .C1(n_1841),
    .C2(fract_denorm[1]),
    .Y(n_2661));
 OAI21xp33_ASAP7_75t_R g52311__8246 (.A1(n_2546),
    .A2(n_2599),
    .B(n_2632),
    .Y(n_2659));
 INVxp33_ASAP7_75t_R g52312 (.A(n_2655),
    .Y(n_2654));
 OAI22xp33_ASAP7_75t_R g52313__7098 (.A1(n_1576),
    .A2(n_2586),
    .B1(n_1914),
    .B2(n_2589),
    .Y(n_2653));
 AOI22xp33_ASAP7_75t_R g52314__6131 (.A1(fract_denorm[26]),
    .A2(n_1822),
    .B1(fract_denorm[25]),
    .B2(n_2595),
    .Y(n_2652));
 AOI22xp33_ASAP7_75t_R g52315__1881 (.A1(fract_denorm[13]),
    .A2(n_1842),
    .B1(fract_denorm[12]),
    .B2(n_1823),
    .Y(n_2651));
 AOI22xp33_ASAP7_75t_R g52316__5115 (.A1(fract_denorm[8]),
    .A2(n_1842),
    .B1(fract_denorm[7]),
    .B2(n_1823),
    .Y(n_2650));
 AOI22xp33_ASAP7_75t_R g52317__7482 (.A1(fract_denorm[12]),
    .A2(n_1842),
    .B1(fract_denorm[11]),
    .B2(n_2595),
    .Y(n_2649));
 AOI22xp33_ASAP7_75t_R g52318__4733 (.A1(fract_denorm[45]),
    .A2(n_1821),
    .B1(fract_denorm[44]),
    .B2(n_2594),
    .Y(n_2648));
 AOI22xp33_ASAP7_75t_R g52319__6161 (.A1(fract_denorm[44]),
    .A2(n_1821),
    .B1(fract_denorm[43]),
    .B2(n_2594),
    .Y(n_2647));
 AOI22xp33_ASAP7_75t_R g52320__9315 (.A1(fract_denorm[21]),
    .A2(n_1841),
    .B1(fract_denorm[19]),
    .B2(n_2595),
    .Y(n_2646));
 AOI22xp33_ASAP7_75t_R g52321__9945 (.A1(fract_denorm[17]),
    .A2(n_1842),
    .B1(fract_denorm[16]),
    .B2(n_2595),
    .Y(n_2645));
 AOI22xp33_ASAP7_75t_R g52322__2883 (.A1(fract_denorm[40]),
    .A2(n_1821),
    .B1(fract_denorm[39]),
    .B2(n_2594),
    .Y(n_2644));
 AOI22xp33_ASAP7_75t_R g52323__2346 (.A1(fract_denorm[16]),
    .A2(n_1842),
    .B1(fract_denorm[15]),
    .B2(n_1823),
    .Y(n_2643));
 OAI22xp33_ASAP7_75t_R g52324__1666 (.A1(n_1852),
    .A2(n_2586),
    .B1(n_1910),
    .B2(n_2589),
    .Y(n_2642));
 OAI22xp33_ASAP7_75t_R g52325__7410 (.A1(n_1568),
    .A2(n_2587),
    .B1(n_1867),
    .B2(n_2590),
    .Y(n_2641));
 OAI22xp33_ASAP7_75t_R g52326__6417 (.A1(n_1923),
    .A2(n_2587),
    .B1(n_1570),
    .B2(n_2590),
    .Y(n_2640));
 OAI22xp33_ASAP7_75t_R g52327__5477 (.A1(n_1850),
    .A2(n_2587),
    .B1(n_1577),
    .B2(n_2590),
    .Y(n_2639));
 OAI22xp33_ASAP7_75t_R g52328__2398 (.A1(n_1903),
    .A2(n_2587),
    .B1(n_1849),
    .B2(n_2590),
    .Y(n_2638));
 OAI22xp33_ASAP7_75t_R g52329__5107 (.A1(n_1591),
    .A2(n_2587),
    .B1(n_1855),
    .B2(n_2590),
    .Y(n_2637));
 OAI22xp33_ASAP7_75t_R g52330__6260 (.A1(n_1590),
    .A2(n_2586),
    .B1(n_1851),
    .B2(n_2589),
    .Y(n_2636));
 OAI22xp33_ASAP7_75t_R g52331__4319 (.A1(n_1845),
    .A2(n_2586),
    .B1(n_1576),
    .B2(n_2589),
    .Y(n_2635));
 AOI22xp33_ASAP7_75t_R g52332__8428 (.A1(fract_denorm[47]),
    .A2(n_1836),
    .B1(fract_denorm[46]),
    .B2(n_1839),
    .Y(n_2634));
 NAND2xp33_ASAP7_75t_R g52333__5526 (.A(n_1830),
    .B(n_2611),
    .Y(n_2655));
 AOI22xp33_ASAP7_75t_R g52334__6783 (.A1(fract_denorm[30]),
    .A2(n_1836),
    .B1(fract_denorm[29]),
    .B2(n_1839),
    .Y(n_2633));
 AOI22xp33_ASAP7_75t_R g52335__3680 (.A1(fract_denorm[3]),
    .A2(n_1838),
    .B1(fract_denorm[2]),
    .B2(n_1841),
    .Y(n_2632));
 AOI22xp33_ASAP7_75t_R g52336__1617 (.A1(fract_denorm[7]),
    .A2(n_1837),
    .B1(fract_denorm[4]),
    .B2(n_1823),
    .Y(n_2631));
 AOI22xp33_ASAP7_75t_R g52337__2802 (.A1(fract_denorm[11]),
    .A2(n_1836),
    .B1(fract_denorm[10]),
    .B2(n_1840),
    .Y(n_2630));
 AOI22xp33_ASAP7_75t_R g52338__1705 (.A1(fract_denorm[23]),
    .A2(n_1838),
    .B1(fract_denorm[21]),
    .B2(n_1842),
    .Y(n_2629));
 OAI22xp33_ASAP7_75t_R g52339__5122 (.A1(n_2587),
    .A2(n_1860),
    .B1(n_2590),
    .B2(n_1589),
    .Y(n_2628));
 OAI22xp33_ASAP7_75t_R g52340__8246 (.A1(n_1851),
    .A2(n_2586),
    .B1(n_1912),
    .B2(n_2589),
    .Y(n_2627));
 AOI22xp33_ASAP7_75t_R g52341__7098 (.A1(fract_denorm[46]),
    .A2(n_1836),
    .B1(fract_denorm[45]),
    .B2(n_1839),
    .Y(n_2626));
 OAI22xp33_ASAP7_75t_R g52342__6131 (.A1(n_1914),
    .A2(n_2586),
    .B1(n_1916),
    .B2(n_2589),
    .Y(n_2625));
 OAI22xp33_ASAP7_75t_R g52343__1881 (.A1(n_1587),
    .A2(n_2586),
    .B1(n_1900),
    .B2(n_2589),
    .Y(n_2624));
 OAI22xp33_ASAP7_75t_R g52344__5115 (.A1(n_2588),
    .A2(n_1925),
    .B1(n_1843),
    .B2(n_1871),
    .Y(n_2623));
 OAI22xp33_ASAP7_75t_R g52345__7482 (.A1(n_2586),
    .A2(n_1910),
    .B1(n_2589),
    .B2(n_1587),
    .Y(n_2622));
 OAI22xp33_ASAP7_75t_R g52346__4733 (.A1(n_1578),
    .A2(n_2586),
    .B1(n_1852),
    .B2(n_2589),
    .Y(n_2621));
 OAI22xp33_ASAP7_75t_R g52347__6161 (.A1(n_2588),
    .A2(n_1567),
    .B1(n_2591),
    .B2(n_1922),
    .Y(n_2620));
 OAI22xp33_ASAP7_75t_R g52348__9315 (.A1(n_2588),
    .A2(n_1917),
    .B1(n_2591),
    .B2(n_1568),
    .Y(n_2619));
 OAI22xp33_ASAP7_75t_R g52349__9945 (.A1(n_2588),
    .A2(n_1915),
    .B1(n_2591),
    .B2(n_1923),
    .Y(n_2618));
 OAI22xp33_ASAP7_75t_R g52350__2883 (.A1(n_1916),
    .A2(n_2586),
    .B1(n_1590),
    .B2(n_2589),
    .Y(n_2617));
 OAI22xp33_ASAP7_75t_R g52351__2346 (.A1(n_1900),
    .A2(n_2586),
    .B1(n_1845),
    .B2(n_2589),
    .Y(n_2616));
 OAI22xp33_ASAP7_75t_R g52352__1666 (.A1(n_2588),
    .A2(n_1920),
    .B1(n_2592),
    .B2(n_1577),
    .Y(n_2615));
 OAI22xp33_ASAP7_75t_R g52353__7410 (.A1(n_1588),
    .A2(n_2587),
    .B1(n_1911),
    .B2(n_2590),
    .Y(n_2614));
 AOI22xp33_ASAP7_75t_R g52354__6417 (.A1(fract_denorm[17]),
    .A2(n_1838),
    .B1(fract_denorm[16]),
    .B2(n_1841),
    .Y(n_2613));
 AOI22xp33_ASAP7_75t_R g52355__5477 (.A1(fract_denorm[21]),
    .A2(n_1838),
    .B1(fract_denorm[18]),
    .B2(n_2595),
    .Y(n_2612));
 NOR2xp33_ASAP7_75t_R g52357__2398 (.A(n_2545),
    .B(n_2581),
    .Y(n_2609));
 NOR2xp33_ASAP7_75t_R g52358__5107 (.A(n_2546),
    .B(n_2581),
    .Y(n_2608));
 NOR2xp33_ASAP7_75t_R g52359__6260 (.A(n_2546),
    .B(n_2580),
    .Y(n_2607));
 NOR2xp33_ASAP7_75t_R g52360__4319 (.A(n_2545),
    .B(n_2599),
    .Y(n_2611));
 NAND2xp33_ASAP7_75t_R g52361__8428 (.A(fract_denorm[0]),
    .B(n_1837),
    .Y(n_2610));
 OAI22xp33_ASAP7_75t_R g52362__5526 (.A1(n_2502),
    .A2(n_2434),
    .B1(n_2553),
    .B2(n_2311),
    .Y(n_2606));
 O2A1O1Ixp33_ASAP7_75t_R g52363__6783 (.A1(n_1920),
    .A2(n_2523),
    .B(n_2559),
    .C(n_2545),
    .Y(n_2605));
 OAI22xp33_ASAP7_75t_R g52364__3680 (.A1(n_2425),
    .A2(n_2516),
    .B1(n_2316),
    .B2(n_2550),
    .Y(n_2604));
 AOI22xp33_ASAP7_75t_R g52365__1617 (.A1(n_2389),
    .A2(n_2532),
    .B1(n_2304),
    .B2(n_2549),
    .Y(n_2603));
 OAI22xp33_ASAP7_75t_R g52366__2802 (.A1(n_2555),
    .A2(n_2302),
    .B1(n_2547),
    .B2(n_2336),
    .Y(n_2602));
 OAI22xp33_ASAP7_75t_R g52367__1705 (.A1(n_2342),
    .A2(n_2547),
    .B1(n_2302),
    .B2(n_2550),
    .Y(n_2601));
 NOR2xp33_ASAP7_75t_R g52368__5122 (.A(n_2546),
    .B(n_2583),
    .Y(n_2600));
 INVxp33_ASAP7_75t_R g52369 (.A(n_2597),
    .Y(n_2596));
 INVxp33_ASAP7_75t_R g52370 (.A(n_2594),
    .Y(n_2593));
 HB1xp67_ASAP7_75t_R g52371 (.A(n_1823),
    .Y(n_2594));
 INVxp33_ASAP7_75t_R g52381 (.A(n_2592),
    .Y(n_1842));
 INVxp33_ASAP7_75t_R g52383 (.A(n_2591),
    .Y(n_1841));
 INVxp33_ASAP7_75t_R g52390 (.A(n_2589),
    .Y(n_1839));
 HB1xp67_ASAP7_75t_R g52394 (.A(n_2590),
    .Y(n_2589));
 INVxp33_ASAP7_75t_R g52395 (.A(n_2590),
    .Y(n_1840));
 HB1xp67_ASAP7_75t_R g52396 (.A(n_2591),
    .Y(n_2590));
 INVxp33_ASAP7_75t_R g52404 (.A(n_2587),
    .Y(n_1837));
 INVxp33_ASAP7_75t_R g52408 (.A(n_2586),
    .Y(n_1836));
 HB1xp67_ASAP7_75t_R g52410 (.A(n_2587),
    .Y(n_2586));
 HB1xp67_ASAP7_75t_R g52411 (.A(n_2588),
    .Y(n_2587));
 INVxp33_ASAP7_75t_R g52412 (.A(n_2588),
    .Y(n_1838));
 NOR2xp33_ASAP7_75t_R g52413__8246 (.A(n_2313),
    .B(n_2547),
    .Y(n_2585));
 OAI21xp33_ASAP7_75t_R g52414__7098 (.A1(n_2335),
    .A2(n_2314),
    .B(n_2549),
    .Y(n_2584));
 AOI22xp33_ASAP7_75t_R g52415__6131 (.A1(fract_denorm[2]),
    .A2(n_2523),
    .B1(fract_denorm[1]),
    .B2(n_2522),
    .Y(n_2583));
 AOI32xp33_ASAP7_75t_R g52416__1881 (.A1(n_2488),
    .A2(u1_signb_r),
    .A3(opb_nan),
    .B1(n_2513),
    .B2(u1_signa_r),
    .Y(n_2582));
 AOI22xp33_ASAP7_75t_R g52417__5115 (.A1(fract_denorm[1]),
    .A2(n_2523),
    .B1(fract_denorm[0]),
    .B2(n_2522),
    .Y(n_2599));
 NAND2xp33_ASAP7_75t_R g52418__7482 (.A(n_2551),
    .B(n_2528),
    .Y(n_2598));
 NAND2xp33_ASAP7_75t_R g52419__4733 (.A(n_2551),
    .B(n_2493),
    .Y(n_2597));
 NOR2xp33_ASAP7_75t_R g52420__6161 (.A(n_2523),
    .B(n_2546),
    .Y(n_2595));
 NAND2xp33_ASAP7_75t_R g52421__9315 (.A(n_2545),
    .B(n_2523),
    .Y(n_2592));
 NAND2xp33_ASAP7_75t_R g52422__9945 (.A(n_2522),
    .B(n_2546),
    .Y(n_2591));
 NAND2xp33_ASAP7_75t_R g52423__2883 (.A(n_2546),
    .B(n_2523),
    .Y(n_2588));
 AOI21xp33_ASAP7_75t_R g52424__2346 (.A1(n_1834),
    .A2(n_2435),
    .B(n_2557),
    .Y(n_2579));
 AOI21xp33_ASAP7_75t_R g52425__1666 (.A1(n_1834),
    .A2(n_2416),
    .B(n_2541),
    .Y(n_2578));
 AOI22xp33_ASAP7_75t_R g52426__7410 (.A1(n_2410),
    .A2(n_1834),
    .B1(n_2390),
    .B2(n_2534),
    .Y(n_2577));
 AOI22xp33_ASAP7_75t_R g52427__6417 (.A1(n_2415),
    .A2(n_1835),
    .B1(n_2405),
    .B2(n_2503),
    .Y(n_2576));
 AOI22xp33_ASAP7_75t_R g52428__5477 (.A1(n_2433),
    .A2(n_1834),
    .B1(n_2389),
    .B2(n_2534),
    .Y(n_2575));
 AOI22xp33_ASAP7_75t_R g52429__2398 (.A1(n_2436),
    .A2(n_1834),
    .B1(n_2253),
    .B2(n_2537),
    .Y(n_2574));
 AOI22xp33_ASAP7_75t_R g52430__5107 (.A1(n_2420),
    .A2(n_1835),
    .B1(n_2430),
    .B2(n_2503),
    .Y(n_2573));
 AOI22xp33_ASAP7_75t_R g52431__6260 (.A1(n_2419),
    .A2(n_1835),
    .B1(n_2402),
    .B2(n_2503),
    .Y(n_2572));
 AOI22xp33_ASAP7_75t_R g52432__4319 (.A1(n_2406),
    .A2(n_1835),
    .B1(n_2408),
    .B2(n_2503),
    .Y(n_2571));
 AOI22xp33_ASAP7_75t_R g52433__8428 (.A1(n_2523),
    .A2(fract_denorm[43]),
    .B1(n_2522),
    .B2(fract_denorm[42]),
    .Y(n_2581));
 AOI22xp33_ASAP7_75t_R g52434__5526 (.A1(n_2523),
    .A2(fract_denorm[42]),
    .B1(n_2522),
    .B2(fract_denorm[41]),
    .Y(n_2580));
 INVxp33_ASAP7_75t_R g52435 (.A(n_2569),
    .Y(n_2568));
 INVxp33_ASAP7_75t_R g52436 (.A(n_2567),
    .Y(n_2566));
 INVxp33_ASAP7_75t_R g52437 (.A(n_2565),
    .Y(n_2564));
 INVxp33_ASAP7_75t_R g52438 (.A(n_2563),
    .Y(n_2562));
 INVxp33_ASAP7_75t_R g52439 (.A(n_2561),
    .Y(n_2560));
 NAND2xp33_ASAP7_75t_R g52441__6783 (.A(fract_denorm[26]),
    .B(n_2523),
    .Y(n_2559));
 NOR2xp33_ASAP7_75t_R g52442__3680 (.A(n_2431),
    .B(n_2516),
    .Y(n_2558));
 NOR2xp33_ASAP7_75t_R g52443__1617 (.A(n_2295),
    .B(n_2535),
    .Y(n_2557));
 NAND2xp33_ASAP7_75t_R g52444__2802 (.A(n_2528),
    .B(n_2527),
    .Y(n_2570));
 NOR2xp33_ASAP7_75t_R g52445__1705 (.A(n_2494),
    .B(n_2526),
    .Y(n_2569));
 NAND2xp33_ASAP7_75t_R g52446__5122 (.A(n_1835),
    .B(n_2294),
    .Y(n_2567));
 NAND2xp33_ASAP7_75t_R g52447__8246 (.A(n_2530),
    .B(n_2524),
    .Y(n_2565));
 NAND2xp33_ASAP7_75t_R g52448__7098 (.A(n_2524),
    .B(n_2528),
    .Y(n_2563));
 NOR2xp33_ASAP7_75t_R g52449__6131 (.A(n_2494),
    .B(n_1816),
    .Y(n_2561));
 INVxp33_ASAP7_75t_R g52450 (.A(n_2556),
    .Y(n_2555));
 INVxp33_ASAP7_75t_R g52451 (.A(n_2554),
    .Y(n_2553));
 INVxp33_ASAP7_75t_R g52452 (.A(n_2552),
    .Y(n_2551));
 INVxp33_ASAP7_75t_R g52453 (.A(n_2550),
    .Y(n_2549));
 INVxp33_ASAP7_75t_R g52454 (.A(n_2548),
    .Y(n_2547));
 INVxp33_ASAP7_75t_R g52455 (.A(n_2546),
    .Y(n_2545));
 INVxp33_ASAP7_75t_R g52456 (.A(n_2544),
    .Y(n_2543));
 AOI22xp33_ASAP7_75t_R g52457__1881 (.A1(n_2419),
    .A2(n_2503),
    .B1(n_2402),
    .B2(n_2505),
    .Y(n_2542));
 NOR2xp33_ASAP7_75t_R g52458__5115 (.A(n_2301),
    .B(n_2538),
    .Y(n_2541));
 AO21x1_ASAP7_75t_R g52459__7482 (.A1(n_2420),
    .A2(n_2503),
    .B(n_2515),
    .Y(n_2540));
 NOR2xp33_ASAP7_75t_R g52460__4733 (.A(n_2329),
    .B(n_2516),
    .Y(n_2556));
 NOR2xp33_ASAP7_75t_R g52461__6161 (.A(n_2328),
    .B(n_2517),
    .Y(n_2554));
 NAND3xp33_ASAP7_75t_R g52462__9315 (.A(n_2506),
    .B(n_2495),
    .C(n_2499),
    .Y(n_2552));
 NAND2xp33_ASAP7_75t_R g52463__9945 (.A(n_2334),
    .B(n_1834),
    .Y(n_2550));
 NOR2xp33_ASAP7_75t_R g52464__2883 (.A(n_2332),
    .B(n_2516),
    .Y(n_2548));
 AOI211xp5_ASAP7_75t_R g52465__2346 (.A1(n_3820),
    .A2(n_1019),
    .B(n_2511),
    .C(n_2447),
    .Y(n_2546));
 NOR2xp33_ASAP7_75t_R g52466__1666 (.A(n_2493),
    .B(n_1816),
    .Y(n_2544));
 INVxp33_ASAP7_75t_R g52467 (.A(underflow_fmul_d[2]),
    .Y(n_2539));
 INVxp33_ASAP7_75t_R g52468 (.A(n_2537),
    .Y(n_2538));
 INVxp33_ASAP7_75t_R g52469 (.A(n_2535),
    .Y(n_2534));
 INVxp33_ASAP7_75t_R g52470 (.A(n_2533),
    .Y(n_2532));
 INVxp33_ASAP7_75t_R g52471 (.A(n_2531),
    .Y(n_2530));
 INVxp33_ASAP7_75t_R g52472 (.A(n_2529),
    .Y(n_2528));
 INVxp33_ASAP7_75t_R g52473 (.A(n_2527),
    .Y(n_2526));
 INVxp33_ASAP7_75t_R g52474 (.A(n_2525),
    .Y(n_2524));
 NOR2xp33_ASAP7_75t_R g52477__7410 (.A(n_2328),
    .B(n_2502),
    .Y(n_2537));
 NAND2xp33_ASAP7_75t_R g52478__6417 (.A(n_2327),
    .B(n_2505),
    .Y(n_2536));
 NAND2xp33_ASAP7_75t_R g52479__5477 (.A(n_2294),
    .B(n_2503),
    .Y(n_2535));
 NAND2xp33_ASAP7_75t_R g52480__2398 (.A(n_2294),
    .B(n_2505),
    .Y(n_2533));
 NAND2xp33_ASAP7_75t_R g52481__5107 (.A(n_2493),
    .B(n_1833),
    .Y(n_2531));
 NAND2xp33_ASAP7_75t_R g52482__6260 (.A(n_2493),
    .B(n_1832),
    .Y(n_2529));
 NOR2xp33_ASAP7_75t_R g52483__4319 (.A(n_2506),
    .B(n_2508),
    .Y(n_2527));
 NAND2xp33_ASAP7_75t_R g52484__8428 (.A(n_2506),
    .B(n_2507),
    .Y(n_2525));
 INVxp33_ASAP7_75t_R g52485 (.A(n_2523),
    .Y(n_2522));
 INVxp33_ASAP7_75t_R g52486 (.A(n_2521),
    .Y(n_2520));
 INVxp33_ASAP7_75t_R g52487 (.A(n_2519),
    .Y(n_2518));
 INVxp33_ASAP7_75t_R g52494 (.A(n_2516),
    .Y(n_1835));
 HB1xp67_ASAP7_75t_R g52497 (.A(n_2517),
    .Y(n_2516));
 INVxp33_ASAP7_75t_R g52501 (.A(n_2517),
    .Y(n_1834));
 AOI21xp33_ASAP7_75t_R g52505__5526 (.A1(n_2429),
    .A2(n_2428),
    .B(n_2504),
    .Y(n_2515));
 NOR2xp33_ASAP7_75t_R g52506__6783 (.A(n_2422),
    .B(n_2502),
    .Y(n_2514));
 OAI311xp33_ASAP7_75t_R g52507__3680 (.A1(n_2193),
    .A2(u1_fracta_lt_fractb),
    .A3(u1_fracta_eq_fractb),
    .B1(opb_nan),
    .C1(n_2011),
    .Y(n_2513));
 AOI31xp33_ASAP7_75t_R g52508__1617 (.A1(n_2418),
    .A2(n_2417),
    .A3(n_2407),
    .B(n_2502),
    .Y(n_2512));
 OAI211xp5_ASAP7_75t_R g52509__2802 (.A1(n_3820),
    .A2(n_2460),
    .B(n_2491),
    .C(n_2105),
    .Y(n_2511));
 AOI21xp33_ASAP7_75t_R g52510__1705 (.A1(n_2413),
    .A2(n_2421),
    .B(n_2502),
    .Y(n_2510));
 AOI221xp5_ASAP7_75t_R g52511__5122 (.A1(n_2468),
    .A2(n_3595),
    .B1(n_2442),
    .B2(n_3717),
    .C(n_2486),
    .Y(n_2523));
 NOR2xp33_ASAP7_75t_R g52512__8246 (.A(n_2493),
    .B(n_1832),
    .Y(n_2521));
 NOR2xp33_ASAP7_75t_R g52513__7098 (.A(n_2493),
    .B(n_1833),
    .Y(n_2519));
 OR3x1_ASAP7_75t_R g52514__6131 (.A(n_2498),
    .B(n_2395),
    .C(n_2362),
    .Y(n_2517));
 INVxp33_ASAP7_75t_R g52515 (.A(underflow_fmul_d[1]),
    .Y(n_2509));
 INVxp33_ASAP7_75t_R g52516 (.A(n_2507),
    .Y(n_2508));
 NOR3xp33_ASAP7_75t_R g52521__1881 (.A(n_2499),
    .B(n_2481),
    .C(n_2482),
    .Y(n_2507));
 INVxp33_ASAP7_75t_R g52522 (.A(n_2505),
    .Y(n_2504));
 INVxp33_ASAP7_75t_R g52523 (.A(n_2503),
    .Y(n_2502));
 INVxp33_ASAP7_75t_R g52533 (.A(n_2501),
    .Y(n_1829));
 HB1xp67_ASAP7_75t_R g52538 (.A(n_1830),
    .Y(n_2501));
 INVxp33_ASAP7_75t_R g52544 (.A(n_1830),
    .Y(n_1831));
 INVxp33_ASAP7_75t_R g52548 (.A(n_1832),
    .Y(n_1833));
 OR3x1_ASAP7_75t_R g52552__5115 (.A(n_2479),
    .B(u2_exp_tmp1[7]),
    .C(n_2139),
    .Y(n_2500));
 AOI221xp5_ASAP7_75t_R g52553__7482 (.A1(n_2442),
    .A2(n_2110),
    .B1(n_2450),
    .B2(exp_r[4]),
    .C(n_2492),
    .Y(n_2506));
 NOR3xp33_ASAP7_75t_R g52554__4733 (.A(n_2498),
    .B(n_2394),
    .C(n_2362),
    .Y(n_2505));
 NOR3xp33_ASAP7_75t_R g52555__6161 (.A(n_2498),
    .B(n_2395),
    .C(n_2361),
    .Y(n_2503));
 AOI221xp5_ASAP7_75t_R g52556__9315 (.A1(n_2442),
    .A2(n_2113),
    .B1(n_2450),
    .B2(exp_r[2]),
    .C(n_2490),
    .Y(n_1832));
 AND2x2_ASAP7_75t_R g52557__9945 (.A(n_2194),
    .B(n_2485),
    .Y(n_2497));
 OR2x2_ASAP7_75t_R g52558__2883 (.A(n_2194),
    .B(n_2485),
    .Y(n_2496));
 OAI221xp5_ASAP7_75t_R g52561__2346 (.A1(n_2467),
    .A2(n_3523),
    .B1(n_2460),
    .B2(n_1069),
    .C(n_2465),
    .Y(n_2499));
 NOR2xp33_ASAP7_75t_R g52562__1666 (.A(n_2482),
    .B(n_2481),
    .Y(n_2495));
 NAND2xp33_ASAP7_75t_R g52563__7410 (.A(n_2426),
    .B(n_2481),
    .Y(n_2498));
 INVxp33_ASAP7_75t_R g52564 (.A(n_2494),
    .Y(n_2493));
 OAI221xp5_ASAP7_75t_R g52565__6417 (.A1(n_2467),
    .A2(n_3516),
    .B1(n_2460),
    .B2(n_14182),
    .C(n_2453),
    .Y(n_2492));
 AOI221xp5_ASAP7_75t_R g52566__5477 (.A1(n_2445),
    .A2(div_opa_ldz_r2[1]),
    .B1(n_2450),
    .B2(exp_r[1]),
    .C(n_2474),
    .Y(n_2491));
 OAI221xp5_ASAP7_75t_R g52567__2398 (.A1(n_2444),
    .A2(n_1130),
    .B1(n_3824),
    .B2(n_3803),
    .C(n_2480),
    .Y(n_2490));
 AOI221xp5_ASAP7_75t_R g52568__5107 (.A1(fracta_mul[23]),
    .A2(opb_r[30]),
    .B1(fractb_mul[23]),
    .B2(opa_r[30]),
    .C(n_2478),
    .Y(n_2489));
 OAI21xp33_ASAP7_75t_R g52569__6260 (.A1(u1_fracta_eq_fractb),
    .A2(n_2477),
    .B(opa_nan),
    .Y(n_2488));
 AOI22xp33_ASAP7_75t_R g52570__4319 (.A1(u0_snan_r_b),
    .A2(u0_expb_ff),
    .B1(u0_snan_r_a),
    .B2(u0_expa_ff),
    .Y(n_2487));
 OAI31xp33_ASAP7_75t_R g52571__8428 (.A1(n_2468),
    .A2(n_2454),
    .A3(n_2442),
    .B(n_2459),
    .Y(n_2486));
 OAI211xp5_ASAP7_75t_R g52572__5526 (.A1(n_98),
    .A2(n_2467),
    .B(n_2473),
    .C(n_2466),
    .Y(n_2494));
 NAND2xp33_ASAP7_75t_R g52573__6783 (.A(u0_fractb_00),
    .B(u0_expb_00),
    .Y(n_2484));
 OR5x1_ASAP7_75t_R g52574__3680 (.A(n_2455),
    .B(n_2126),
    .C(n_1983),
    .D(fract_denorm[37]),
    .E(fract_denorm[38]),
    .Y(n_2483));
 NAND2xp33_ASAP7_75t_R g52576__1617 (.A(u0_infb_f_r),
    .B(u0_expb_ff),
    .Y(n_2485));
 AOI22xp33_ASAP7_75t_R g52577__2802 (.A1(n_1685),
    .A2(n_2468),
    .B1(n_3771),
    .B2(n_2461),
    .Y(n_2480));
 OAI322xp33_ASAP7_75t_R g52578__1705 (.A1(n_2443),
    .A2(n_1854),
    .A3(n_792),
    .B1(n_2460),
    .B2(n_1968),
    .C1(n_2155),
    .C2(n_3803),
    .Y(n_2482));
 OAI22xp33_ASAP7_75t_R g52579__5122 (.A1(fractb_mul[23]),
    .A2(n_2472),
    .B1(fracta_mul[23]),
    .B2(n_2458),
    .Y(n_2479));
 OAI22xp33_ASAP7_75t_R g52580__8246 (.A1(fractb_mul[23]),
    .A2(n_2471),
    .B1(n_13884),
    .B2(n_2457),
    .Y(n_2478));
 OA21x2_ASAP7_75t_R g52581__7098 (.A1(u4_n_1091),
    .A2(n_2462),
    .B(n_2476),
    .Y(n_2481));
 INVxp33_ASAP7_75t_R g52582 (.A(u1_fracta_lt_fractb),
    .Y(n_2477));
 OAI311xp33_ASAP7_75t_R g52587__6131 (.A1(n_2140),
    .A2(n_13920),
    .A3(n_14180),
    .B1(n_2101),
    .C1(n_2462),
    .Y(n_2476));
 NAND2xp33_ASAP7_75t_R g52588__1881 (.A(n_2166),
    .B(n_2472),
    .Y(n_2475));
 NOR2xp33_ASAP7_75t_R g52589__5115 (.A(n_3514),
    .B(n_2467),
    .Y(n_2474));
 AOI22xp33_ASAP7_75t_R g52590__7482 (.A1(n_3768),
    .A2(n_2461),
    .B1(div_opa_ldz_r2[3]),
    .B2(n_2445),
    .Y(n_2473));
 INVxp33_ASAP7_75t_R g52591 (.A(n_2471),
    .Y(n_2472));
 OR2x2_ASAP7_75t_R g52592__4733 (.A(n_14164),
    .B(n_2463),
    .Y(n_2470));
 OAI321xp33_ASAP7_75t_R g52593__6161 (.A1(n_2452),
    .A2(n_2077),
    .A3(n_2087),
    .B1(n_2084),
    .B2(n_2083),
    .C(n_2211),
    .Y(n_2469));
 NOR2xp33_ASAP7_75t_R g52594__9315 (.A(n_14164),
    .B(n_2464),
    .Y(n_2471));
 INVxp33_ASAP7_75t_R g52595 (.A(n_2468),
    .Y(n_2467));
 AOI221xp5_ASAP7_75t_R g52596__9945 (.A1(n_2450),
    .A2(exp_r[3]),
    .B1(n_3751),
    .B2(n_1019),
    .C(n_2448),
    .Y(n_2466));
 AOI221xp5_ASAP7_75t_R g52597__2883 (.A1(n_2450),
    .A2(n_13946),
    .B1(n_3753),
    .B2(n_1019),
    .C(n_2451),
    .Y(n_2465));
 NAND4xp25_ASAP7_75t_R g52598__2346 (.A(n_2462),
    .B(n_2440),
    .C(n_2099),
    .D(n_3594),
    .Y(n_2468));
 INVxp33_ASAP7_75t_R g52599 (.A(n_2463),
    .Y(n_2464));
 NOR5xp2_ASAP7_75t_R g52600__1666 (.A(n_2439),
    .B(n_14128),
    .C(n_14130),
    .D(n_14126),
    .E(n_3303),
    .Y(n_2463));
 NAND3xp33_ASAP7_75t_R g52601__7410 (.A(n_3495),
    .B(n_3502),
    .C(n_23),
    .Y(n_2462));
 INVxp33_ASAP7_75t_R g52602 (.A(n_2461),
    .Y(n_2460));
 AOI22xp33_ASAP7_75t_R g52603__6417 (.A1(div_opa_ldz_r2[0]),
    .A2(n_2445),
    .B1(n_13972),
    .B2(n_2450),
    .Y(n_2459));
 OAI22xp33_ASAP7_75t_R g52604__5477 (.A1(n_2012),
    .A2(n_2446),
    .B1(n_3850),
    .B2(n_3495),
    .Y(n_2461));
 INVxp33_ASAP7_75t_R g52605 (.A(n_2457),
    .Y(n_2458));
 INVxp33_ASAP7_75t_R g52606 (.A(n_2455),
    .Y(n_2456));
 NOR5xp2_ASAP7_75t_R g52607__2398 (.A(n_2424),
    .B(n_3386),
    .C(n_3432),
    .D(n_3476),
    .E(n_3409),
    .Y(n_2457));
 OAI21xp33_ASAP7_75t_R g52608__5107 (.A1(u4_exp_out1_co),
    .A2(n_3567),
    .B(n_1844),
    .Y(n_2455));
 NAND4xp25_ASAP7_75t_R g52609__6260 (.A(n_2449),
    .B(n_2444),
    .C(n_2105),
    .D(u4_sll_315_50_n_29),
    .Y(n_2454));
 AOI22xp33_ASAP7_75t_R g52610__4319 (.A1(div_opa_ldz_r2[4]),
    .A2(n_2445),
    .B1(n_1019),
    .B2(n_3752),
    .Y(n_2453));
 A2O1A1Ixp33_ASAP7_75t_R g52611__8428 (.A1(n_2153),
    .A2(n_2427),
    .B(n_2169),
    .C(n_2137),
    .Y(n_2452));
 O2A1O1Ixp33_ASAP7_75t_R g52612__5526 (.A1(n_13946),
    .A2(n_1988),
    .B(n_2097),
    .C(n_2443),
    .Y(n_2451));
 OAI21xp33_ASAP7_75t_R g52613__6783 (.A1(u4_exp_out1_co),
    .A2(n_2437),
    .B(n_26),
    .Y(n_3495));
 INVxp33_ASAP7_75t_R g52614 (.A(n_2450),
    .Y(n_2449));
 O2A1O1Ixp33_ASAP7_75t_R g52615__3680 (.A1(n_3569),
    .A2(n_1974),
    .B(n_2096),
    .C(n_2443),
    .Y(n_2448));
 O2A1O1Ixp33_ASAP7_75t_R g52616__1617 (.A1(n_1975),
    .A2(n_3720),
    .B(n_2094),
    .C(n_2443),
    .Y(n_2447));
 NOR3xp33_ASAP7_75t_R g52617__2802 (.A(u4_n_1722),
    .B(n_13919),
    .C(u4_op_dn),
    .Y(n_2450));
 NOR2xp33_ASAP7_75t_R g52619__1705 (.A(n_2134),
    .B(n_2437),
    .Y(n_2446));
 NAND2xp33_ASAP7_75t_R g52620__5122 (.A(u4_n_1722),
    .B(n_2140),
    .Y(n_3567));
 INVxp33_ASAP7_75t_R g52621 (.A(n_2445),
    .Y(n_2444));
 INVxp33_ASAP7_75t_R g52622 (.A(n_2443),
    .Y(n_2442));
 OAI221xp5_ASAP7_75t_R g52623__8246 (.A1(n_2329),
    .A2(n_2275),
    .B1(n_2297),
    .B2(n_2332),
    .C(n_2423),
    .Y(n_2441));
 A2O1A1Ixp33_ASAP7_75t_R g52624__7098 (.A1(n_2013),
    .A2(n_3494),
    .B(n_1844),
    .C(u4_n_1722),
    .Y(n_2440));
 NOR3xp33_ASAP7_75t_R g52625__6131 (.A(u4_n_1722),
    .B(n_3502),
    .C(n_2104),
    .Y(n_2445));
 NAND3xp33_ASAP7_75t_R g52626__1881 (.A(n_2437),
    .B(n_3502),
    .C(n_2103),
    .Y(n_2443));
 OR5x1_ASAP7_75t_R g52627__5115 (.A(n_2367),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .C(n_14136),
    .D(n_14146),
    .E(n_14132),
    .Y(n_2439));
 OAI31xp33_ASAP7_75t_R g52628__7482 (.A1(n_2385),
    .A2(n_3395),
    .A3(n_3409),
    .B(n_802),
    .Y(n_2438));
 INVxp33_ASAP7_75t_R g52629 (.A(n_2437),
    .Y(u4_n_1722));
 NAND5xp2_ASAP7_75t_R g52630__4733 (.A(n_2358),
    .B(n_3724),
    .C(n_3722),
    .D(n_3723),
    .E(n_3726),
    .Y(u4_n_1438));
 NOR5xp2_ASAP7_75t_R g52631__6161 (.A(n_2360),
    .B(n_3721),
    .C(n_3722),
    .D(n_3723),
    .E(n_3724),
    .Y(n_2437));
 INVxp33_ASAP7_75t_R g52632 (.A(n_2432),
    .Y(n_2433));
 INVxp33_ASAP7_75t_R g52633 (.A(n_2430),
    .Y(n_2429));
 OAI322xp33_ASAP7_75t_R g52634__9315 (.A1(n_2357),
    .A2(n_2138),
    .A3(n_1996),
    .B1(n_2088),
    .B2(n_2008),
    .C1(n_2009),
    .C2(n_2082),
    .Y(n_2427));
 AOI222xp33_ASAP7_75t_R g52635__9945 (.A1(n_2359),
    .A2(n_792),
    .B1(n_3811),
    .B2(n_13920),
    .C1(n_13840),
    .C2(exp_r[6]),
    .Y(n_2426));
 AOI321xp33_ASAP7_75t_R g52636__2883 (.A1(n_2330),
    .A2(n_2217),
    .A3(n_1994),
    .B1(n_2312),
    .B2(n_2334),
    .C(n_2388),
    .Y(n_2425));
 OR5x1_ASAP7_75t_R g52637__2346 (.A(n_2326),
    .B(n_3395),
    .C(n_3438),
    .D(n_2896),
    .E(n_3466),
    .Y(n_2424));
 AOI221xp5_ASAP7_75t_R g52638__1666 (.A1(n_2234),
    .A2(fract_denorm[13]),
    .B1(n_1826),
    .B2(fract_denorm[14]),
    .C(n_2403),
    .Y(n_2423));
 OAI222xp33_ASAP7_75t_R g52639__7410 (.A1(n_2337),
    .A2(n_2332),
    .B1(n_2381),
    .B2(n_2293),
    .C1(n_2343),
    .C2(n_2333),
    .Y(n_2436));
 OAI222xp33_ASAP7_75t_R g52640__6417 (.A1(n_2310),
    .A2(n_2332),
    .B1(n_2378),
    .B2(n_2293),
    .C1(n_2345),
    .C2(n_2333),
    .Y(n_2435));
 AOI21xp33_ASAP7_75t_R g52641__5477 (.A1(n_2294),
    .A2(n_2377),
    .B(n_2372),
    .Y(n_2434));
 AOI222xp33_ASAP7_75t_R g52642__2398 (.A1(n_2320),
    .A2(n_2331),
    .B1(n_2338),
    .B2(n_2334),
    .C1(n_2396),
    .C2(n_2294),
    .Y(n_2432));
 AOI222xp33_ASAP7_75t_R g52643__5107 (.A1(n_2322),
    .A2(n_2327),
    .B1(n_2307),
    .B2(n_2330),
    .C1(n_2390),
    .C2(n_2293),
    .Y(n_2431));
 OAI222xp33_ASAP7_75t_R g52644__6260 (.A1(n_2323),
    .A2(n_2328),
    .B1(n_2392),
    .B2(n_2294),
    .C1(n_2310),
    .C2(n_2329),
    .Y(n_2430));
 AOI222xp33_ASAP7_75t_R g52645__4319 (.A1(n_2389),
    .A2(n_2293),
    .B1(n_2320),
    .B2(n_2327),
    .C1(n_2338),
    .C2(n_2330),
    .Y(n_2428));
 INVxp33_ASAP7_75t_R g52646 (.A(n_2414),
    .Y(n_2415));
 INVxp33_ASAP7_75t_R g52647 (.A(n_2411),
    .Y(n_2412));
 INVxp33_ASAP7_75t_R g52648 (.A(n_2408),
    .Y(n_2409));
 AOI21xp33_ASAP7_75t_R g52649__8428 (.A1(n_2375),
    .A2(n_2293),
    .B(n_2373),
    .Y(n_2422));
 AOI222xp33_ASAP7_75t_R g52650__5526 (.A1(n_2314),
    .A2(n_2327),
    .B1(n_2304),
    .B2(n_2330),
    .C1(n_2396),
    .C2(n_2293),
    .Y(n_2421));
 OAI222xp33_ASAP7_75t_R g52651__6783 (.A1(n_2302),
    .A2(n_2328),
    .B1(n_2382),
    .B2(n_2294),
    .C1(n_2336),
    .C2(n_2329),
    .Y(n_2420));
 OAI221xp5_ASAP7_75t_R g52652__3680 (.A1(n_2381),
    .A2(n_2294),
    .B1(n_2303),
    .B2(n_2328),
    .C(n_2363),
    .Y(n_2419));
 AOI21xp33_ASAP7_75t_R g52653__1617 (.A1(n_2397),
    .A2(n_2293),
    .B(n_2374),
    .Y(n_2418));
 AOI222xp33_ASAP7_75t_R g52654__2802 (.A1(n_2335),
    .A2(n_2327),
    .B1(n_2309),
    .B2(n_2330),
    .C1(n_2380),
    .C2(n_2293),
    .Y(n_2417));
 OAI222xp33_ASAP7_75t_R g52655__1705 (.A1(n_2325),
    .A2(n_2332),
    .B1(n_2398),
    .B2(n_2293),
    .C1(n_2344),
    .C2(n_2333),
    .Y(n_2416));
 AOI222xp33_ASAP7_75t_R g52656__5122 (.A1(n_2309),
    .A2(n_2327),
    .B1(n_2330),
    .B2(n_2318),
    .C1(n_2377),
    .C2(n_2293),
    .Y(n_2414));
 OA222x2_ASAP7_75t_R g52657__8246 (.A1(n_2336),
    .A2(n_2328),
    .B1(n_2329),
    .B2(n_2319),
    .C1(n_2378),
    .C2(n_2294),
    .Y(n_2413));
 OAI222xp33_ASAP7_75t_R g52658__7098 (.A1(n_2323),
    .A2(n_2332),
    .B1(n_2382),
    .B2(n_2293),
    .C1(n_2310),
    .C2(n_2333),
    .Y(n_2411));
 OAI21xp33_ASAP7_75t_R g52659__6131 (.A1(n_2293),
    .A2(n_2379),
    .B(n_2370),
    .Y(n_2410));
 OAI22xp33_ASAP7_75t_R g52660__1881 (.A1(n_2293),
    .A2(n_2376),
    .B1(n_2294),
    .B2(n_2391),
    .Y(n_2408));
 INVxp33_ASAP7_75t_R g52661 (.A(n_2406),
    .Y(n_2407));
 INVxp33_ASAP7_75t_R g52662 (.A(n_2404),
    .Y(n_2405));
 OAI222xp33_ASAP7_75t_R g52663__5115 (.A1(n_2233),
    .A2(n_1923),
    .B1(n_2299),
    .B2(n_2328),
    .C1(n_1828),
    .C2(n_1849),
    .Y(n_2403));
 OAI221xp5_ASAP7_75t_R g52664__7482 (.A1(n_2316),
    .A2(n_2328),
    .B1(n_2315),
    .B2(n_2329),
    .C(n_2383),
    .Y(n_2406));
 AOI221xp5_ASAP7_75t_R g52665__4733 (.A1(n_2307),
    .A2(n_2327),
    .B1(n_2346),
    .B2(n_2330),
    .C(n_2364),
    .Y(n_2404));
 INVxp33_ASAP7_75t_R g52666 (.A(n_2400),
    .Y(n_2401));
 OAI222xp33_ASAP7_75t_R g52667__6161 (.A1(n_2337),
    .A2(n_2328),
    .B1(n_2254),
    .B2(n_2332),
    .C1(n_2343),
    .C2(n_2329),
    .Y(n_2402));
 OAI222xp33_ASAP7_75t_R g52668__9315 (.A1(n_2310),
    .A2(n_2328),
    .B1(n_2295),
    .B2(n_2294),
    .C1(n_2345),
    .C2(n_2329),
    .Y(n_2400));
 OA222x2_ASAP7_75t_R g52669__9945 (.A1(n_2325),
    .A2(n_2328),
    .B1(n_2344),
    .B2(n_2329),
    .C1(n_2301),
    .C2(n_2332),
    .Y(n_2399));
 INVxp33_ASAP7_75t_R g52670 (.A(n_2397),
    .Y(n_2398));
 INVxp33_ASAP7_75t_R g52671 (.A(n_2394),
    .Y(n_2395));
 INVxp33_ASAP7_75t_R g52672 (.A(n_2393),
    .Y(n_2392));
 INVxp33_ASAP7_75t_R g52673 (.A(n_2384),
    .Y(n_2391));
 OAI22xp33_ASAP7_75t_R g52674__2883 (.A1(n_2283),
    .A2(n_2328),
    .B1(n_2332),
    .B2(n_2284),
    .Y(n_2388));
 OAI22xp33_ASAP7_75t_R g52675__2346 (.A1(n_2239),
    .A2(n_2342),
    .B1(n_2240),
    .B2(n_2355),
    .Y(n_2387));
 OAI22xp33_ASAP7_75t_R g52676__1666 (.A1(n_2239),
    .A2(n_2324),
    .B1(n_2240),
    .B2(n_2354),
    .Y(n_2386));
 OR5x1_ASAP7_75t_R g52677__7410 (.A(n_2247),
    .B(n_3466),
    .C(n_3476),
    .D(n_3468),
    .E(n_3432),
    .Y(n_2385));
 OAI22xp33_ASAP7_75t_R g52678__6417 (.A1(n_2240),
    .A2(n_2339),
    .B1(n_2241),
    .B2(n_2352),
    .Y(n_2397));
 OAI22xp33_ASAP7_75t_R g52679__5477 (.A1(n_1827),
    .A2(n_2340),
    .B1(n_2241),
    .B2(n_2351),
    .Y(n_2396));
 AOI222xp33_ASAP7_75t_R g52680__2398 (.A1(n_2296),
    .A2(n_1854),
    .B1(n_3816),
    .B2(n_13919),
    .C1(n_2279),
    .C2(n_13946),
    .Y(n_2394));
 OAI22xp33_ASAP7_75t_R g52681__5107 (.A1(n_1827),
    .A2(n_2345),
    .B1(n_2241),
    .B2(n_2257),
    .Y(n_2393));
 OAI22xp33_ASAP7_75t_R g52682__6260 (.A1(n_2240),
    .A2(n_2344),
    .B1(n_2239),
    .B2(n_2301),
    .Y(n_2384));
 OAI22xp33_ASAP7_75t_R g52683__4319 (.A1(n_1827),
    .A2(n_2347),
    .B1(n_2241),
    .B2(n_2300),
    .Y(n_2390));
 OAI22xp33_ASAP7_75t_R g52684__8428 (.A1(n_1827),
    .A2(n_2343),
    .B1(n_2241),
    .B2(n_2254),
    .Y(n_2389));
 INVxp33_ASAP7_75t_R g52685 (.A(n_2371),
    .Y(n_2383));
 INVxp33_ASAP7_75t_R g52686 (.A(n_2369),
    .Y(n_2382));
 INVxp33_ASAP7_75t_R g52687 (.A(n_2379),
    .Y(n_2380));
 INVxp33_ASAP7_75t_R g52688 (.A(n_2368),
    .Y(n_2378));
 INVxp33_ASAP7_75t_R g52689 (.A(n_2375),
    .Y(n_2376));
 OAI22xp33_ASAP7_75t_R g52690__5526 (.A1(n_2328),
    .A2(n_2315),
    .B1(n_2329),
    .B2(n_2305),
    .Y(n_2374));
 OAI22xp33_ASAP7_75t_R g52691__6783 (.A1(n_2329),
    .A2(n_2339),
    .B1(n_2328),
    .B2(n_2305),
    .Y(n_2373));
 OAI22xp33_ASAP7_75t_R g52692__3680 (.A1(n_2332),
    .A2(n_2306),
    .B1(n_2333),
    .B2(n_2347),
    .Y(n_2372));
 OAI22xp33_ASAP7_75t_R g52693__1617 (.A1(n_2333),
    .A2(n_2339),
    .B1(n_2332),
    .B2(n_2305),
    .Y(n_2371));
 AOI22xp33_ASAP7_75t_R g52694__2802 (.A1(n_2331),
    .A2(n_2322),
    .B1(n_2334),
    .B2(n_2307),
    .Y(n_2370));
 OAI22xp33_ASAP7_75t_R g52695__1705 (.A1(n_2241),
    .A2(n_2356),
    .B1(n_2240),
    .B2(n_2319),
    .Y(n_2369));
 AOI22xp33_ASAP7_75t_R g52696__5122 (.A1(n_2239),
    .A2(n_2350),
    .B1(n_2240),
    .B2(n_2320),
    .Y(n_2381));
 AOI22xp33_ASAP7_75t_R g52697__8246 (.A1(n_1827),
    .A2(n_2348),
    .B1(n_2241),
    .B2(n_2318),
    .Y(n_2379));
 OAI22xp33_ASAP7_75t_R g52698__7098 (.A1(n_2356),
    .A2(n_2240),
    .B1(n_2323),
    .B2(n_2239),
    .Y(n_2368));
 OAI22xp33_ASAP7_75t_R g52699__6131 (.A1(n_2240),
    .A2(n_2349),
    .B1(n_2239),
    .B2(n_2321),
    .Y(n_2377));
 OAI22xp33_ASAP7_75t_R g52700__1881 (.A1(n_2240),
    .A2(n_2352),
    .B1(n_2239),
    .B2(n_2325),
    .Y(n_2375));
 OR5x1_ASAP7_75t_R g52701__5115 (.A(n_2231),
    .B(n_14160),
    .C(u5_mul_69_18_n_143),
    .D(n_14156),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(n_2367));
 NOR4xp25_ASAP7_75t_R g52703__4733 (.A(n_2249),
    .B(n_1994),
    .C(fract_denorm[4]),
    .D(fract_denorm[3]),
    .Y(n_2365));
 NOR2xp33_ASAP7_75t_R g52704__6161 (.A(n_2332),
    .B(n_2300),
    .Y(n_2364));
 NAND2xp33_ASAP7_75t_R g52705__9315 (.A(n_2330),
    .B(n_2341),
    .Y(n_2363));
 NAND2xp33_ASAP7_75t_R g52706__9945 (.A(n_1844),
    .B(n_3556),
    .Y(n_3555));
 INVxp33_ASAP7_75t_R g52707 (.A(n_2362),
    .Y(n_2361));
 OR4x1_ASAP7_75t_R g52708__2883 (.A(n_3725),
    .B(n_3726),
    .C(u4_exp_out[0]),
    .D(u4_exp_out[7]),
    .Y(n_2360));
 AO21x1_ASAP7_75t_R g52709__2346 (.A1(n_13946),
    .A2(n_2296),
    .B(exp_r[7]),
    .Y(n_2359));
 AND4x1_ASAP7_75t_R g52710__1666 (.A(n_3721),
    .B(n_3725),
    .C(n_2255),
    .D(u4_exp_out[7]),
    .Y(n_2358));
 NOR3xp33_ASAP7_75t_R g52711__7410 (.A(n_2277),
    .B(n_2015),
    .C(n_2010),
    .Y(n_2357));
 OAI311xp33_ASAP7_75t_R g52712__6417 (.A1(u4_exp_zero),
    .A2(n_2162),
    .A3(n_1936),
    .B1(n_3562),
    .C1(n_2285),
    .Y(n_3723));
 OAI21xp33_ASAP7_75t_R g52713__5477 (.A1(n_2207),
    .A2(n_2136),
    .B(n_2298),
    .Y(n_2362));
 INVxp33_ASAP7_75t_R g52714 (.A(n_2353),
    .Y(n_2354));
 INVxp33_ASAP7_75t_R g52715 (.A(n_2350),
    .Y(n_2351));
 INVxp33_ASAP7_75t_R g52716 (.A(n_2348),
    .Y(n_2349));
 INVxp33_ASAP7_75t_R g52717 (.A(n_2346),
    .Y(n_2347));
 INVxp33_ASAP7_75t_R g52718 (.A(n_2341),
    .Y(n_2340));
 INVxp33_ASAP7_75t_R g52719 (.A(n_2338),
    .Y(n_2337));
 INVxp33_ASAP7_75t_R g52720 (.A(n_2334),
    .Y(n_2333));
 INVxp33_ASAP7_75t_R g52721 (.A(n_2332),
    .Y(n_2331));
 INVxp33_ASAP7_75t_R g52722 (.A(n_2330),
    .Y(n_2329));
 INVxp33_ASAP7_75t_R g52723 (.A(n_2328),
    .Y(n_2327));
 OR4x1_ASAP7_75t_R g52724__2398 (.A(n_2232),
    .B(n_2079),
    .C(n_3468),
    .D(n_3434),
    .Y(n_2326));
 AOI221xp5_ASAP7_75t_R g52725__5107 (.A1(n_2235),
    .A2(fract_denorm[31]),
    .B1(n_2244),
    .B2(fract_denorm[33]),
    .C(n_2264),
    .Y(n_2356));
 AOI221xp5_ASAP7_75t_R g52726__6260 (.A1(n_1826),
    .A2(fract_denorm[13]),
    .B1(n_2243),
    .B2(fract_denorm[14]),
    .C(fract_denorm[11]),
    .Y(n_2355));
 OAI221xp5_ASAP7_75t_R g52727__4319 (.A1(n_2233),
    .A2(n_1913),
    .B1(n_1828),
    .B2(n_1915),
    .C(n_1923),
    .Y(n_2353));
 AOI221xp5_ASAP7_75t_R g52728__8428 (.A1(n_2235),
    .A2(fract_denorm[33]),
    .B1(n_2243),
    .B2(fract_denorm[35]),
    .C(n_2266),
    .Y(n_2352));
 OAI221xp5_ASAP7_75t_R g52729__5526 (.A1(n_1820),
    .A2(n_1851),
    .B1(n_2237),
    .B2(n_1916),
    .C(n_2289),
    .Y(n_2350));
 OAI221xp5_ASAP7_75t_R g52730__6783 (.A1(n_1820),
    .A2(n_1588),
    .B1(n_2237),
    .B2(n_1851),
    .C(n_2288),
    .Y(n_2348));
 OAI221xp5_ASAP7_75t_R g52731__3680 (.A1(n_2233),
    .A2(n_1578),
    .B1(n_2237),
    .B2(n_1861),
    .C(n_2287),
    .Y(n_2346));
 AOI221xp5_ASAP7_75t_R g52732__1617 (.A1(n_1819),
    .A2(fract_denorm[43]),
    .B1(n_2244),
    .B2(fract_denorm[45]),
    .C(n_2272),
    .Y(n_2345));
 AOI221xp5_ASAP7_75t_R g52733__2802 (.A1(n_1819),
    .A2(fract_denorm[41]),
    .B1(n_2243),
    .B2(fract_denorm[43]),
    .C(n_2271),
    .Y(n_2344));
 AOI221xp5_ASAP7_75t_R g52734__1705 (.A1(n_2235),
    .A2(fract_denorm[44]),
    .B1(n_2244),
    .B2(fract_denorm[46]),
    .C(n_2273),
    .Y(n_2343));
 AOI221xp5_ASAP7_75t_R g52735__5122 (.A1(n_1824),
    .A2(fract_denorm[15]),
    .B1(n_2234),
    .B2(fract_denorm[16]),
    .C(n_2274),
    .Y(n_2342));
 OAI311xp33_ASAP7_75t_R g52736__8246 (.A1(u4_exp_zero),
    .A2(n_2162),
    .A3(n_1935),
    .B1(n_3562),
    .C1(n_2246),
    .Y(n_3724));
 OAI221xp5_ASAP7_75t_R g52737__7098 (.A1(n_2233),
    .A2(n_1860),
    .B1(n_2237),
    .B2(n_1588),
    .C(n_2291),
    .Y(n_2341));
 AOI221xp5_ASAP7_75t_R g52738__6131 (.A1(n_1819),
    .A2(fract_denorm[29]),
    .B1(n_2243),
    .B2(fract_denorm[31]),
    .C(n_2263),
    .Y(n_2339));
 OAI221xp5_ASAP7_75t_R g52739__1881 (.A1(n_1820),
    .A2(n_1910),
    .B1(n_2236),
    .B2(n_1578),
    .C(n_2290),
    .Y(n_2338));
 AOI221xp5_ASAP7_75t_R g52740__5115 (.A1(n_1824),
    .A2(fract_denorm[22]),
    .B1(n_2234),
    .B2(fract_denorm[23]),
    .C(n_2261),
    .Y(n_2336));
 OAI221xp5_ASAP7_75t_R g52741__7482 (.A1(n_2236),
    .A2(n_1855),
    .B1(n_1828),
    .B2(n_1591),
    .C(n_2282),
    .Y(n_2335));
 NOR2xp33_ASAP7_75t_R g52742__4733 (.A(n_2294),
    .B(n_2239),
    .Y(n_2334));
 NAND2xp33_ASAP7_75t_R g52743__6161 (.A(n_2241),
    .B(n_2293),
    .Y(n_2332));
 NOR2xp33_ASAP7_75t_R g52744__9315 (.A(n_2293),
    .B(n_2239),
    .Y(n_2330));
 NAND2xp33_ASAP7_75t_R g52745__9945 (.A(n_2294),
    .B(n_2241),
    .Y(n_2328));
 INVxp33_ASAP7_75t_R g52746 (.A(n_2322),
    .Y(n_2321));
 INVxp33_ASAP7_75t_R g52747 (.A(n_2317),
    .Y(n_2316));
 INVxp33_ASAP7_75t_R g52748 (.A(n_2314),
    .Y(n_2313));
 INVxp33_ASAP7_75t_R g52749 (.A(n_2312),
    .Y(n_2311));
 INVxp33_ASAP7_75t_R g52750 (.A(n_2309),
    .Y(n_2308));
 INVxp33_ASAP7_75t_R g52751 (.A(n_2307),
    .Y(n_2306));
 INVxp33_ASAP7_75t_R g52752 (.A(n_2304),
    .Y(n_2303));
 AOI222xp33_ASAP7_75t_R g52753__2883 (.A1(n_1824),
    .A2(fract_denorm[0]),
    .B1(n_2234),
    .B2(fract_denorm[1]),
    .C1(n_1826),
    .C2(fract_denorm[2]),
    .Y(n_2299));
 AOI211xp5_ASAP7_75t_R g52754__2346 (.A1(n_3826),
    .A2(n_13919),
    .B(n_2173),
    .C(n_2245),
    .Y(n_2298));
 AOI222xp33_ASAP7_75t_R g52755__1666 (.A1(n_2234),
    .A2(fract_denorm[9]),
    .B1(n_1826),
    .B2(fract_denorm[10]),
    .C1(n_1817),
    .C2(fract_denorm[8]),
    .Y(n_2297));
 OR5x1_ASAP7_75t_R g52756__7410 (.A(n_2258),
    .B(remainder[9]),
    .C(remainder[10]),
    .D(remainder[11]),
    .E(remainder[12]),
    .Y(n_3556));
 AOI221xp5_ASAP7_75t_R g52757__6417 (.A1(n_2235),
    .A2(fract_denorm[37]),
    .B1(n_2243),
    .B2(fract_denorm[39]),
    .C(n_2268),
    .Y(n_2325));
 AOI221xp5_ASAP7_75t_R g52758__5477 (.A1(n_1824),
    .A2(fract_denorm[14]),
    .B1(n_2234),
    .B2(fract_denorm[15]),
    .C(n_2262),
    .Y(n_2324));
 AOI221xp5_ASAP7_75t_R g52759__2398 (.A1(n_1819),
    .A2(fract_denorm[35]),
    .B1(n_2244),
    .B2(fract_denorm[37]),
    .C(n_2267),
    .Y(n_2323));
 OAI221xp5_ASAP7_75t_R g52760__5107 (.A1(n_1820),
    .A2(n_1916),
    .B1(n_2237),
    .B2(n_1576),
    .C(n_2259),
    .Y(n_2322));
 OAI221xp5_ASAP7_75t_R g52761__6260 (.A1(n_2233),
    .A2(n_1576),
    .B1(n_2236),
    .B2(n_1900),
    .C(n_2276),
    .Y(n_2320));
 AOI221xp5_ASAP7_75t_R g52762__4319 (.A1(n_1826),
    .A2(fract_denorm[28]),
    .B1(n_2244),
    .B2(fract_denorm[29]),
    .C(n_2250),
    .Y(n_2319));
 OAI222xp33_ASAP7_75t_R g52763__8428 (.A1(n_2227),
    .A2(n_2218),
    .B1(n_2237),
    .B2(n_1860),
    .C1(n_2242),
    .C2(n_1911),
    .Y(n_2318));
 OAI221xp5_ASAP7_75t_R g52764__5526 (.A1(n_2236),
    .A2(n_1853),
    .B1(n_1828),
    .B2(n_1855),
    .C(n_2281),
    .Y(n_2317));
 AOI221xp5_ASAP7_75t_R g52765__6783 (.A1(n_1817),
    .A2(fract_denorm[20]),
    .B1(n_2234),
    .B2(fract_denorm[21]),
    .C(n_2260),
    .Y(n_2315));
 OAI221xp5_ASAP7_75t_R g52766__3680 (.A1(n_2233),
    .A2(n_1855),
    .B1(n_1825),
    .B2(n_1591),
    .C(n_2270),
    .Y(n_2314));
 OAI221xp5_ASAP7_75t_R g52767__1617 (.A1(n_2236),
    .A2(n_1849),
    .B1(n_1828),
    .B2(n_1903),
    .C(n_2280),
    .Y(n_2312));
 AOI221xp5_ASAP7_75t_R g52768__2802 (.A1(n_2235),
    .A2(fract_denorm[39]),
    .B1(n_2244),
    .B2(fract_denorm[41]),
    .C(n_2269),
    .Y(n_2310));
 OAI221xp5_ASAP7_75t_R g52769__1705 (.A1(n_2236),
    .A2(n_1577),
    .B1(n_1828),
    .B2(n_1850),
    .C(n_2286),
    .Y(n_2309));
 OAI221xp5_ASAP7_75t_R g52770__5122 (.A1(n_1820),
    .A2(n_1900),
    .B1(n_2237),
    .B2(n_1910),
    .C(n_2292),
    .Y(n_2307));
 AOI221xp5_ASAP7_75t_R g52771__8246 (.A1(n_1817),
    .A2(fract_denorm[24]),
    .B1(n_2234),
    .B2(fract_denorm[25]),
    .C(n_2251),
    .Y(n_2305));
 OAI222xp33_ASAP7_75t_R g52772__7098 (.A1(n_2227),
    .A2(n_2217),
    .B1(n_2233),
    .B2(n_1577),
    .C1(n_1825),
    .C2(n_1850),
    .Y(n_2304));
 AOI221xp5_ASAP7_75t_R g52773__6131 (.A1(n_1824),
    .A2(fract_denorm[18]),
    .B1(n_2234),
    .B2(fract_denorm[19]),
    .C(n_2265),
    .Y(n_2302));
 AOI221xp5_ASAP7_75t_R g52774__1881 (.A1(n_1824),
    .A2(fract_denorm[44]),
    .B1(n_2235),
    .B2(fract_denorm[45]),
    .C(n_2252),
    .Y(n_2301));
 AOI222xp33_ASAP7_75t_R g52775__5115 (.A1(n_1819),
    .A2(fract_denorm[46]),
    .B1(n_1824),
    .B2(fract_denorm[45]),
    .C1(n_2238),
    .C2(fract_denorm[47]),
    .Y(n_2300));
 INVxp33_ASAP7_75t_R g52776 (.A(n_2294),
    .Y(n_2293));
 AOI22xp33_ASAP7_75t_R g52777__7482 (.A1(fract_denorm[38]),
    .A2(n_1819),
    .B1(fract_denorm[40]),
    .B2(n_2244),
    .Y(n_2292));
 AOI22xp33_ASAP7_75t_R g52778__4733 (.A1(fract_denorm[28]),
    .A2(n_2235),
    .B1(fract_denorm[30]),
    .B2(n_2244),
    .Y(n_2291));
 AOI22xp33_ASAP7_75t_R g52779__6161 (.A1(fract_denorm[40]),
    .A2(n_1819),
    .B1(fract_denorm[42]),
    .B2(n_2244),
    .Y(n_2290));
 AOI22xp33_ASAP7_75t_R g52780__9315 (.A1(fract_denorm[32]),
    .A2(n_1819),
    .B1(fract_denorm[34]),
    .B2(n_2244),
    .Y(n_2289));
 AOI22xp33_ASAP7_75t_R g52781__9945 (.A1(fract_denorm[30]),
    .A2(n_2235),
    .B1(fract_denorm[32]),
    .B2(n_2244),
    .Y(n_2288));
 AOI22xp33_ASAP7_75t_R g52782__2883 (.A1(fract_denorm[42]),
    .A2(n_1819),
    .B1(fract_denorm[44]),
    .B2(n_2244),
    .Y(n_2287));
 AOI22xp33_ASAP7_75t_R g52783__2346 (.A1(fract_denorm[21]),
    .A2(n_1817),
    .B1(fract_denorm[22]),
    .B2(n_2234),
    .Y(n_2286));
 AOI222xp33_ASAP7_75t_R g52784__1666 (.A1(n_3746),
    .A2(n_3597),
    .B1(u4_exp_div[3]),
    .B2(n_1844),
    .C1(n_2057),
    .C2(n_3598),
    .Y(n_2285));
 AOI22xp33_ASAP7_75t_R g52785__7410 (.A1(fract_denorm[9]),
    .A2(n_1817),
    .B1(fract_denorm[10]),
    .B2(n_2234),
    .Y(n_2284));
 AOI22xp33_ASAP7_75t_R g52786__6417 (.A1(fract_denorm[1]),
    .A2(n_1824),
    .B1(fract_denorm[2]),
    .B2(n_2234),
    .Y(n_2283));
 AOI22xp33_ASAP7_75t_R g52787__5477 (.A1(fract_denorm[17]),
    .A2(n_1824),
    .B1(fract_denorm[18]),
    .B2(n_2234),
    .Y(n_2282));
 AOI22xp33_ASAP7_75t_R g52788__2398 (.A1(fract_denorm[16]),
    .A2(n_1824),
    .B1(fract_denorm[17]),
    .B2(n_2234),
    .Y(n_2281));
 AOI22xp33_ASAP7_75t_R g52789__5107 (.A1(fract_denorm[13]),
    .A2(n_1817),
    .B1(fract_denorm[14]),
    .B2(n_2234),
    .Y(n_2280));
 OAI22xp33_ASAP7_75t_R g52791__6260 (.A1(n_2101),
    .A2(n_2229),
    .B1(n_2089),
    .B2(n_2149),
    .Y(n_2296));
 NAND2xp33_ASAP7_75t_R g52792__4319 (.A(n_3562),
    .B(n_2248),
    .Y(n_3721));
 OAI311xp33_ASAP7_75t_R g52793__8428 (.A1(u4_exp_zero),
    .A2(n_2162),
    .A3(n_1945),
    .B1(n_2025),
    .C1(n_2225),
    .Y(n_3726));
 OAI311xp33_ASAP7_75t_R g52794__5526 (.A1(u4_exp_zero),
    .A2(n_2162),
    .A3(n_1943),
    .B1(n_2025),
    .C1(n_2222),
    .Y(n_3725));
 OAI311xp33_ASAP7_75t_R g52795__6783 (.A1(u4_exp_zero),
    .A2(n_2162),
    .A3(n_3805),
    .B1(n_3562),
    .C1(n_2220),
    .Y(n_3722));
 NAND2xp33_ASAP7_75t_R g52796__3680 (.A(n_2239),
    .B(n_2256),
    .Y(n_2295));
 AOI211xp5_ASAP7_75t_R g52797__1617 (.A1(n_3822),
    .A2(n_13920),
    .B(n_13842),
    .C(n_2230),
    .Y(n_2294));
 INVxp33_ASAP7_75t_R g52798 (.A(n_2278),
    .Y(n_2279));
 OAI221xp5_ASAP7_75t_R g52799__2802 (.A1(n_2085),
    .A2(n_2016),
    .B1(n_1999),
    .B2(n_2027),
    .C(n_2223),
    .Y(n_2277));
 AOI22xp33_ASAP7_75t_R g52800__1705 (.A1(fract_denorm[36]),
    .A2(n_1819),
    .B1(fract_denorm[38]),
    .B2(n_2244),
    .Y(n_2276));
 AOI22xp33_ASAP7_75t_R g52801__5122 (.A1(fract_denorm[4]),
    .A2(n_1817),
    .B1(fract_denorm[6]),
    .B2(n_1826),
    .Y(n_2275));
 OAI22xp33_ASAP7_75t_R g52802__8246 (.A1(n_1585),
    .A2(n_2236),
    .B1(n_1853),
    .B2(n_1828),
    .Y(n_2274));
 OAI22xp33_ASAP7_75t_R g52803__7098 (.A1(n_1861),
    .A2(n_1820),
    .B1(n_1918),
    .B2(n_2237),
    .Y(n_2273));
 OAI22xp33_ASAP7_75t_R g52804__6131 (.A1(n_1866),
    .A2(n_1820),
    .B1(n_1586),
    .B2(n_2237),
    .Y(n_2272));
 OAI22xp33_ASAP7_75t_R g52805__1881 (.A1(n_1852),
    .A2(n_2233),
    .B1(n_1866),
    .B2(n_2236),
    .Y(n_2271));
 AOI22xp33_ASAP7_75t_R g52806__5115 (.A1(fract_denorm[21]),
    .A2(n_1826),
    .B1(fract_denorm[22]),
    .B2(n_2243),
    .Y(n_2270));
 OAI22xp33_ASAP7_75t_R g52807__7482 (.A1(n_1587),
    .A2(n_2233),
    .B1(n_1852),
    .B2(n_2237),
    .Y(n_2269));
 OAI22xp33_ASAP7_75t_R g52808__4733 (.A1(n_1845),
    .A2(n_1820),
    .B1(n_1587),
    .B2(n_2236),
    .Y(n_2268));
 OAI22xp33_ASAP7_75t_R g52809__6161 (.A1(n_1914),
    .A2(n_1820),
    .B1(n_1845),
    .B2(n_2237),
    .Y(n_2267));
 OAI22xp33_ASAP7_75t_R g52810__9315 (.A1(n_1590),
    .A2(n_2233),
    .B1(n_1914),
    .B2(n_2237),
    .Y(n_2266));
 OAI22xp33_ASAP7_75t_R g52811__9945 (.A1(n_1591),
    .A2(n_2236),
    .B1(n_1847),
    .B2(n_1828),
    .Y(n_2265));
 OAI22xp33_ASAP7_75t_R g52812__2883 (.A1(n_1912),
    .A2(n_2233),
    .B1(n_1590),
    .B2(n_2237),
    .Y(n_2264));
 OAI22xp33_ASAP7_75t_R g52813__2346 (.A1(n_1911),
    .A2(n_2233),
    .B1(n_1912),
    .B2(n_2236),
    .Y(n_2263));
 OAI22xp33_ASAP7_75t_R g52814__1666 (.A1(n_1903),
    .A2(n_2236),
    .B1(n_1585),
    .B2(n_1828),
    .Y(n_2262));
 OAI22xp33_ASAP7_75t_R g52815__7410 (.A1(n_1850),
    .A2(n_2236),
    .B1(n_1920),
    .B2(n_1828),
    .Y(n_2261));
 OAI22xp33_ASAP7_75t_R g52816__6417 (.A1(n_1846),
    .A2(n_2236),
    .B1(n_1577),
    .B2(n_1828),
    .Y(n_2260));
 AOI22xp33_ASAP7_75t_R g52817__5477 (.A1(fract_denorm[34]),
    .A2(n_2235),
    .B1(fract_denorm[36]),
    .B2(n_2244),
    .Y(n_2259));
 OR5x1_ASAP7_75t_R g52818__2398 (.A(n_2214),
    .B(remainder[14]),
    .C(remainder[8]),
    .D(remainder[15]),
    .E(remainder[13]),
    .Y(n_2258));
 AOI22xp33_ASAP7_75t_R g52819__5107 (.A1(n_2102),
    .A2(n_2229),
    .B1(n_2089),
    .B2(n_2148),
    .Y(n_2278));
 INVxp33_ASAP7_75t_R g52820 (.A(n_2256),
    .Y(n_2257));
 INVxp33_ASAP7_75t_R g52821 (.A(u4_exp_out[0]),
    .Y(n_2255));
 INVxp33_ASAP7_75t_R g52822 (.A(n_2254),
    .Y(n_2253));
 NOR2xp33_ASAP7_75t_R g52823__6260 (.A(n_2217),
    .B(n_2228),
    .Y(n_2252));
 NOR2xp33_ASAP7_75t_R g52824__4319 (.A(n_2217),
    .B(n_2226),
    .Y(n_2251));
 NOR2xp33_ASAP7_75t_R g52825__8428 (.A(n_2218),
    .B(n_2226),
    .Y(n_2250));
 NOR2xp33_ASAP7_75t_R g52826__5526 (.A(n_2218),
    .B(n_2228),
    .Y(n_2256));
 NAND2xp33_ASAP7_75t_R g52827__6783 (.A(n_3513),
    .B(n_2221),
    .Y(u4_exp_out[0]));
 NAND2xp33_ASAP7_75t_R g52828__3680 (.A(fract_denorm[47]),
    .B(n_1824),
    .Y(n_2254));
 NOR2xp33_ASAP7_75t_R g52829__1617 (.A(n_1571),
    .B(n_2233),
    .Y(n_2249));
 AOI221xp5_ASAP7_75t_R g52830__2802 (.A1(n_3766),
    .A2(n_3598),
    .B1(n_3744),
    .B2(n_3597),
    .C(n_2212),
    .Y(n_2248));
 OR5x1_ASAP7_75t_R g52831__1705 (.A(n_2210),
    .B(n_3566),
    .C(n_2079),
    .D(n_3570),
    .E(n_3434),
    .Y(n_2247));
 AOI221xp5_ASAP7_75t_R g52832__5122 (.A1(u4_exp_div[4]),
    .A2(n_1844),
    .B1(n_3747),
    .B2(n_3597),
    .C(n_2128),
    .Y(n_2246));
 O2A1O1Ixp33_ASAP7_75t_R g52833__8246 (.A1(n_1977),
    .A2(n_2205),
    .B(n_2216),
    .C(n_2101),
    .Y(n_2245));
 OR2x2_ASAP7_75t_R g52834__7098 (.A(n_2077),
    .B(n_2224),
    .Y(u1_n_4702));
 INVxp33_ASAP7_75t_R g52844 (.A(n_2243),
    .Y(n_1828));
 HB1xp67_ASAP7_75t_R g52846 (.A(n_2244),
    .Y(n_2243));
 INVxp33_ASAP7_75t_R g52847 (.A(n_2244),
    .Y(n_2242));
 INVxp33_ASAP7_75t_R g52850 (.A(n_2241),
    .Y(n_1827));
 INVxp33_ASAP7_75t_R g52851 (.A(n_2239),
    .Y(n_2240));
 HB1xp67_ASAP7_75t_R g52859 (.A(n_2241),
    .Y(n_2239));
 INVxp33_ASAP7_75t_R g52863 (.A(n_2237),
    .Y(n_2238));
 INVxp33_ASAP7_75t_R g52866 (.A(n_2236),
    .Y(n_1826));
 HB1xp67_ASAP7_75t_R g52870 (.A(n_2237),
    .Y(n_2236));
 INVxp33_ASAP7_75t_R g52873 (.A(n_2234),
    .Y(n_1825));
 HB1xp67_ASAP7_75t_R g52874 (.A(n_2235),
    .Y(n_2234));
 OR3x1_ASAP7_75t_R g52884__6131 (.A(n_2210),
    .B(n_3411),
    .C(n_3440),
    .Y(n_2232));
 OR5x1_ASAP7_75t_R g52886__1881 (.A(n_2181),
    .B(n_14152),
    .C(n_14154),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .E(n_14134),
    .Y(n_2231));
 OAI22xp33_ASAP7_75t_R g52887__5115 (.A1(n_2201),
    .A2(n_2101),
    .B1(n_2136),
    .B2(n_2186),
    .Y(n_2230));
 NOR2xp33_ASAP7_75t_R g52888__7482 (.A(n_2202),
    .B(n_2217),
    .Y(n_2244));
 AOI21xp33_ASAP7_75t_R g52889__4733 (.A1(n_3824),
    .A2(n_13920),
    .B(n_2213),
    .Y(n_2241));
 NAND2xp33_ASAP7_75t_R g52890__6161 (.A(n_2202),
    .B(n_2218),
    .Y(n_2237));
 NOR2xp33_ASAP7_75t_R g52891__9315 (.A(n_2202),
    .B(n_2218),
    .Y(n_2235));
 NAND2xp33_ASAP7_75t_R g52892__9945 (.A(n_2202),
    .B(n_2217),
    .Y(n_2233));
 AOI22xp33_ASAP7_75t_R g52893__2883 (.A1(n_1844),
    .A2(n_2208),
    .B1(n_3597),
    .B2(n_3749),
    .Y(n_2225));
 NAND5xp2_ASAP7_75t_R g52894__2346 (.A(n_2191),
    .B(n_2147),
    .C(n_2153),
    .D(n_2146),
    .E(n_2081),
    .Y(n_2224));
 A2O1A1Ixp33_ASAP7_75t_R g52895__1666 (.A1(n_2001),
    .A2(n_2192),
    .B(n_2024),
    .C(n_2123),
    .Y(n_2223));
 AOI22xp33_ASAP7_75t_R g52896__7410 (.A1(n_1844),
    .A2(n_2200),
    .B1(n_3597),
    .B2(n_3748),
    .Y(n_2222));
 AOI221xp5_ASAP7_75t_R g52897__6417 (.A1(n_3595),
    .A2(n_3598),
    .B1(n_3743),
    .B2(n_3597),
    .C(n_2215),
    .Y(n_2221));
 AOI221xp5_ASAP7_75t_R g52898__5477 (.A1(u4_exp_div[2]),
    .A2(n_1844),
    .B1(n_3745),
    .B2(n_3597),
    .C(n_2127),
    .Y(n_2220));
 MAJIxp5_ASAP7_75t_R g52899__2398 (.A(n_2204),
    .B(div_opa_ldz_r2[4]),
    .C(exp_r[4]),
    .Y(n_2229));
 AOI22xp33_ASAP7_75t_R g52900__5107 (.A1(fract_denorm[46]),
    .A2(n_2202),
    .B1(fract_denorm[47]),
    .B2(n_2203),
    .Y(n_2228));
 AOI22xp33_ASAP7_75t_R g52901__6260 (.A1(fract_denorm[25]),
    .A2(n_2202),
    .B1(fract_denorm[26]),
    .B2(n_2203),
    .Y(n_2227));
 AOI22xp33_ASAP7_75t_R g52902__4319 (.A1(fract_denorm[26]),
    .A2(n_2202),
    .B1(fract_denorm[27]),
    .B2(n_2203),
    .Y(n_2226));
 INVxp33_ASAP7_75t_R g52903 (.A(inf_mul),
    .Y(n_2219));
 INVxp33_ASAP7_75t_R g52904 (.A(n_2218),
    .Y(n_2217));
 NAND2xp33_ASAP7_75t_R g52909__8428 (.A(n_1977),
    .B(n_2205),
    .Y(n_2216));
 OAI221xp5_ASAP7_75t_R g52910__5526 (.A1(n_2136),
    .A2(n_2116),
    .B1(n_2114),
    .B2(n_2101),
    .C(n_2187),
    .Y(n_2218));
 OAI22xp33_ASAP7_75t_R g52911__6783 (.A1(n_2188),
    .A2(u4_exp_zero),
    .B1(n_13919),
    .B2(n_2129),
    .Y(n_2215));
 OR5x1_ASAP7_75t_R g52912__3680 (.A(n_2196),
    .B(remainder[16]),
    .C(remainder[17]),
    .D(remainder[22]),
    .E(remainder[23]),
    .Y(n_2214));
 OAI221xp5_ASAP7_75t_R g52913__1617 (.A1(n_2149),
    .A2(n_2059),
    .B1(n_2136),
    .B2(n_2142),
    .C(n_2190),
    .Y(n_2213));
 OAI22xp33_ASAP7_75t_R g52914__2802 (.A1(n_2189),
    .A2(u4_exp_zero),
    .B1(n_13920),
    .B2(n_2177),
    .Y(n_2212));
 O2A1O1Ixp33_ASAP7_75t_R g52915__1705 (.A1(n_2003),
    .A2(n_2170),
    .B(n_2137),
    .C(n_1998),
    .Y(n_2211));
 OAI21xp33_ASAP7_75t_R g52916__5122 (.A1(n_3527),
    .A2(n_2150),
    .B(n_2197),
    .Y(u4_exp_div[3]));
 AOI32xp33_ASAP7_75t_R g52917__8246 (.A1(n_2156),
    .A2(rmode_r2[0]),
    .A3(rmode_r2[1]),
    .B1(n_2121),
    .B2(u1_signa_r),
    .Y(n_2209));
 OAI21xp33_ASAP7_75t_R g52919__7098 (.A1(n_3529),
    .A2(n_2111),
    .B(n_2185),
    .Y(n_2208));
 A2O1A1Ixp33_ASAP7_75t_R g52920__6131 (.A1(n_3580),
    .A2(n_2163),
    .B(n_1952),
    .C(n_1977),
    .Y(n_2207));
 NAND3xp33_ASAP7_75t_R g52922__1881 (.A(n_620),
    .B(n_2193),
    .C(fpu_op_r2[0]),
    .Y(n_2206));
 OR5x1_ASAP7_75t_R g52923__5115 (.A(n_2131),
    .B(n_3415),
    .C(n_3472),
    .D(n_3456),
    .E(n_3454),
    .Y(n_2210));
 OAI221xp5_ASAP7_75t_R g52924__7482 (.A1(n_2073),
    .A2(n_3529),
    .B1(n_2118),
    .B2(n_3528),
    .C(n_2167),
    .Y(u4_exp_div[4]));
 INVxp33_ASAP7_75t_R g52925 (.A(n_2205),
    .Y(n_2204));
 INVxp33_ASAP7_75t_R g52926 (.A(n_2203),
    .Y(n_2202));
 XOR2xp5_ASAP7_75t_R g52927__4733 (.A(n_1974),
    .B(n_2175),
    .Y(n_2201));
 OAI221xp5_ASAP7_75t_R g52928__6161 (.A1(n_2143),
    .A2(n_3528),
    .B1(n_2108),
    .B2(n_3529),
    .C(n_2184),
    .Y(n_2200));
 AOI31xp33_ASAP7_75t_R g52929__9315 (.A1(n_2164),
    .A2(u2_n_710),
    .A3(u2_n_606),
    .B(n_2074),
    .Y(n_2199));
 AOI22xp33_ASAP7_75t_R g52930__9945 (.A1(u0_qnan_r_a),
    .A2(u0_expa_ff),
    .B1(u0_qnan_r_b),
    .B2(u0_expb_ff),
    .Y(n_2198));
 AOI211xp5_ASAP7_75t_R g52931__2883 (.A1(n_1863),
    .A2(n_3737),
    .B(n_2159),
    .C(n_2174),
    .Y(n_2197));
 OR5x1_ASAP7_75t_R g52932__2346 (.A(n_2183),
    .B(remainder[20]),
    .C(remainder[19]),
    .D(remainder[21]),
    .E(remainder[18]),
    .Y(n_2196));
 MAJIxp5_ASAP7_75t_R g52933__1666 (.A(n_2176),
    .B(div_opa_ldz_r2[3]),
    .C(exp_r[3]),
    .Y(n_2205));
 OAI221xp5_ASAP7_75t_R g52934__7410 (.A1(n_2149),
    .A2(u4_sll_315_50_n_29),
    .B1(n_13972),
    .B2(n_1844),
    .C(n_2179),
    .Y(n_2203));
 INVxp33_ASAP7_75t_R g52935 (.A(underflow_fmul_d[0]),
    .Y(n_2195));
 INVxp33_ASAP7_75t_R g52936 (.A(opa_nan),
    .Y(n_2193));
 OAI221xp5_ASAP7_75t_R g52938__6417 (.A1(n_2122),
    .A2(n_2075),
    .B1(n_1986),
    .B2(n_1991),
    .C(n_2026),
    .Y(n_2192));
 NOR5xp2_ASAP7_75t_R g52939__5477 (.A(n_2160),
    .B(n_2144),
    .C(n_2145),
    .D(n_2109),
    .E(n_2122),
    .Y(n_2191));
 A2O1A1Ixp33_ASAP7_75t_R g52940__2398 (.A1(n_2120),
    .A2(n_1976),
    .B(n_2157),
    .C(n_2102),
    .Y(n_2190));
 NAND2xp33_ASAP7_75t_R g52941__5107 (.A(u0_infa_f_r),
    .B(u0_expa_ff),
    .Y(n_2194));
 AOI32xp33_ASAP7_75t_R g52943__6260 (.A1(n_2134),
    .A2(n_3599),
    .A3(fract_denorm[47]),
    .B1(n_2161),
    .B2(n_3808),
    .Y(n_2189));
 AOI31xp33_ASAP7_75t_R g52944__4319 (.A1(n_2134),
    .A2(n_3599),
    .A3(fract_denorm[46]),
    .B(n_2180),
    .Y(n_2188));
 AOI22xp33_ASAP7_75t_R g52945__8428 (.A1(n_2148),
    .A2(n_716),
    .B1(n_3820),
    .B2(n_13920),
    .Y(n_2187));
 XOR2xp5_ASAP7_75t_R g52946__5526 (.A(n_2163),
    .B(n_1974),
    .Y(n_2186));
 AOI221xp5_ASAP7_75t_R g52947__6783 (.A1(n_1863),
    .A2(n_3731),
    .B1(n_3809),
    .B2(n_1024),
    .C(n_2158),
    .Y(n_2185));
 AOI22xp33_ASAP7_75t_R g52948__3680 (.A1(n_1024),
    .A2(n_3814),
    .B1(n_3733),
    .B2(n_1863),
    .Y(n_2184));
 OAI221xp5_ASAP7_75t_R g52949__1617 (.A1(n_2115),
    .A2(n_3528),
    .B1(n_2069),
    .B2(n_3529),
    .C(n_2067),
    .Y(u4_exp_div[2]));
 OR5x1_ASAP7_75t_R g52950__2802 (.A(n_2141),
    .B(remainder[0]),
    .C(remainder[1]),
    .D(remainder[2]),
    .E(remainder[3]),
    .Y(n_2183));
 OR3x1_ASAP7_75t_R g52951__1705 (.A(n_2164),
    .B(n_2056),
    .C(u2_n_775),
    .Y(n_2182));
 OR4x1_ASAP7_75t_R g52952__5122 (.A(n_2072),
    .B(n_14124),
    .C(n_14142),
    .D(n_14140),
    .Y(n_2181));
 NOR2xp33_ASAP7_75t_R g52953__8246 (.A(n_3727),
    .B(n_2162),
    .Y(n_2180));
 OAI21xp33_ASAP7_75t_R g52955__7098 (.A1(n_2102),
    .A2(n_2135),
    .B(n_3717),
    .Y(n_2179));
 OAI31xp33_ASAP7_75t_R g52956__6131 (.A1(u0_n_321),
    .A2(n_3544),
    .A3(n_2079),
    .B(n_2152),
    .Y(n_2178));
 INVxp33_ASAP7_75t_R g52959 (.A(n_2177),
    .Y(u4_exp_div[1]));
 INVxp33_ASAP7_75t_R g52960 (.A(n_2175),
    .Y(n_2176));
 O2A1O1Ixp33_ASAP7_75t_R g52961__1881 (.A1(n_1993),
    .A2(n_2080),
    .B(n_2130),
    .C(n_3528),
    .Y(n_2174));
 O2A1O1Ixp33_ASAP7_75t_R g52962__5115 (.A1(exp_r[4]),
    .A2(n_3715),
    .B(n_1971),
    .C(n_2149),
    .Y(n_2173));
 OR5x1_ASAP7_75t_R g52964__4733 (.A(u4_n_1819),
    .B(u4_n_1820),
    .C(u4_n_1818),
    .D(u4_n_1827),
    .E(n_2062),
    .Y(n_2171));
 OAI22xp33_ASAP7_75t_R g52965__6161 (.A1(n_2117),
    .A2(n_2077),
    .B1(n_2017),
    .B2(n_2014),
    .Y(n_2170));
 OAI22xp33_ASAP7_75t_R g52966__9315 (.A1(n_2112),
    .A2(n_2090),
    .B1(n_2081),
    .B2(n_1995),
    .Y(n_2169));
 AND5x1_ASAP7_75t_R g52967__9945 (.A(u4_n_1834),
    .B(u4_n_1833),
    .C(n_2125),
    .D(u4_n_1836),
    .E(u4_n_1835),
    .Y(n_2168));
 AOI22xp33_ASAP7_75t_R g52968__2883 (.A1(n_1024),
    .A2(n_3813),
    .B1(n_3732),
    .B2(n_1863),
    .Y(n_2167));
 AOI221xp5_ASAP7_75t_R g52969__2346 (.A1(n_3808),
    .A2(n_1024),
    .B1(n_3730),
    .B2(n_1919),
    .C(n_2154),
    .Y(n_2177));
 MAJIxp5_ASAP7_75t_R g52970__1666 (.A(n_2119),
    .B(div_opa_ldz_r2[2]),
    .C(exp_r[2]),
    .Y(n_2175));
 INVxp33_ASAP7_75t_R g52971 (.A(n_2165),
    .Y(n_2166));
 INVxp33_ASAP7_75t_R g52972 (.A(n_2162),
    .Y(n_2161));
 NAND2xp33_ASAP7_75t_R g52973__7410 (.A(n_2123),
    .B(n_2137),
    .Y(n_2160));
 O2A1O1Ixp33_ASAP7_75t_R g52974__6417 (.A1(n_1985),
    .A2(n_3761),
    .B(n_2095),
    .C(n_3529),
    .Y(n_2159));
 O2A1O1Ixp33_ASAP7_75t_R g52975__5477 (.A1(n_1992),
    .A2(n_2023),
    .B(n_2093),
    .C(n_3528),
    .Y(n_2158));
 NOR2xp33_ASAP7_75t_R g52976__2398 (.A(n_2120),
    .B(n_1976),
    .Y(n_2157));
 OR2x2_ASAP7_75t_R g52977__5107 (.A(u1_signa_r),
    .B(n_2121),
    .Y(n_2156));
 NOR3xp33_ASAP7_75t_R g52978__6260 (.A(u4_f2i_zero),
    .B(n_2058),
    .C(n_2068),
    .Y(n_2155));
 OAI21xp33_ASAP7_75t_R g52980__4319 (.A1(n_3531),
    .A2(n_3730),
    .B(n_2132),
    .Y(n_2154));
 NAND5xp2_ASAP7_75t_R g52981__8428 (.A(n_2063),
    .B(opb_r[30]),
    .C(opb_r[23]),
    .D(opb_r[27]),
    .E(opb_r[26]),
    .Y(n_2165));
 NAND2xp33_ASAP7_75t_R g52982__5526 (.A(n_2139),
    .B(n_1896),
    .Y(n_2164));
 OAI21xp33_ASAP7_75t_R g52983__6783 (.A1(n_1139),
    .A2(n_2076),
    .B(n_3563),
    .Y(n_2163));
 NAND2xp33_ASAP7_75t_R g52984__3680 (.A(n_3599),
    .B(n_3494),
    .Y(n_2162));
 INVxp33_ASAP7_75t_R g52985 (.A(n_2151),
    .Y(n_2152));
 INVxp33_ASAP7_75t_R g52986 (.A(n_2150),
    .Y(n_3806));
 INVxp33_ASAP7_75t_R g52987 (.A(n_2149),
    .Y(n_2148));
 NOR5xp2_ASAP7_75t_R g52988__1617 (.A(n_2138),
    .B(n_2019),
    .C(n_2007),
    .D(n_2003),
    .E(n_2002),
    .Y(n_2147));
 AND5x1_ASAP7_75t_R g52989__2802 (.A(n_2086),
    .B(n_2084),
    .C(n_2082),
    .D(n_1989),
    .E(n_2017),
    .Y(n_2146));
 NAND4xp25_ASAP7_75t_R g52990__1705 (.A(n_1997),
    .B(n_2001),
    .C(n_2016),
    .D(n_2027),
    .Y(n_2145));
 NAND4xp25_ASAP7_75t_R g52991__5122 (.A(n_2107),
    .B(n_2026),
    .C(n_2000),
    .D(n_1991),
    .Y(n_2144));
 NOR3xp33_ASAP7_75t_R g52992__8246 (.A(u4_exp_zero),
    .B(n_2134),
    .C(n_1955),
    .Y(u4_n_1266));
 XNOR2xp5_ASAP7_75t_R g52993__7098 (.A(n_2053),
    .B(n_1963),
    .Y(n_2143));
 XNOR2xp5_ASAP7_75t_R g52994__6131 (.A(n_1976),
    .B(n_2076),
    .Y(n_2142));
 OR4x1_ASAP7_75t_R g52995__1881 (.A(remainder[7]),
    .B(remainder[4]),
    .C(remainder[6]),
    .D(remainder[5]),
    .Y(n_2141));
 XOR2xp5_ASAP7_75t_R g52996__5115 (.A(n_2054),
    .B(n_1962),
    .Y(n_3814));
 AOI211xp5_ASAP7_75t_R g52997__7482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .A2(n_1933),
    .B(n_2090),
    .C(n_2021),
    .Y(n_2153));
 NAND5xp2_ASAP7_75t_R g52998__4733 (.A(n_2060),
    .B(opa_r[30]),
    .C(opa_r[28]),
    .D(opa_r[27]),
    .E(opa_r[26]),
    .Y(n_2151));
 XNOR2xp5_ASAP7_75t_R g52999__6161 (.A(n_2055),
    .B(n_1966),
    .Y(n_2150));
 NAND3xp33_ASAP7_75t_R g53000__9315 (.A(n_2078),
    .B(n_1844),
    .C(n_1983),
    .Y(n_2149));
 INVxp33_ASAP7_75t_R g53001 (.A(n_2124),
    .Y(n_3513));
 INVxp33_ASAP7_75t_R g53002 (.A(n_2135),
    .Y(n_2136));
 INVxp33_ASAP7_75t_R g53003 (.A(n_2134),
    .Y(n_3494));
 NAND5xp2_ASAP7_75t_R g53004__9945 (.A(n_2061),
    .B(exp_mul[3]),
    .C(exp_mul[2]),
    .D(exp_mul[0]),
    .E(exp_mul[1]),
    .Y(n_2133));
 AO21x1_ASAP7_75t_R g53006__2883 (.A1(n_3521),
    .A2(n_3807),
    .B(n_3529),
    .Y(n_2132));
 OR4x1_ASAP7_75t_R g53007__2346 (.A(n_3452),
    .B(n_3444),
    .C(n_3474),
    .D(n_3401),
    .Y(n_2131));
 NAND2xp33_ASAP7_75t_R g53008__1666 (.A(n_1993),
    .B(n_2080),
    .Y(n_2130));
 O2A1O1Ixp33_ASAP7_75t_R g53009__7410 (.A1(n_1919),
    .A2(n_1863),
    .B(n_3740),
    .C(n_2070),
    .Y(n_2129));
 AOI21xp33_ASAP7_75t_R g53010__6417 (.A1(n_3568),
    .A2(n_1969),
    .B(n_1865),
    .Y(n_2128));
 O2A1O1Ixp33_ASAP7_75t_R g53011__5477 (.A1(n_1685),
    .A2(n_3480),
    .B(n_3565),
    .C(n_1865),
    .Y(n_2127));
 OR5x1_ASAP7_75t_R g53012__2398 (.A(n_3505),
    .B(n_2071),
    .C(u4_n_1944),
    .D(u4_n_1942),
    .E(u4_n_1934),
    .Y(n_2126));
 AND5x1_ASAP7_75t_R g53014__5107 (.A(n_2066),
    .B(u4_n_1844),
    .C(u4_n_1843),
    .D(u4_n_1846),
    .E(u4_n_1845),
    .Y(n_2125));
 AND2x2_ASAP7_75t_R g53015__6260 (.A(n_26),
    .B(n_2078),
    .Y(n_2140));
 NAND5xp2_ASAP7_75t_R g53016__4319 (.A(u2_exp_tmp1[6]),
    .B(n_1957),
    .C(n_14295),
    .D(n_1990),
    .E(u2_exp_tmp1[2]),
    .Y(n_2139));
 O2A1O1Ixp33_ASAP7_75t_R g53017__8428 (.A1(opas_r2),
    .A2(n_3754),
    .B(n_3512),
    .C(n_3803),
    .Y(n_2124));
 AO21x1_ASAP7_75t_R g53018__5526 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .A2(n_1875),
    .B(n_2088),
    .Y(n_2138));
 AOI21xp33_ASAP7_75t_R g53019__6783 (.A1(n_14160),
    .A2(n_1884),
    .B(n_2083),
    .Y(n_2137));
 NOR2xp33_ASAP7_75t_R g53020__3680 (.A(n_1982),
    .B(n_2078),
    .Y(n_2135));
 O2A1O1Ixp33_ASAP7_75t_R g53021__1617 (.A1(fract_denorm[47]),
    .A2(n_1801),
    .B(n_3502),
    .C(n_3801),
    .Y(n_2134));
 INVxp33_ASAP7_75t_R g53022 (.A(n_2120),
    .Y(n_2119));
 XOR2xp5_ASAP7_75t_R g53023__2802 (.A(n_3585),
    .B(n_1965),
    .Y(n_2118));
 OA21x2_ASAP7_75t_R g53024__1705 (.A1(n_1989),
    .A2(n_2006),
    .B(n_2005),
    .Y(n_2117));
 XOR2xp5_ASAP7_75t_R g53025__5122 (.A(n_1975),
    .B(n_3576),
    .Y(n_2116));
 XOR2xp5_ASAP7_75t_R g53026__8246 (.A(n_3590),
    .B(n_1967),
    .Y(n_2115));
 XOR2xp5_ASAP7_75t_R g53027__7098 (.A(n_1975),
    .B(n_1980),
    .Y(n_2114));
 XNOR2xp5_ASAP7_75t_R g53028__6131 (.A(n_1976),
    .B(n_3719),
    .Y(n_2113));
 AOI21xp33_ASAP7_75t_R g53029__1881 (.A1(n_2019),
    .A2(n_2022),
    .B(n_2020),
    .Y(n_2112));
 OAI32xp33_ASAP7_75t_R g53030__5115 (.A1(n_1945),
    .A2(n_3729),
    .A3(n_3728),
    .B1(n_3764),
    .B2(n_1961),
    .Y(n_2111));
 XNOR2xp5_ASAP7_75t_R g53031__7482 (.A(n_3718),
    .B(n_1977),
    .Y(n_2110));
 OAI21xp33_ASAP7_75t_R g53032__4733 (.A1(n_3303),
    .A2(u5_mul_69_18_n_54),
    .B(n_2100),
    .Y(n_2109));
 XNOR2xp5_ASAP7_75t_R g53033__6161 (.A(n_1984),
    .B(n_3763),
    .Y(n_2108));
 NOR4xp25_ASAP7_75t_R g53034__9315 (.A(n_2020),
    .B(n_2024),
    .C(n_2010),
    .D(n_2004),
    .Y(n_2107));
 AOI21xp33_ASAP7_75t_R g53035__9945 (.A1(n_1873),
    .A2(n_14130),
    .B(n_2085),
    .Y(n_2123));
 XNOR2xp5_ASAP7_75t_R g53036__2883 (.A(n_3817),
    .B(n_1964),
    .Y(n_3813));
 AO221x1_ASAP7_75t_R g53037__2346 (.A1(n_1944),
    .A2(n_14124),
    .B1(n_1877),
    .B2(n_14178),
    .C(n_1986),
    .Y(n_2122));
 XOR2xp5_ASAP7_75t_R g53038__1666 (.A(n_2011),
    .B(u1_add_r),
    .Y(n_2121));
 XNOR2xp5_ASAP7_75t_R g53039__7410 (.A(n_3571),
    .B(n_1960),
    .Y(n_3809));
 MAJIxp5_ASAP7_75t_R g53040__6417 (.A(n_1981),
    .B(div_opa_ldz_r2[1]),
    .C(exp_r[1]),
    .Y(n_2120));
 INVxp33_ASAP7_75t_R g53041 (.A(sign_exe),
    .Y(n_2106));
 INVxp33_ASAP7_75t_R g53042 (.A(n_2103),
    .Y(n_2104));
 INVxp33_ASAP7_75t_R g53043 (.A(n_2102),
    .Y(n_2101));
 NOR2xp33_ASAP7_75t_R g53044__5477 (.A(n_2015),
    .B(n_1996),
    .Y(n_2100));
 NAND2xp33_ASAP7_75t_R g53070__2398 (.A(exp_ovf_r[0]),
    .B(n_1978),
    .Y(n_2099));
 NAND2xp33_ASAP7_75t_R g53071__5107 (.A(u0_fracta_00),
    .B(u0_expa_00),
    .Y(n_2098));
 NAND2xp33_ASAP7_75t_R g53072__6260 (.A(n_13946),
    .B(n_1988),
    .Y(n_2097));
 NAND2xp33_ASAP7_75t_R g53074__4319 (.A(n_1974),
    .B(n_3569),
    .Y(n_2096));
 NAND2xp33_ASAP7_75t_R g53075__8428 (.A(n_1985),
    .B(n_3761),
    .Y(n_2095));
 NAND2xp33_ASAP7_75t_R g53076__5526 (.A(n_3720),
    .B(n_1975),
    .Y(n_2094));
 NAND2xp33_ASAP7_75t_R g53077__6783 (.A(n_1992),
    .B(n_2023),
    .Y(n_2093));
 NAND2xp33_ASAP7_75t_R g53078__3680 (.A(n_2013),
    .B(n_36),
    .Y(n_2105));
 NOR2xp33_ASAP7_75t_R g53079__1617 (.A(exp_ovf_r[0]),
    .B(n_1979),
    .Y(n_2103));
 NOR2xp33_ASAP7_75t_R g53080__2802 (.A(n_26),
    .B(n_1979),
    .Y(n_2102));
 INVxp33_ASAP7_75t_R g53081 (.A(n_2091),
    .Y(n_2092));
 INVxp33_ASAP7_75t_R g53082 (.A(n_2086),
    .Y(n_2087));
 NOR2xp33_ASAP7_75t_R g53083__1705 (.A(n_2000),
    .B(n_2002),
    .Y(n_2075));
 NOR3xp33_ASAP7_75t_R g53084__5122 (.A(fractb_mul[23]),
    .B(n_13981),
    .C(opa_r[30]),
    .Y(n_2074));
 AOI21xp33_ASAP7_75t_R g53085__8246 (.A1(n_3728),
    .A2(n_3762),
    .B(n_1984),
    .Y(n_2073));
 OR3x1_ASAP7_75t_R g53086__7098 (.A(n_14150),
    .B(n_14148),
    .C(n_14178),
    .Y(n_2072));
 OR3x1_ASAP7_75t_R g53087__6131 (.A(u4_n_1938),
    .B(u4_n_1948),
    .C(u4_n_1946),
    .Y(n_2071));
 AOI22xp33_ASAP7_75t_R g53088__1881 (.A1(n_3527),
    .A2(n_1931),
    .B1(n_3529),
    .B2(n_3727),
    .Y(n_2070));
 OA21x2_ASAP7_75t_R g53089__5115 (.A1(n_3805),
    .A2(n_1949),
    .B(n_1985),
    .Y(n_2069));
 XOR2xp5_ASAP7_75t_R g53090__7482 (.A(n_3774),
    .B(n_792),
    .Y(n_2068));
 AOI22xp33_ASAP7_75t_R g53091__4733 (.A1(n_1024),
    .A2(n_3805),
    .B1(n_3736),
    .B2(n_1863),
    .Y(n_2067));
 AND4x1_ASAP7_75t_R g53092__6161 (.A(u4_n_1840),
    .B(u4_n_1839),
    .C(u4_n_1842),
    .D(u4_n_1841),
    .Y(n_2066));
 OR4x1_ASAP7_75t_R g53093__9315 (.A(u4_n_1826),
    .B(u4_n_1829),
    .C(u4_n_1828),
    .D(u4_n_1821),
    .Y(n_2065));
 AND4x1_ASAP7_75t_R g53094__9945 (.A(u4_n_1838),
    .B(u4_n_1837),
    .C(u4_n_1832),
    .D(u4_n_1831),
    .Y(n_2064));
 AND4x1_ASAP7_75t_R g53095__2883 (.A(opb_r[29]),
    .B(opb_r[25]),
    .C(opb_r[28]),
    .D(opb_r[24]),
    .Y(n_2063));
 OR4x1_ASAP7_75t_R g53096__2346 (.A(u4_n_1823),
    .B(u4_n_1822),
    .C(u4_n_1825),
    .D(u4_n_1824),
    .Y(n_2062));
 AND4x1_ASAP7_75t_R g53097__1666 (.A(exp_mul[7]),
    .B(exp_mul[6]),
    .C(exp_mul[5]),
    .D(exp_mul[4]),
    .Y(n_2061));
 AND4x1_ASAP7_75t_R g53098__7410 (.A(opa_r[25]),
    .B(opa_r[24]),
    .C(opa_r[29]),
    .D(opa_r[23]),
    .Y(n_2060));
 XOR2xp5_ASAP7_75t_R g53099__6417 (.A(n_716),
    .B(exp_r[2]),
    .Y(n_2059));
 XOR2xp5_ASAP7_75t_R g53100__5477 (.A(n_3500),
    .B(exp_r[7]),
    .Y(n_2058));
 XNOR2xp5_ASAP7_75t_R g53101__2398 (.A(n_3565),
    .B(n_98),
    .Y(n_2057));
 XNOR2xp5_ASAP7_75t_R g53102__5107 (.A(u2_n_710),
    .B(n_13981),
    .Y(n_2056));
 NOR3xp33_ASAP7_75t_R g53103__6260 (.A(fract_denorm[10]),
    .B(fract_denorm[9]),
    .C(fract_denorm[7]),
    .Y(n_2091));
 AO21x1_ASAP7_75t_R g53104__4319 (.A1(n_14148),
    .A2(n_1939),
    .B(n_1995),
    .Y(n_2090));
 NAND3xp33_ASAP7_75t_R g53105__8428 (.A(n_1950),
    .B(exp_r[3]),
    .C(exp_r[4]),
    .Y(n_2089));
 AO21x1_ASAP7_75t_R g53106__5526 (.A1(n_14140),
    .A2(u5_mul_69_18_n_106),
    .B(n_2009),
    .Y(n_2088));
 AOI21xp33_ASAP7_75t_R g53107__6783 (.A1(n_14152),
    .A2(n_1879),
    .B(n_2006),
    .Y(n_2086));
 AO21x1_ASAP7_75t_R g53108__3680 (.A1(n_14132),
    .A2(n_1930),
    .B(n_1999),
    .Y(n_2085));
 AOI21xp33_ASAP7_75t_R g53109__1617 (.A1(n_3818),
    .A2(n_3517),
    .B(n_1686),
    .Y(n_2055));
 AOI22xp33_ASAP7_75t_R g53110__2802 (.A1(n_3474),
    .A2(n_1937),
    .B1(n_3444),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .Y(n_2084));
 OAI22xp33_ASAP7_75t_R g53111__1705 (.A1(n_3444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B1(n_3386),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_584),
    .Y(n_2083));
 AOI22xp33_ASAP7_75t_R g53112__5122 (.A1(n_3432),
    .A2(n_1889),
    .B1(n_3468),
    .B2(u5_mul_69_18_n_125),
    .Y(n_2082));
 AOI22xp33_ASAP7_75t_R g53113__8246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .A2(n_3415),
    .B1(n_3454),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(n_2081));
 NAND2xp33_ASAP7_75t_R g53114__7098 (.A(n_3591),
    .B(n_1970),
    .Y(n_2080));
 AOI21xp33_ASAP7_75t_R g53115__6131 (.A1(n_3817),
    .A2(n_3509),
    .B(n_1891),
    .Y(n_2054));
 AOI21xp33_ASAP7_75t_R g53116__1881 (.A1(n_3585),
    .A2(n_3511),
    .B(n_1951),
    .Y(n_2053));
 NAND3xp33_ASAP7_75t_R g53117__5115 (.A(u5_mul_69_18_n_54),
    .B(n_1944),
    .C(n_1877),
    .Y(n_2079));
 OR3x1_ASAP7_75t_R g53118__7482 (.A(n_3592),
    .B(n_36),
    .C(n_1020),
    .Y(n_2078));
 AO21x1_ASAP7_75t_R g53119__4733 (.A1(n_14156),
    .A2(n_1940),
    .B(n_2014),
    .Y(n_2077));
 AOI21xp33_ASAP7_75t_R g53120__6161 (.A1(n_3584),
    .A2(n_3576),
    .B(n_1895),
    .Y(n_2076));
 INVxp33_ASAP7_75t_R g53130 (.A(fasu_op_r1),
    .Y(n_2043));
 INVxp33_ASAP7_75t_R g53146 (.A(n_2021),
    .Y(n_2022));
 INVxp33_ASAP7_75t_R g53148 (.A(n_2013),
    .Y(n_2012));
 INVxp33_ASAP7_75t_R g53149 (.A(u1_signb_r),
    .Y(n_2011));
 OR2x2_ASAP7_75t_R g53181 (.A(n_1930),
    .B(n_14132),
    .Y(n_2027));
 NAND2xp33_ASAP7_75t_R g53183 (.A(n_3411),
    .B(u5_mul_69_18_n_89),
    .Y(n_2026));
 OR2x2_ASAP7_75t_R g53184 (.A(n_1865),
    .B(n_3757),
    .Y(n_2025));
 NOR2xp33_ASAP7_75t_R g53185 (.A(n_14128),
    .B(n_1883),
    .Y(n_2024));
 NAND2xp33_ASAP7_75t_R g53186 (.A(n_3560),
    .B(n_14181),
    .Y(n_2023));
 NOR2xp33_ASAP7_75t_R g53187 (.A(n_3476),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .Y(n_2021));
 NOR2xp33_ASAP7_75t_R g53188 (.A(n_14146),
    .B(n_1932),
    .Y(n_2020));
 NOR2xp33_ASAP7_75t_R g53189 (.A(n_1933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .Y(n_2019));
 NAND2xp33_ASAP7_75t_R g53190 (.A(fpu_op_r2[1]),
    .B(n_727),
    .Y(n_3557));
 OR2x2_ASAP7_75t_R g53191 (.A(n_14156),
    .B(n_1940),
    .Y(n_2017));
 OR2x2_ASAP7_75t_R g53192 (.A(n_14130),
    .B(n_1873),
    .Y(n_2016));
 NOR2xp33_ASAP7_75t_R g53193 (.A(n_14136),
    .B(n_80),
    .Y(n_2015));
 NAND2xp33_ASAP7_75t_R g53194 (.A(n_3808),
    .B(n_1931),
    .Y(n_3807));
 NOR2xp33_ASAP7_75t_R g53195 (.A(n_3401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .Y(n_2014));
 NOR2xp33_ASAP7_75t_R g53196 (.A(n_682),
    .B(n_3801),
    .Y(n_2013));
 INVxp33_ASAP7_75t_R g53199 (.A(n_2007),
    .Y(n_2008));
 INVxp33_ASAP7_75t_R g53200 (.A(n_2004),
    .Y(n_2005));
 INVxp33_ASAP7_75t_R g53201 (.A(n_1997),
    .Y(n_1998));
 INVxp33_ASAP7_75t_R g53202 (.A(u2_n_1493),
    .Y(n_1990));
 INVxp33_ASAP7_75t_R g53204 (.A(n_1983),
    .Y(n_1982));
 INVxp33_ASAP7_75t_R g53205 (.A(n_1980),
    .Y(n_1981));
 INVxp33_ASAP7_75t_R g53206 (.A(n_1979),
    .Y(n_1978));
 NAND2xp33_ASAP7_75t_R g53208 (.A(opb_r[31]),
    .B(opa_r[31]),
    .Y(n_1972));
 NAND2xp33_ASAP7_75t_R g53209 (.A(n_3715),
    .B(exp_r[4]),
    .Y(n_1971));
 NAND2xp33_ASAP7_75t_R g53210 (.A(n_3518),
    .B(n_3590),
    .Y(n_1970));
 NAND2xp33_ASAP7_75t_R g53211 (.A(n_3516),
    .B(n_3758),
    .Y(n_1969));
 NOR2xp33_ASAP7_75t_R g53212 (.A(n_3773),
    .B(n_3772),
    .Y(n_1968));
 NOR2xp33_ASAP7_75t_R g53213 (.A(n_1934),
    .B(n_14134),
    .Y(n_2010));
 NOR2xp33_ASAP7_75t_R g53214 (.A(n_3468),
    .B(u5_mul_69_18_n_125),
    .Y(n_2009));
 NOR2xp33_ASAP7_75t_R g53215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B(n_1875),
    .Y(n_2007));
 NOR2xp33_ASAP7_75t_R g53216 (.A(u5_mul_69_18_n_130),
    .B(n_3456),
    .Y(n_2006));
 NOR2xp33_ASAP7_75t_R g53217 (.A(n_14154),
    .B(n_1942),
    .Y(n_2004));
 AND2x2_ASAP7_75t_R g53218 (.A(n_3401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .Y(n_2003));
 NOR2xp33_ASAP7_75t_R g53219 (.A(n_14124),
    .B(n_1944),
    .Y(n_2002));
 NAND2xp33_ASAP7_75t_R g53220 (.A(n_14128),
    .B(n_1883),
    .Y(n_2001));
 NAND2xp33_ASAP7_75t_R g53221 (.A(n_3303),
    .B(u5_mul_69_18_n_54),
    .Y(n_2000));
 NOR2xp33_ASAP7_75t_R g53222 (.A(n_3434),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .Y(n_1999));
 NAND2xp33_ASAP7_75t_R g53223 (.A(n_3386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_584),
    .Y(n_1997));
 NAND2xp33_ASAP7_75t_R g53224 (.A(n_3591),
    .B(n_3518),
    .Y(n_1967));
 NAND2xp33_ASAP7_75t_R g53225 (.A(n_3502),
    .B(n_26),
    .Y(u4_n_1091));
 AND2x2_ASAP7_75t_R g53226 (.A(n_14136),
    .B(n_80),
    .Y(n_1996));
 NAND2xp33_ASAP7_75t_R g53227 (.A(n_3821),
    .B(n_3519),
    .Y(n_1966));
 NOR2xp33_ASAP7_75t_R g53228 (.A(n_3454),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(n_1995));
 NAND2xp33_ASAP7_75t_R g53229 (.A(n_1567),
    .B(n_1925),
    .Y(n_1994));
 NAND2xp33_ASAP7_75t_R g53230 (.A(n_3589),
    .B(n_3520),
    .Y(n_1993));
 NAND2xp33_ASAP7_75t_R g53231 (.A(n_3526),
    .B(n_3586),
    .Y(n_1992));
 OR2x2_ASAP7_75t_R g53232 (.A(n_1877),
    .B(n_14178),
    .Y(n_1991));
 NAND2xp33_ASAP7_75t_R g53233 (.A(u2_exp_tmp1[0]),
    .B(u2_exp_tmp1[1]),
    .Y(u2_n_1493));
 OR2x2_ASAP7_75t_R g53234 (.A(n_1879),
    .B(n_14152),
    .Y(n_1989));
 NAND2xp33_ASAP7_75t_R g53235 (.A(n_3588),
    .B(n_3511),
    .Y(n_1965));
 NAND2xp33_ASAP7_75t_R g53236 (.A(n_3583),
    .B(n_3581),
    .Y(n_1988));
 NAND2xp33_ASAP7_75t_R g53237 (.A(n_3509),
    .B(n_3825),
    .Y(n_1964));
 NAND2xp33_ASAP7_75t_R g53238 (.A(n_3587),
    .B(n_3510),
    .Y(n_1963));
 NOR2xp33_ASAP7_75t_R g53240 (.A(n_3411),
    .B(u5_mul_69_18_n_89),
    .Y(n_1986));
 NAND2xp33_ASAP7_75t_R g53241 (.A(n_3815),
    .B(n_3574),
    .Y(n_1962));
 OR2x2_ASAP7_75t_R g53242 (.A(n_3572),
    .B(n_3755),
    .Y(n_3512));
 NAND2xp33_ASAP7_75t_R g53243 (.A(fractb_mul[23]),
    .B(n_13883),
    .Y(u2_n_775));
 NOR2xp33_ASAP7_75t_R g53244 (.A(n_3728),
    .B(n_3729),
    .Y(n_1961));
 NAND2xp33_ASAP7_75t_R g53245 (.A(n_3522),
    .B(n_3810),
    .Y(n_1960));
 NAND2xp33_ASAP7_75t_R g53246 (.A(n_3812),
    .B(n_3561),
    .Y(n_3571));
 NAND2xp33_ASAP7_75t_R g53247 (.A(n_3805),
    .B(n_1949),
    .Y(n_1985));
 NOR2xp33_ASAP7_75t_R g53248 (.A(n_3762),
    .B(n_3728),
    .Y(n_1984));
 NAND2xp33_ASAP7_75t_R g53249 (.A(exp_ovf_r[1]),
    .B(u4_op_dn),
    .Y(n_1983));
 NAND2xp33_ASAP7_75t_R g53250 (.A(div_opa_ldz_r2[0]),
    .B(n_13972),
    .Y(n_1980));
 NAND2xp33_ASAP7_75t_R g53251 (.A(u4_op_dn),
    .B(n_1844),
    .Y(n_1979));
 NAND2xp33_ASAP7_75t_R g53252 (.A(n_3507),
    .B(n_3583),
    .Y(n_1977));
 NAND2xp33_ASAP7_75t_R g53253 (.A(n_3582),
    .B(n_3563),
    .Y(n_1976));
 NAND2xp33_ASAP7_75t_R g53254 (.A(n_3584),
    .B(n_3575),
    .Y(n_1975));
 NAND2xp33_ASAP7_75t_R g53255 (.A(n_3506),
    .B(n_3580),
    .Y(n_1974));
 INVxp33_ASAP7_75t_R g53256 (.A(n_3775),
    .Y(n_1069));
 INVxp33_ASAP7_75t_R g53258 (.A(u2_n_1487),
    .Y(n_1957));
 INVxp33_ASAP7_75t_R g53259 (.A(sign_mul),
    .Y(n_1956));
 INVxp33_ASAP7_75t_R g53260 (.A(n_3765),
    .Y(n_1955));
 INVxp33_ASAP7_75t_R g53261 (.A(sign_fasu),
    .Y(n_1954));
 INVxp33_ASAP7_75t_R g53263 (.A(n_3506),
    .Y(n_1952));
 INVxp33_ASAP7_75t_R g53264 (.A(n_3588),
    .Y(n_1951));
 INVxp33_ASAP7_75t_R g53265 (.A(n_3716),
    .Y(n_1950));
 INVxp33_ASAP7_75t_R g53266 (.A(n_3521),
    .Y(n_1949));
 INVxp33_ASAP7_75t_R g53270 (.A(n_3764),
    .Y(n_1945));
 INVxp33_ASAP7_75t_R g53271 (.A(n_3436),
    .Y(n_1944));
 INVxp33_ASAP7_75t_R g53272 (.A(n_3763),
    .Y(n_1943));
 INVxp33_ASAP7_75t_R g53273 (.A(n_3456),
    .Y(n_1942));
 INVxp33_ASAP7_75t_R g53275 (.A(n_3472),
    .Y(n_1940));
 INVxp33_ASAP7_75t_R g53276 (.A(n_3415),
    .Y(n_1939));
 INVxp33_ASAP7_75t_R g53278 (.A(n_14160),
    .Y(n_1937));
 INVxp33_ASAP7_75t_R g53279 (.A(n_3761),
    .Y(n_1936));
 INVxp33_ASAP7_75t_R g53280 (.A(n_3762),
    .Y(n_1935));
 INVxp33_ASAP7_75t_R g53281 (.A(n_3434),
    .Y(n_1934));
 INVxp33_ASAP7_75t_R g53282 (.A(n_3466),
    .Y(n_1933));
 INVxp33_ASAP7_75t_R g53283 (.A(n_3476),
    .Y(n_1932));
 INVxp33_ASAP7_75t_R g53284 (.A(n_3727),
    .Y(n_1931));
 INVxp33_ASAP7_75t_R g53285 (.A(n_3409),
    .Y(n_1930));
 INVxp33_ASAP7_75t_R g53286 (.A(exp_r[0]),
    .Y(u4_sll_315_50_n_29));
 INVxp33_ASAP7_75t_R g53287 (.A(fract_denorm[5]),
    .Y(n_1567));
 INVxp33_ASAP7_75t_R g53290 (.A(fract_denorm[6]),
    .Y(n_1925));
 INVxp33_ASAP7_75t_R g53292 (.A(fract_denorm[12]),
    .Y(n_1923));
 INVxp33_ASAP7_75t_R g53293 (.A(fract_denorm[4]),
    .Y(n_1922));
 INVxp33_ASAP7_75t_R g53294 (.A(fract_denorm[41]),
    .Y(n_1578));
 INVxp33_ASAP7_75t_R g53295 (.A(fract_denorm[25]),
    .Y(n_1920));
 INVxp33_ASAP7_75t_R g53296 (.A(n_3528),
    .Y(n_1919));
 INVxp33_ASAP7_75t_R g53297 (.A(fract_denorm[45]),
    .Y(n_1918));
 INVxp33_ASAP7_75t_R g53298 (.A(fract_denorm[9]),
    .Y(n_1917));
 INVxp33_ASAP7_75t_R g53299 (.A(fract_denorm[33]),
    .Y(n_1916));
 INVxp33_ASAP7_75t_R g53300 (.A(fract_denorm[13]),
    .Y(n_1915));
 INVxp33_ASAP7_75t_R g53301 (.A(fract_denorm[34]),
    .Y(n_1914));
 INVxp33_ASAP7_75t_R g53302 (.A(fract_denorm[10]),
    .Y(n_1913));
 INVxp33_ASAP7_75t_R g53303 (.A(fract_denorm[30]),
    .Y(n_1912));
 INVxp33_ASAP7_75t_R g53304 (.A(fract_denorm[28]),
    .Y(n_1911));
 INVxp33_ASAP7_75t_R g53305 (.A(fract_denorm[39]),
    .Y(n_1910));
 INVxp33_ASAP7_75t_R g53306 (.A(fract_denorm[14]),
    .Y(n_1569));
 INVxp33_ASAP7_75t_R g53307 (.A(fract_denorm[32]),
    .Y(n_1590));
 INVxp33_ASAP7_75t_R g53308 (.A(fract_denorm[29]),
    .Y(n_1588));
 INVxp33_ASAP7_75t_R g53309 (.A(fract_denorm[23]),
    .Y(n_1577));
 INVxp33_ASAP7_75t_R g53310 (.A(fract_denorm[17]),
    .Y(n_1585));
 INVxp33_ASAP7_75t_R g53311 (.A(fract_denorm[20]),
    .Y(n_1591));
 INVxp33_ASAP7_75t_R g53312 (.A(fract_denorm[16]),
    .Y(n_1903));
 INVxp33_ASAP7_75t_R g53313 (.A(fract_denorm[38]),
    .Y(n_1587));
 INVxp33_ASAP7_75t_R g53314 (.A(fract_denorm[35]),
    .Y(n_1576));
 INVxp33_ASAP7_75t_R g53315 (.A(fract_denorm[37]),
    .Y(n_1900));
 INVxp33_ASAP7_75t_R g53319 (.A(u2_exp_tmp1[7]),
    .Y(n_1896));
 INVxp33_ASAP7_75t_R g53320 (.A(n_3575),
    .Y(n_1895));
 INVxp33_ASAP7_75t_R g53322 (.A(opa_r[31]),
    .Y(n_725));
 INVxp33_ASAP7_75t_R g53323 (.A(opb_r[31]),
    .Y(n_728));
 INVxp33_ASAP7_75t_R g53324 (.A(n_3825),
    .Y(n_1891));
 INVxp33_ASAP7_75t_R g53325 (.A(n_3515),
    .Y(n_1685));
 INVxp33_ASAP7_75t_R g53326 (.A(n_14140),
    .Y(n_1889));
 INVxp33_ASAP7_75t_R g53331 (.A(n_3474),
    .Y(n_1884));
 INVxp33_ASAP7_75t_R g53332 (.A(n_3440),
    .Y(n_1883));
 INVxp33_ASAP7_75t_R g53336 (.A(n_3452),
    .Y(n_1879));
 INVxp33_ASAP7_75t_R g53337 (.A(n_3593),
    .Y(n_98));
 INVxp33_ASAP7_75t_R g53338 (.A(n_3427),
    .Y(n_1877));
 INVxp33_ASAP7_75t_R g53340 (.A(n_3438),
    .Y(n_1875));
 INVxp33_ASAP7_75t_R g53342 (.A(n_3395),
    .Y(n_1873));
 INVxp33_ASAP7_75t_R g53344 (.A(fract_denorm[3]),
    .Y(n_1871));
 INVxp33_ASAP7_75t_R g53346 (.A(n_3386),
    .Y(n_802));
 INVxp33_ASAP7_75t_R g53347 (.A(n_14164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_584));
 INVxp33_ASAP7_75t_R g53348 (.A(fract_denorm[7]),
    .Y(n_1867));
 INVxp33_ASAP7_75t_R g53349 (.A(fract_denorm[42]),
    .Y(n_1866));
 INVxp33_ASAP7_75t_R g53350 (.A(n_3598),
    .Y(n_1865));
 INVxp33_ASAP7_75t_R g53351 (.A(exp_r[1]),
    .Y(n_716));
 INVxp33_ASAP7_75t_R g53352 (.A(n_3531),
    .Y(n_1863));
 INVxp33_ASAP7_75t_R g53353 (.A(n_3803),
    .Y(n_1019));
 INVxp33_ASAP7_75t_R g53354 (.A(fract_denorm[43]),
    .Y(n_1861));
 INVxp33_ASAP7_75t_R g53355 (.A(fract_denorm[27]),
    .Y(n_1860));
 INVxp33_ASAP7_75t_R g53359 (.A(fract_denorm[8]),
    .Y(n_1568));
 INVxp33_ASAP7_75t_R g53360 (.A(fract_denorm[19]),
    .Y(n_1855));
 INVxp33_ASAP7_75t_R g53361 (.A(n_13946),
    .Y(n_1854));
 INVxp33_ASAP7_75t_R g53362 (.A(fract_denorm[18]),
    .Y(n_1853));
 INVxp33_ASAP7_75t_R g53363 (.A(fract_denorm[40]),
    .Y(n_1852));
 INVxp33_ASAP7_75t_R g53364 (.A(fract_denorm[31]),
    .Y(n_1851));
 INVxp33_ASAP7_75t_R g53365 (.A(fract_denorm[24]),
    .Y(n_1850));
 INVxp33_ASAP7_75t_R g53366 (.A(fract_denorm[15]),
    .Y(n_1849));
 INVxp33_ASAP7_75t_R g53368 (.A(fract_denorm[21]),
    .Y(n_1847));
 INVxp33_ASAP7_75t_R g53369 (.A(fract_denorm[22]),
    .Y(n_1846));
 INVxp33_ASAP7_75t_R g53370 (.A(fract_denorm[36]),
    .Y(n_1845));
 INVxp33_ASAP7_75t_R g53371 (.A(n_13919),
    .Y(n_1844));
 AO222x2_ASAP7_75t_R g53503 (.A1(n_680),
    .A2(fract_i2f[17]),
    .B1(n_677),
    .B2(quo[19]),
    .C1(n_671),
    .C2(prod[17]),
    .Y(n_651));
 INVxp33_ASAP7_75t_R g92 (.A(n_14055),
    .Y(n_14056));
 INVxp33_ASAP7_75t_R g94 (.A(u6_remainder[1]),
    .Y(n_14057));
 INVxp33_ASAP7_75t_R g96 (.A(u6_remainder[3]),
    .Y(n_14059));
 INVxp33_ASAP7_75t_R g98 (.A(u6_remainder[7]),
    .Y(n_14063));
 XOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g2 (.A(inc_u4_add_230_34_n_221),
    .B(u4_fract_out[13]),
    .Y(n_3790));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g291 (.A1(inc_u4_add_230_34_n_185),
    .A2(inc_u4_add_230_34_n_272),
    .B(u4_fract_out_pl1[23]),
    .Y(n_3799));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g292 (.A(inc_u4_add_230_34_n_272),
    .B(inc_u4_add_230_34_n_185),
    .Y(u4_fract_out_pl1[23]));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g293 (.A1(u4_fract_out[21]),
    .A2(inc_u4_add_230_34_n_189),
    .B(inc_u4_add_230_34_n_185),
    .Y(n_3798));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g294 (.A(u4_fract_out[21]),
    .B(inc_u4_add_230_34_n_189),
    .Y(inc_u4_add_230_34_n_185));
 XNOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g295 (.A(inc_u4_add_230_34_n_192),
    .B(u4_fract_out[20]),
    .Y(n_3797));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g296 (.A(inc_u4_add_230_34_n_278),
    .B(inc_u4_add_230_34_n_192),
    .Y(inc_u4_add_230_34_n_189));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g297 (.A1(u4_fract_out[19]),
    .A2(inc_u4_add_230_34_n_196),
    .B(inc_u4_add_230_34_n_192),
    .Y(n_3796));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g298 (.A(u4_fract_out[19]),
    .B(inc_u4_add_230_34_n_196),
    .Y(inc_u4_add_230_34_n_192));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g299 (.A1(inc_u4_add_230_34_n_200),
    .A2(inc_u4_add_230_34_n_270),
    .B(inc_u4_add_230_34_n_196),
    .Y(n_3795));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g300 (.A(inc_u4_add_230_34_n_270),
    .B(inc_u4_add_230_34_n_200),
    .Y(inc_u4_add_230_34_n_196));
 XNOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g301 (.A(inc_u4_add_230_34_n_204),
    .B(u4_fract_out[17]),
    .Y(n_3794));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g302 (.A(inc_u4_add_230_34_n_203),
    .B(u4_fract_out[17]),
    .Y(inc_u4_add_230_34_n_200));
 XNOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g303 (.A(inc_u4_add_230_34_n_208),
    .B(u4_fract_out[16]),
    .Y(n_3793));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g304 (.A(inc_u4_add_230_34_n_204),
    .Y(inc_u4_add_230_34_n_203));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g305 (.A(u4_fract_out[16]),
    .B(inc_u4_add_230_34_n_209),
    .Y(inc_u4_add_230_34_n_204));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g306 (.A1(u4_fract_out[15]),
    .A2(inc_u4_add_230_34_n_213),
    .B(inc_u4_add_230_34_n_208),
    .Y(n_3792));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g307 (.A(inc_u4_add_230_34_n_208),
    .Y(inc_u4_add_230_34_n_209));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g308 (.A(u4_fract_out[15]),
    .B(inc_u4_add_230_34_n_213),
    .Y(inc_u4_add_230_34_n_208));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g309 (.A1(inc_u4_add_230_34_n_217),
    .A2(inc_u4_add_230_34_n_277),
    .B(inc_u4_add_230_34_n_213),
    .Y(n_3791));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g310 (.A(inc_u4_add_230_34_n_277),
    .B(inc_u4_add_230_34_n_217),
    .Y(inc_u4_add_230_34_n_213));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g312 (.A(u4_fract_out[13]),
    .B(inc_u4_add_230_34_n_221),
    .Y(inc_u4_add_230_34_n_217));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g313 (.A1(inc_u4_add_230_34_n_226),
    .A2(inc_u4_add_230_34_n_284),
    .B(inc_u4_add_230_34_n_221),
    .Y(n_3789));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g315 (.A(inc_u4_add_230_34_n_284),
    .B(inc_u4_add_230_34_n_226),
    .Y(inc_u4_add_230_34_n_221));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g317 (.A(u4_fract_out[11]),
    .B(inc_u4_add_230_34_n_230),
    .Y(inc_u4_add_230_34_n_226));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g318 (.A1(inc_u4_add_230_34_n_235),
    .A2(inc_u4_add_230_34_n_286),
    .B(inc_u4_add_230_34_n_230),
    .Y(n_3787));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g320 (.A(inc_u4_add_230_34_n_286),
    .B(inc_u4_add_230_34_n_235),
    .Y(inc_u4_add_230_34_n_230));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g321 (.A1(u4_fract_out[9]),
    .A2(inc_u4_add_230_34_n_239),
    .B(inc_u4_add_230_34_n_235),
    .Y(n_3786));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g322 (.A(u4_fract_out[9]),
    .B(inc_u4_add_230_34_n_239),
    .Y(inc_u4_add_230_34_n_235));
 XNOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g323 (.A(inc_u4_add_230_34_n_242),
    .B(u4_fract_out[8]),
    .Y(n_3785));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g324 (.A(inc_u4_add_230_34_n_280),
    .B(inc_u4_add_230_34_n_242),
    .Y(inc_u4_add_230_34_n_239));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g325 (.A1(u4_fract_out[7]),
    .A2(inc_u4_add_230_34_n_246),
    .B(inc_u4_add_230_34_n_242),
    .Y(n_3784));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g326 (.A(u4_fract_out[7]),
    .B(inc_u4_add_230_34_n_246),
    .Y(inc_u4_add_230_34_n_242));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g327 (.A1(inc_u4_add_230_34_n_250),
    .A2(inc_u4_add_230_34_n_289),
    .B(inc_u4_add_230_34_n_246),
    .Y(n_3783));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g328 (.A(inc_u4_add_230_34_n_289),
    .B(inc_u4_add_230_34_n_250),
    .Y(inc_u4_add_230_34_n_246));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g330 (.A(u4_fract_out[5]),
    .B(inc_u4_add_230_34_n_254),
    .Y(inc_u4_add_230_34_n_250));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g331 (.A1(inc_u4_add_230_34_n_259),
    .A2(inc_u4_add_230_34_n_290),
    .B(inc_u4_add_230_34_n_254),
    .Y(n_3781));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g333 (.A(inc_u4_add_230_34_n_290),
    .B(inc_u4_add_230_34_n_259),
    .Y(inc_u4_add_230_34_n_254));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g334 (.A1(u4_fract_out[3]),
    .A2(inc_u4_add_230_34_n_263),
    .B(inc_u4_add_230_34_n_259),
    .Y(n_3780));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g335 (.A(u4_fract_out[3]),
    .B(inc_u4_add_230_34_n_263),
    .Y(inc_u4_add_230_34_n_259));
 AOI21xp33_ASAP7_75t_R inc_u4_add_230_34_g336 (.A1(inc_u4_add_230_34_n_267),
    .A2(inc_u4_add_230_34_n_274),
    .B(inc_u4_add_230_34_n_263),
    .Y(n_3779));
 NOR2xp33_ASAP7_75t_R inc_u4_add_230_34_g337 (.A(inc_u4_add_230_34_n_274),
    .B(inc_u4_add_230_34_n_267),
    .Y(inc_u4_add_230_34_n_263));
 OA21x2_ASAP7_75t_R inc_u4_add_230_34_g338 (.A1(u4_fract_out[1]),
    .A2(u4_g),
    .B(inc_u4_add_230_34_n_267),
    .Y(n_3778));
 NAND2xp33_ASAP7_75t_R inc_u4_add_230_34_g339 (.A(u4_fract_out[1]),
    .B(u4_g),
    .Y(inc_u4_add_230_34_n_267));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g340 (.A(u4_fract_out[18]),
    .Y(inc_u4_add_230_34_n_270));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g341 (.A(u4_fract_out[22]),
    .Y(inc_u4_add_230_34_n_272));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g342 (.A(u4_fract_out[2]),
    .Y(inc_u4_add_230_34_n_274));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g343 (.A(u4_fract_out[14]),
    .Y(inc_u4_add_230_34_n_277));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g344 (.A(u4_fract_out[20]),
    .Y(inc_u4_add_230_34_n_278));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g345 (.A(u4_fract_out[8]),
    .Y(inc_u4_add_230_34_n_280));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g346 (.A(u4_fract_out[12]),
    .Y(inc_u4_add_230_34_n_284));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g347 (.A(u4_fract_out[10]),
    .Y(inc_u4_add_230_34_n_286));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g348 (.A(u4_fract_out[6]),
    .Y(inc_u4_add_230_34_n_289));
 INVxp33_ASAP7_75t_R inc_u4_add_230_34_g349 (.A(u4_fract_out[4]),
    .Y(inc_u4_add_230_34_n_290));
 XOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g350 (.A(inc_u4_add_230_34_n_230),
    .B(u4_fract_out[11]),
    .Y(n_3788));
 XOR2xp5_ASAP7_75t_R inc_u4_add_230_34_g351 (.A(inc_u4_add_230_34_n_254),
    .B(u4_fract_out[5]),
    .Y(n_3782));
 DFFHQNx1_ASAP7_75t_R ine_reg (.CLK(clk),
    .D(n_609),
    .QN(ine));
 DFFHQNx1_ASAP7_75t_R inf_mul2_reg (.CLK(clk),
    .D(n_2133),
    .QN(inf_mul2));
 DFFHQNx1_ASAP7_75t_R inf_mul_r_reg (.CLK(clk),
    .D(n_2219),
    .QN(inf_mul_r));
 DFFHQNx1_ASAP7_75t_R inf_reg (.CLK(clk),
    .D(n_610),
    .QN(inf));
 DFFHQNx1_ASAP7_75t_R opa_nan_r_reg (.CLK(clk),
    .D(n_2206),
    .QN(opa_nan_r));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[0]  (.CLK(clk),
    .D(n_88),
    .QN(opa_r1[0]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[10]  (.CLK(clk),
    .D(n_84),
    .QN(opa_r1[10]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[11]  (.CLK(clk),
    .D(n_77),
    .QN(opa_r1[11]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[12]  (.CLK(clk),
    .D(n_89),
    .QN(opa_r1[12]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[13]  (.CLK(clk),
    .D(n_73),
    .QN(opa_r1[13]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[14]  (.CLK(clk),
    .D(n_72),
    .QN(opa_r1[14]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[15]  (.CLK(clk),
    .D(n_81),
    .QN(opa_r1[15]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[16]  (.CLK(clk),
    .D(n_95),
    .QN(opa_r1[16]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[17]  (.CLK(clk),
    .D(n_83),
    .QN(opa_r1[17]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[18]  (.CLK(clk),
    .D(n_86),
    .QN(opa_r1[18]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[19]  (.CLK(clk),
    .D(n_85),
    .QN(opa_r1[19]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[1]  (.CLK(clk),
    .D(n_91),
    .QN(opa_r1[1]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[20]  (.CLK(clk),
    .D(n_93),
    .QN(opa_r1[20]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[21]  (.CLK(clk),
    .D(n_96),
    .QN(opa_r1[21]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[22]  (.CLK(clk),
    .D(n_76),
    .QN(opa_r1[22]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[23]  (.CLK(clk),
    .D(n_54),
    .QN(opa_r1[23]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[24]  (.CLK(clk),
    .D(n_71),
    .QN(opa_r1[24]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[25]  (.CLK(clk),
    .D(n_44),
    .QN(opa_r1[25]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[26]  (.CLK(clk),
    .D(n_41),
    .QN(opa_r1[26]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[27]  (.CLK(clk),
    .D(n_45),
    .QN(opa_r1[27]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[28]  (.CLK(clk),
    .D(n_49),
    .QN(opa_r1[28]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[29]  (.CLK(clk),
    .D(n_42),
    .QN(opa_r1[29]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[2]  (.CLK(clk),
    .D(n_78),
    .QN(opa_r1[2]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[30]  (.CLK(clk),
    .D(n_62),
    .QN(opa_r1[30]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[3]  (.CLK(clk),
    .D(n_87),
    .QN(opa_r1[3]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[4]  (.CLK(clk),
    .D(n_74),
    .QN(opa_r1[4]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[5]  (.CLK(clk),
    .D(n_82),
    .QN(opa_r1[5]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[6]  (.CLK(clk),
    .D(n_75),
    .QN(opa_r1[6]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[7]  (.CLK(clk),
    .D(n_90),
    .QN(opa_r1[7]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[8]  (.CLK(clk),
    .D(n_80),
    .QN(opa_r1[8]));
 DFFHQNx1_ASAP7_75t_R \opa_r1_reg[9]  (.CLK(clk),
    .D(n_79),
    .QN(opa_r1[9]));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[0]  (.CLK(clk),
    .D(n_14087),
    .QN(n_14088));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[10]  (.CLK(clk),
    .D(n_14107),
    .QN(n_14108));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[11]  (.CLK(clk),
    .D(n_14109),
    .QN(n_14110));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[12]  (.CLK(clk),
    .D(n_14111),
    .QN(n_14112));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[13]  (.CLK(clk),
    .D(n_14113),
    .QN(n_14114));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[14]  (.CLK(clk),
    .D(n_14115),
    .QN(n_14116));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[15]  (.CLK(clk),
    .D(n_14165),
    .QN(n_14166));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[16]  (.CLK(clk),
    .D(n_14167),
    .QN(n_14168));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[17]  (.CLK(clk),
    .D(n_14169),
    .QN(n_14170));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[18]  (.CLK(clk),
    .D(n_14171),
    .QN(n_14172));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[19]  (.CLK(clk),
    .D(n_14173),
    .QN(n_14174));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[1]  (.CLK(clk),
    .D(n_14089),
    .QN(n_14090));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[20]  (.CLK(clk),
    .D(n_14117),
    .QN(n_14118));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[21]  (.CLK(clk),
    .D(n_14119),
    .QN(n_14120));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[22]  (.CLK(clk),
    .D(n_14175),
    .QN(n_14176));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[23]  (.CLK(clk),
    .D(n_2958),
    .QN(opa_r[23]));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[24]  (.CLK(clk),
    .D(n_2962),
    .QN(opa_r[24]));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[25]  (.CLK(clk),
    .D(n_2963),
    .QN(opa_r[25]));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[26]  (.CLK(clk),
    .D(n_2975),
    .QN(opa_r[26]));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[27]  (.CLK(clk),
    .D(n_2979),
    .QN(opa_r[27]));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[28]  (.CLK(clk),
    .D(n_2977),
    .QN(opa_r[28]));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[29]  (.CLK(clk),
    .D(n_2976),
    .QN(opa_r[29]));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[2]  (.CLK(clk),
    .D(n_14091),
    .QN(n_14092));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[30]  (.CLK(clk),
    .D(n_2978),
    .QN(opa_r[30]));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[31]  (.CLK(clk),
    .D(n_2964),
    .QN(opa_r[31]));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[3]  (.CLK(clk),
    .D(n_14093),
    .QN(n_14094));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[4]  (.CLK(clk),
    .D(n_14095),
    .QN(n_14096));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[5]  (.CLK(clk),
    .D(n_14097),
    .QN(n_14098));
 DFFHQNx1_ASAP7_75t_R \opa_r_reg[6]  (.CLK(clk),
    .D(n_14099),
    .QN(n_14100));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[7]  (.CLK(clk),
    .D(n_14101),
    .QN(n_14102));
 DFFHQNx1_ASAP7_75t_SL \opa_r_reg[8]  (.CLK(clk),
    .D(n_14103),
    .QN(n_2896));
 DFFHQNx1_ASAP7_75t_L \opa_r_reg[9]  (.CLK(clk),
    .D(n_14105),
    .QN(n_14106));
 DFFHQNx1_ASAP7_75t_R opas_r1_reg (.CLK(clk),
    .D(n_725),
    .QN(opas_r1));
 DFFHQNx1_ASAP7_75t_R opas_r2_reg (.CLK(clk),
    .D(n_884),
    .QN(opas_r2));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[0]  (.CLK(clk),
    .D(n_14121),
    .QN(u6_rem_96_22_Y_u6_div_90_17_n_70));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[10]  (.CLK(clk),
    .D(n_14139),
    .QN(n_14140));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[11]  (.CLK(clk),
    .D(n_14141),
    .QN(n_14142));
 DFFHQNx2_ASAP7_75t_SL \opb_r_reg[12]  (.CLK(clk),
    .D(n_14143),
    .QN(u6_rem_96_22_Y_u6_div_90_17_n_643));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[13]  (.CLK(clk),
    .D(n_14145),
    .QN(n_14146));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[14]  (.CLK(clk),
    .D(n_14147),
    .QN(n_14148));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[15]  (.CLK(clk),
    .D(n_14149),
    .QN(n_14150));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[16]  (.CLK(clk),
    .D(n_14151),
    .QN(n_14152));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[17]  (.CLK(clk),
    .D(n_14153),
    .QN(n_14154));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[18]  (.CLK(clk),
    .D(n_14155),
    .QN(n_14156));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[19]  (.CLK(clk),
    .D(n_14157),
    .QN(u6_rem_96_22_Y_u6_div_90_17_n_674));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[1]  (.CLK(clk),
    .D(n_14123),
    .QN(n_14124));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[20]  (.CLK(clk),
    .D(n_14159),
    .QN(n_14160));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[21]  (.CLK(clk),
    .D(n_14161),
    .QN(u5_mul_69_18_n_143));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[22]  (.CLK(clk),
    .D(n_14163),
    .QN(n_14164));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[23]  (.CLK(clk),
    .D(n_2972),
    .QN(opb_r[23]));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[24]  (.CLK(clk),
    .D(n_2973),
    .QN(opb_r[24]));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[25]  (.CLK(clk),
    .D(n_2959),
    .QN(opb_r[25]));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[26]  (.CLK(clk),
    .D(n_2960),
    .QN(opb_r[26]));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[27]  (.CLK(clk),
    .D(n_2971),
    .QN(opb_r[27]));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[28]  (.CLK(clk),
    .D(n_2974),
    .QN(opb_r[28]));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[29]  (.CLK(clk),
    .D(n_2957),
    .QN(opb_r[29]));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[2]  (.CLK(clk),
    .D(n_14177),
    .QN(n_14178));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[30]  (.CLK(clk),
    .D(n_2980),
    .QN(opb_r[30]));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[31]  (.CLK(clk),
    .D(n_2961),
    .QN(opb_r[31]));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[3]  (.CLK(clk),
    .D(n_14125),
    .QN(n_14126));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[4]  (.CLK(clk),
    .D(n_14127),
    .QN(n_14128));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[5]  (.CLK(clk),
    .D(n_14129),
    .QN(n_14130));
 DFFHQNx1_ASAP7_75t_SL \opb_r_reg[6]  (.CLK(clk),
    .D(n_14131),
    .QN(n_14132));
 DFFHQNx1_ASAP7_75t_R \opb_r_reg[7]  (.CLK(clk),
    .D(n_14133),
    .QN(n_14134));
 DFFHQNx1_ASAP7_75t_L \opb_r_reg[8]  (.CLK(clk),
    .D(n_14135),
    .QN(n_14136));
 DFFHQNx2_ASAP7_75t_SL \opb_r_reg[9]  (.CLK(clk),
    .D(n_14137),
    .QN(u6_rem_96_22_Y_u6_div_90_17_n_155));
 DFFHQNx1_ASAP7_75t_R \out_reg[0]  (.CLK(clk),
    .D(n_590),
    .QN(out[0]));
 DFFHQNx1_ASAP7_75t_R \out_reg[10]  (.CLK(clk),
    .D(n_578),
    .QN(out[10]));
 DFFHQNx1_ASAP7_75t_R \out_reg[11]  (.CLK(clk),
    .D(n_577),
    .QN(out[11]));
 DFFHQNx1_ASAP7_75t_R \out_reg[12]  (.CLK(clk),
    .D(n_573),
    .QN(out[12]));
 DFFHQNx1_ASAP7_75t_R \out_reg[13]  (.CLK(clk),
    .D(n_571),
    .QN(out[13]));
 DFFHQNx1_ASAP7_75t_R \out_reg[14]  (.CLK(clk),
    .D(n_575),
    .QN(out[14]));
 DFFHQNx1_ASAP7_75t_R \out_reg[15]  (.CLK(clk),
    .D(n_574),
    .QN(out[15]));
 DFFHQNx1_ASAP7_75t_R \out_reg[16]  (.CLK(clk),
    .D(n_572),
    .QN(out[16]));
 DFFHQNx1_ASAP7_75t_R \out_reg[17]  (.CLK(clk),
    .D(n_576),
    .QN(out[17]));
 DFFHQNx1_ASAP7_75t_R \out_reg[18]  (.CLK(clk),
    .D(n_570),
    .QN(out[18]));
 DFFHQNx1_ASAP7_75t_R \out_reg[19]  (.CLK(clk),
    .D(n_569),
    .QN(out[19]));
 DFFHQNx1_ASAP7_75t_R \out_reg[1]  (.CLK(clk),
    .D(n_584),
    .QN(out[1]));
 DFFHQNx1_ASAP7_75t_R \out_reg[20]  (.CLK(clk),
    .D(n_568),
    .QN(out[20]));
 DFFHQNx1_ASAP7_75t_R \out_reg[21]  (.CLK(clk),
    .D(n_567),
    .QN(out[21]));
 SDFHx1_ASAP7_75t_R \out_reg[22]  (.CLK(clk),
    .QN(out[22]),
    .D(n_385),
    .SE(n_13),
    .SI(n_553));
 DFFHQNx1_ASAP7_75t_R \out_reg[23]  (.CLK(clk),
    .D(n_516),
    .QN(out[23]));
 DFFHQNx1_ASAP7_75t_R \out_reg[24]  (.CLK(clk),
    .D(n_523),
    .QN(out[24]));
 DFFHQNx1_ASAP7_75t_R \out_reg[25]  (.CLK(clk),
    .D(n_522),
    .QN(out[25]));
 DFFHQNx1_ASAP7_75t_R \out_reg[26]  (.CLK(clk),
    .D(n_524),
    .QN(out[26]));
 DFFHQNx1_ASAP7_75t_R \out_reg[27]  (.CLK(clk),
    .D(n_525),
    .QN(out[27]));
 DFFHQNx1_ASAP7_75t_R \out_reg[28]  (.CLK(clk),
    .D(n_521),
    .QN(out[28]));
 DFFHQNx1_ASAP7_75t_R \out_reg[29]  (.CLK(clk),
    .D(n_520),
    .QN(out[29]));
 DFFHQNx1_ASAP7_75t_R \out_reg[2]  (.CLK(clk),
    .D(n_586),
    .QN(out[2]));
 DFFHQNx1_ASAP7_75t_R \out_reg[30]  (.CLK(clk),
    .D(n_526),
    .QN(out[30]));
 DFFHQNx1_ASAP7_75t_R \out_reg[31]  (.CLK(clk),
    .D(n_619),
    .QN(out[31]));
 DFFHQNx1_ASAP7_75t_R \out_reg[3]  (.CLK(clk),
    .D(n_585),
    .QN(out[3]));
 DFFHQNx1_ASAP7_75t_R \out_reg[4]  (.CLK(clk),
    .D(n_583),
    .QN(out[4]));
 DFFHQNx1_ASAP7_75t_R \out_reg[5]  (.CLK(clk),
    .D(n_582),
    .QN(out[5]));
 DFFHQNx1_ASAP7_75t_R \out_reg[6]  (.CLK(clk),
    .D(n_581),
    .QN(out[6]));
 DFFHQNx1_ASAP7_75t_R \out_reg[7]  (.CLK(clk),
    .D(n_566),
    .QN(out[7]));
 DFFHQNx1_ASAP7_75t_R \out_reg[8]  (.CLK(clk),
    .D(n_580),
    .QN(out[8]));
 DFFHQNx1_ASAP7_75t_R \out_reg[9]  (.CLK(clk),
    .D(n_579),
    .QN(out[9]));
 DFFHQNx1_ASAP7_75t_R overflow_reg (.CLK(clk),
    .D(n_536),
    .QN(overflow));
 DFFHQNx1_ASAP7_75t_R qnan_reg (.CLK(clk),
    .D(n_397),
    .QN(qnan));
 DFFHQNx1_ASAP7_75t_R \rmode_r1_reg[0]  (.CLK(clk),
    .D(n_746),
    .QN(rmode_r1[0]));
 DFFHQNx1_ASAP7_75t_R \rmode_r1_reg[1]  (.CLK(clk),
    .D(n_743),
    .QN(rmode_r1[1]));
 DFFHQNx1_ASAP7_75t_R \rmode_r2_reg[0]  (.CLK(clk),
    .D(n_940),
    .QN(rmode_r2[0]));
 DFFHQNx1_ASAP7_75t_R \rmode_r2_reg[1]  (.CLK(clk),
    .D(n_942),
    .QN(rmode_r2[1]));
 DFFHQNx1_ASAP7_75t_R \rmode_r3_reg[0]  (.CLK(clk),
    .D(n_996),
    .QN(rmode_r3[0]));
 DFFHQNx1_ASAP7_75t_R \rmode_r3_reg[1]  (.CLK(clk),
    .D(n_1003),
    .QN(rmode_r3[1]));
 DFFHQNx1_ASAP7_75t_R sign_exe_r_reg (.CLK(clk),
    .D(n_2106),
    .QN(sign_exe_r));
 DFFHQNx1_ASAP7_75t_R sign_fasu_r_reg (.CLK(clk),
    .D(n_1954),
    .QN(sign_fasu_r));
 DFFHQNx1_ASAP7_75t_R sign_mul_r_reg (.CLK(clk),
    .D(n_1956),
    .QN(sign_mul_r));
 SDFHx1_ASAP7_75t_R sign_reg (.CLK(clk),
    .QN(sign),
    .D(n_1430),
    .SE(n_1017),
    .SI(n_1431));
 DFFHQNx1_ASAP7_75t_R snan_reg (.CLK(clk),
    .D(n_92),
    .QN(snan));
 XNOR2xp5_ASAP7_75t_R sub_327_16_g585 (.A(sub_327_16_n_450),
    .B(opa_r1[30]),
    .Y(n_3666));
 AOI21xp33_ASAP7_75t_R sub_327_16_g586 (.A1(sub_327_16_n_454),
    .A2(opa_r1[29]),
    .B(sub_327_16_n_450),
    .Y(n_3665));
 NOR2xp33_ASAP7_75t_R sub_327_16_g587 (.A(opa_r1[29]),
    .B(sub_327_16_n_454),
    .Y(sub_327_16_n_450));
 AOI21xp33_ASAP7_75t_R sub_327_16_g588 (.A1(sub_327_16_n_459),
    .A2(opa_r1[28]),
    .B(sub_327_16_n_455),
    .Y(n_3664));
 INVxp33_ASAP7_75t_R sub_327_16_g589 (.A(sub_327_16_n_455),
    .Y(sub_327_16_n_454));
 NOR2xp33_ASAP7_75t_R sub_327_16_g590 (.A(opa_r1[28]),
    .B(sub_327_16_n_459),
    .Y(sub_327_16_n_455));
 AOI21xp33_ASAP7_75t_R sub_327_16_g591 (.A1(sub_327_16_n_464),
    .A2(opa_r1[27]),
    .B(sub_327_16_n_460),
    .Y(n_3663));
 INVxp33_ASAP7_75t_R sub_327_16_g592 (.A(sub_327_16_n_460),
    .Y(sub_327_16_n_459));
 NOR2xp33_ASAP7_75t_R sub_327_16_g593 (.A(opa_r1[27]),
    .B(sub_327_16_n_464),
    .Y(sub_327_16_n_460));
 AOI21xp33_ASAP7_75t_R sub_327_16_g594 (.A1(sub_327_16_n_469),
    .A2(opa_r1[26]),
    .B(sub_327_16_n_465),
    .Y(n_3662));
 INVxp33_ASAP7_75t_R sub_327_16_g595 (.A(sub_327_16_n_465),
    .Y(sub_327_16_n_464));
 NOR2xp33_ASAP7_75t_R sub_327_16_g596 (.A(opa_r1[26]),
    .B(sub_327_16_n_469),
    .Y(sub_327_16_n_465));
 AOI21xp33_ASAP7_75t_R sub_327_16_g597 (.A1(sub_327_16_n_474),
    .A2(opa_r1[25]),
    .B(sub_327_16_n_470),
    .Y(n_3661));
 INVxp33_ASAP7_75t_R sub_327_16_g598 (.A(sub_327_16_n_470),
    .Y(sub_327_16_n_469));
 NOR2xp33_ASAP7_75t_R sub_327_16_g599 (.A(opa_r1[25]),
    .B(sub_327_16_n_474),
    .Y(sub_327_16_n_470));
 AOI21xp33_ASAP7_75t_R sub_327_16_g600 (.A1(sub_327_16_n_479),
    .A2(opa_r1[24]),
    .B(sub_327_16_n_475),
    .Y(n_3660));
 INVxp33_ASAP7_75t_R sub_327_16_g601 (.A(sub_327_16_n_475),
    .Y(sub_327_16_n_474));
 NOR2xp33_ASAP7_75t_R sub_327_16_g602 (.A(opa_r1[24]),
    .B(sub_327_16_n_479),
    .Y(sub_327_16_n_475));
 AOI21xp33_ASAP7_75t_R sub_327_16_g603 (.A1(sub_327_16_n_484),
    .A2(opa_r1[23]),
    .B(sub_327_16_n_480),
    .Y(n_3659));
 INVxp33_ASAP7_75t_R sub_327_16_g604 (.A(sub_327_16_n_480),
    .Y(sub_327_16_n_479));
 NOR2xp33_ASAP7_75t_R sub_327_16_g605 (.A(opa_r1[23]),
    .B(sub_327_16_n_484),
    .Y(sub_327_16_n_480));
 AOI21xp33_ASAP7_75t_R sub_327_16_g606 (.A1(sub_327_16_n_489),
    .A2(opa_r1[22]),
    .B(sub_327_16_n_485),
    .Y(n_3658));
 INVxp33_ASAP7_75t_R sub_327_16_g607 (.A(sub_327_16_n_485),
    .Y(sub_327_16_n_484));
 NOR2xp33_ASAP7_75t_R sub_327_16_g608 (.A(opa_r1[22]),
    .B(sub_327_16_n_489),
    .Y(sub_327_16_n_485));
 AOI21xp33_ASAP7_75t_R sub_327_16_g609 (.A1(sub_327_16_n_494),
    .A2(opa_r1[21]),
    .B(sub_327_16_n_490),
    .Y(n_3657));
 INVxp33_ASAP7_75t_R sub_327_16_g610 (.A(sub_327_16_n_490),
    .Y(sub_327_16_n_489));
 NOR2xp33_ASAP7_75t_R sub_327_16_g611 (.A(opa_r1[21]),
    .B(sub_327_16_n_494),
    .Y(sub_327_16_n_490));
 AOI21xp33_ASAP7_75t_R sub_327_16_g612 (.A1(sub_327_16_n_499),
    .A2(opa_r1[20]),
    .B(sub_327_16_n_495),
    .Y(n_3656));
 INVxp33_ASAP7_75t_R sub_327_16_g613 (.A(sub_327_16_n_495),
    .Y(sub_327_16_n_494));
 NOR2xp33_ASAP7_75t_R sub_327_16_g614 (.A(opa_r1[20]),
    .B(sub_327_16_n_499),
    .Y(sub_327_16_n_495));
 AOI21xp33_ASAP7_75t_R sub_327_16_g615 (.A1(sub_327_16_n_504),
    .A2(opa_r1[19]),
    .B(sub_327_16_n_500),
    .Y(n_3655));
 INVxp33_ASAP7_75t_R sub_327_16_g616 (.A(sub_327_16_n_500),
    .Y(sub_327_16_n_499));
 NOR2xp33_ASAP7_75t_R sub_327_16_g617 (.A(opa_r1[19]),
    .B(sub_327_16_n_504),
    .Y(sub_327_16_n_500));
 AOI21xp33_ASAP7_75t_R sub_327_16_g618 (.A1(sub_327_16_n_509),
    .A2(opa_r1[18]),
    .B(sub_327_16_n_505),
    .Y(n_3654));
 INVxp33_ASAP7_75t_R sub_327_16_g619 (.A(sub_327_16_n_505),
    .Y(sub_327_16_n_504));
 NOR2xp33_ASAP7_75t_R sub_327_16_g620 (.A(opa_r1[18]),
    .B(sub_327_16_n_509),
    .Y(sub_327_16_n_505));
 AOI21xp33_ASAP7_75t_R sub_327_16_g621 (.A1(sub_327_16_n_514),
    .A2(opa_r1[17]),
    .B(sub_327_16_n_510),
    .Y(n_3653));
 INVxp33_ASAP7_75t_R sub_327_16_g622 (.A(sub_327_16_n_510),
    .Y(sub_327_16_n_509));
 NOR2xp33_ASAP7_75t_R sub_327_16_g623 (.A(opa_r1[17]),
    .B(sub_327_16_n_514),
    .Y(sub_327_16_n_510));
 AOI21xp33_ASAP7_75t_R sub_327_16_g624 (.A1(sub_327_16_n_519),
    .A2(opa_r1[16]),
    .B(sub_327_16_n_515),
    .Y(n_3652));
 INVxp33_ASAP7_75t_R sub_327_16_g625 (.A(sub_327_16_n_515),
    .Y(sub_327_16_n_514));
 NOR2xp33_ASAP7_75t_R sub_327_16_g626 (.A(opa_r1[16]),
    .B(sub_327_16_n_519),
    .Y(sub_327_16_n_515));
 AOI21xp33_ASAP7_75t_R sub_327_16_g627 (.A1(sub_327_16_n_524),
    .A2(opa_r1[15]),
    .B(sub_327_16_n_520),
    .Y(n_3651));
 INVxp33_ASAP7_75t_R sub_327_16_g628 (.A(sub_327_16_n_520),
    .Y(sub_327_16_n_519));
 NOR2xp33_ASAP7_75t_R sub_327_16_g629 (.A(opa_r1[15]),
    .B(sub_327_16_n_524),
    .Y(sub_327_16_n_520));
 AOI21xp33_ASAP7_75t_R sub_327_16_g630 (.A1(sub_327_16_n_529),
    .A2(opa_r1[14]),
    .B(sub_327_16_n_525),
    .Y(n_3650));
 INVxp33_ASAP7_75t_R sub_327_16_g631 (.A(sub_327_16_n_525),
    .Y(sub_327_16_n_524));
 NOR2xp33_ASAP7_75t_R sub_327_16_g632 (.A(opa_r1[14]),
    .B(sub_327_16_n_529),
    .Y(sub_327_16_n_525));
 AOI21xp33_ASAP7_75t_R sub_327_16_g633 (.A1(sub_327_16_n_534),
    .A2(opa_r1[13]),
    .B(sub_327_16_n_530),
    .Y(n_3649));
 INVxp33_ASAP7_75t_R sub_327_16_g634 (.A(sub_327_16_n_530),
    .Y(sub_327_16_n_529));
 NOR2xp33_ASAP7_75t_R sub_327_16_g635 (.A(opa_r1[13]),
    .B(sub_327_16_n_534),
    .Y(sub_327_16_n_530));
 AOI21xp33_ASAP7_75t_R sub_327_16_g636 (.A1(sub_327_16_n_539),
    .A2(opa_r1[12]),
    .B(sub_327_16_n_535),
    .Y(n_3648));
 INVxp33_ASAP7_75t_R sub_327_16_g637 (.A(sub_327_16_n_535),
    .Y(sub_327_16_n_534));
 NOR2xp33_ASAP7_75t_R sub_327_16_g638 (.A(opa_r1[12]),
    .B(sub_327_16_n_539),
    .Y(sub_327_16_n_535));
 AOI21xp33_ASAP7_75t_R sub_327_16_g639 (.A1(sub_327_16_n_544),
    .A2(opa_r1[11]),
    .B(sub_327_16_n_540),
    .Y(n_3837));
 INVxp33_ASAP7_75t_R sub_327_16_g640 (.A(sub_327_16_n_540),
    .Y(sub_327_16_n_539));
 NOR2xp33_ASAP7_75t_R sub_327_16_g641 (.A(opa_r1[11]),
    .B(sub_327_16_n_544),
    .Y(sub_327_16_n_540));
 AOI21xp33_ASAP7_75t_R sub_327_16_g642 (.A1(sub_327_16_n_549),
    .A2(opa_r1[10]),
    .B(sub_327_16_n_545),
    .Y(n_3836));
 INVxp33_ASAP7_75t_R sub_327_16_g643 (.A(sub_327_16_n_545),
    .Y(sub_327_16_n_544));
 NOR2xp33_ASAP7_75t_R sub_327_16_g644 (.A(opa_r1[10]),
    .B(sub_327_16_n_549),
    .Y(sub_327_16_n_545));
 AOI21xp33_ASAP7_75t_R sub_327_16_g645 (.A1(sub_327_16_n_554),
    .A2(opa_r1[9]),
    .B(sub_327_16_n_550),
    .Y(n_3835));
 INVxp33_ASAP7_75t_R sub_327_16_g646 (.A(sub_327_16_n_550),
    .Y(sub_327_16_n_549));
 NOR2xp33_ASAP7_75t_R sub_327_16_g647 (.A(opa_r1[9]),
    .B(sub_327_16_n_554),
    .Y(sub_327_16_n_550));
 AOI21xp33_ASAP7_75t_R sub_327_16_g648 (.A1(sub_327_16_n_559),
    .A2(opa_r1[8]),
    .B(sub_327_16_n_555),
    .Y(n_3834));
 INVxp33_ASAP7_75t_R sub_327_16_g649 (.A(sub_327_16_n_555),
    .Y(sub_327_16_n_554));
 NOR2xp33_ASAP7_75t_R sub_327_16_g650 (.A(opa_r1[8]),
    .B(sub_327_16_n_559),
    .Y(sub_327_16_n_555));
 AOI21xp33_ASAP7_75t_R sub_327_16_g651 (.A1(sub_327_16_n_564),
    .A2(opa_r1[7]),
    .B(sub_327_16_n_560),
    .Y(n_3833));
 INVxp33_ASAP7_75t_R sub_327_16_g652 (.A(sub_327_16_n_560),
    .Y(sub_327_16_n_559));
 NOR2xp33_ASAP7_75t_R sub_327_16_g653 (.A(opa_r1[7]),
    .B(sub_327_16_n_564),
    .Y(sub_327_16_n_560));
 AOI21xp33_ASAP7_75t_R sub_327_16_g654 (.A1(sub_327_16_n_569),
    .A2(opa_r1[6]),
    .B(sub_327_16_n_565),
    .Y(n_3832));
 INVxp33_ASAP7_75t_R sub_327_16_g655 (.A(sub_327_16_n_565),
    .Y(sub_327_16_n_564));
 NOR2xp33_ASAP7_75t_R sub_327_16_g656 (.A(opa_r1[6]),
    .B(sub_327_16_n_569),
    .Y(sub_327_16_n_565));
 AOI21xp33_ASAP7_75t_R sub_327_16_g657 (.A1(sub_327_16_n_574),
    .A2(opa_r1[5]),
    .B(sub_327_16_n_570),
    .Y(n_3831));
 INVxp33_ASAP7_75t_R sub_327_16_g658 (.A(sub_327_16_n_570),
    .Y(sub_327_16_n_569));
 NOR2xp33_ASAP7_75t_R sub_327_16_g659 (.A(opa_r1[5]),
    .B(sub_327_16_n_574),
    .Y(sub_327_16_n_570));
 AOI21xp33_ASAP7_75t_R sub_327_16_g660 (.A1(sub_327_16_n_579),
    .A2(opa_r1[4]),
    .B(sub_327_16_n_575),
    .Y(n_3830));
 INVxp33_ASAP7_75t_R sub_327_16_g661 (.A(sub_327_16_n_575),
    .Y(sub_327_16_n_574));
 NOR2xp33_ASAP7_75t_R sub_327_16_g662 (.A(opa_r1[4]),
    .B(sub_327_16_n_579),
    .Y(sub_327_16_n_575));
 AOI21xp33_ASAP7_75t_R sub_327_16_g663 (.A1(sub_327_16_n_584),
    .A2(opa_r1[3]),
    .B(sub_327_16_n_580),
    .Y(n_3829));
 INVxp33_ASAP7_75t_R sub_327_16_g664 (.A(sub_327_16_n_580),
    .Y(sub_327_16_n_579));
 NOR2xp33_ASAP7_75t_R sub_327_16_g665 (.A(opa_r1[3]),
    .B(sub_327_16_n_584),
    .Y(sub_327_16_n_580));
 AOI21xp33_ASAP7_75t_R sub_327_16_g666 (.A1(sub_327_16_n_589),
    .A2(opa_r1[2]),
    .B(n_14564),
    .Y(n_3828));
 INVxp33_ASAP7_75t_R sub_327_16_g667 (.A(n_14564),
    .Y(sub_327_16_n_584));
 AOI21xp33_ASAP7_75t_R sub_327_16_g669 (.A1(opa_r1[1]),
    .A2(opa_r1[0]),
    .B(n_14033),
    .Y(n_3827));
 INVxp33_ASAP7_75t_R sub_327_16_g670 (.A(n_14033),
    .Y(sub_327_16_n_589));
 DFFHQNx1_ASAP7_75t_R u0_expa_00_reg (.CLK(clk),
    .D(n_13883),
    .QN(u0_expa_00));
 DFFHQNx1_ASAP7_75t_R u0_expa_ff_reg (.CLK(clk),
    .D(n_2151),
    .QN(u0_expa_ff));
 DFFHQNx1_ASAP7_75t_R u0_expb_00_reg (.CLK(clk),
    .D(fractb_mul[23]),
    .QN(u0_expb_00));
 DFFHQNx1_ASAP7_75t_R u0_expb_ff_reg (.CLK(clk),
    .D(n_2165),
    .QN(u0_expb_ff));
 DFFHQNx1_ASAP7_75t_R u0_fracta_00_reg (.CLK(clk),
    .D(n_3545),
    .QN(u0_fracta_00));
 DFFHQNx1_ASAP7_75t_R u0_fractb_00_reg (.CLK(clk),
    .D(n_2472),
    .QN(u0_fractb_00));
 DFFHQNx1_ASAP7_75t_R u0_ind_reg (.CLK(clk),
    .D(n_2496),
    .QN(ind_d));
 DFFHQNx1_ASAP7_75t_R u0_inf_reg (.CLK(clk),
    .D(n_2497),
    .QN(inf_d));
 DFFHQNx1_ASAP7_75t_R u0_infa_f_r_reg (.CLK(clk),
    .D(n_3545),
    .QN(u0_infa_f_r));
 DFFHQNx1_ASAP7_75t_R u0_infb_f_r_reg (.CLK(clk),
    .D(n_2472),
    .QN(u0_infb_f_r));
 DFFHQNx1_ASAP7_75t_R u0_opa_00_reg (.CLK(clk),
    .D(n_2098),
    .QN(opa_00));
 DFFHQNx1_ASAP7_75t_R u0_opa_dn_reg (.CLK(clk),
    .D(n_880),
    .QN(opa_dn));
 DFFHQNx1_ASAP7_75t_R u0_opa_inf_reg (.CLK(clk),
    .D(n_2194),
    .QN(opa_inf));
 DFFHQNx1_ASAP7_75t_R u0_opa_nan_reg (.CLK(clk),
    .D(n_2178),
    .QN(opa_nan));
 DFFHQNx1_ASAP7_75t_R u0_opb_00_reg (.CLK(clk),
    .D(n_2484),
    .QN(opb_00));
 DFFHQNx1_ASAP7_75t_R u0_opb_dn_reg (.CLK(clk),
    .D(n_881),
    .QN(opb_dn));
 DFFHQNx1_ASAP7_75t_R u0_opb_inf_reg (.CLK(clk),
    .D(n_2485),
    .QN(opb_inf));
 DFFHQNx1_ASAP7_75t_R u0_opb_nan_reg (.CLK(clk),
    .D(n_2475),
    .QN(opb_nan));
 DFFHQNx1_ASAP7_75t_R u0_qnan_r_a_reg (.CLK(clk),
    .D(n_802),
    .QN(u0_qnan_r_a));
 DFFHQNx1_ASAP7_75t_R u0_qnan_r_b_reg (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_584),
    .QN(u0_qnan_r_b));
 DFFHQNx1_ASAP7_75t_R u0_qnan_reg (.CLK(clk),
    .D(n_2198),
    .QN(qnan_d));
 DFFHQNx1_ASAP7_75t_R u0_snan_r_a_reg (.CLK(clk),
    .D(n_2438),
    .QN(u0_snan_r_a));
 DFFHQNx1_ASAP7_75t_R u0_snan_r_b_reg (.CLK(clk),
    .D(n_2470),
    .QN(u0_snan_r_b));
 DFFHQNx1_ASAP7_75t_R u0_snan_reg (.CLK(clk),
    .D(n_2487),
    .QN(snan_d));
 DFFHQNx1_ASAP7_75t_R u1_add_r_reg (.CLK(clk),
    .D(fpu_op_r1[0]),
    .QN(u1_add_r));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[0]  (.CLK(clk),
    .D(n_448),
    .QN(exp_fasu[0]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[1]  (.CLK(clk),
    .D(n_447),
    .QN(exp_fasu[1]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[2]  (.CLK(clk),
    .D(n_446),
    .QN(exp_fasu[2]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[3]  (.CLK(clk),
    .D(n_449),
    .QN(exp_fasu[3]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[4]  (.CLK(clk),
    .D(n_441),
    .QN(exp_fasu[4]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[5]  (.CLK(clk),
    .D(n_444),
    .QN(exp_fasu[5]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[6]  (.CLK(clk),
    .D(n_443),
    .QN(exp_fasu[6]));
 DFFHQNx1_ASAP7_75t_R \u1_exp_dn_out_reg[7]  (.CLK(clk),
    .D(n_442),
    .QN(exp_fasu[7]));
 DFFHQNx1_ASAP7_75t_R u1_fasu_op_reg (.CLK(clk),
    .D(n_3074),
    .QN(fasu_op));
 DFFHQNx1_ASAP7_75t_R u1_fracta_eq_fractb_reg (.CLK(clk),
    .D(u1_n_4702),
    .QN(u1_fracta_eq_fractb));
 DFFHQNx1_ASAP7_75t_R u1_fracta_lt_fractb_reg (.CLK(clk),
    .D(n_2469),
    .QN(u1_fracta_lt_fractb));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[10]  (.CLK(clk),
    .D(n_214),
    .QN(fracta[10]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[11]  (.CLK(clk),
    .D(n_222),
    .QN(fracta[11]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[12]  (.CLK(clk),
    .D(n_223),
    .QN(fracta[12]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[13]  (.CLK(clk),
    .D(n_224),
    .QN(fracta[13]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[14]  (.CLK(clk),
    .D(n_226),
    .QN(fracta[14]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[15]  (.CLK(clk),
    .D(n_227),
    .QN(fracta[15]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[16]  (.CLK(clk),
    .D(n_166),
    .QN(fracta[16]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[17]  (.CLK(clk),
    .D(n_187),
    .QN(fracta[17]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[18]  (.CLK(clk),
    .D(n_169),
    .QN(fracta[18]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[19]  (.CLK(clk),
    .D(n_195),
    .QN(fracta[19]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[20]  (.CLK(clk),
    .D(n_194),
    .QN(fracta[20]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[21]  (.CLK(clk),
    .D(n_193),
    .QN(fracta[21]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[22]  (.CLK(clk),
    .D(n_192),
    .QN(fracta[22]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[23]  (.CLK(clk),
    .D(n_191),
    .QN(fracta[23]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[24]  (.CLK(clk),
    .D(n_167),
    .QN(fracta[24]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[25]  (.CLK(clk),
    .D(n_190),
    .QN(fracta[25]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[26]  (.CLK(clk),
    .D(n_55),
    .QN(fracta[26]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[3]  (.CLK(clk),
    .D(n_215),
    .QN(fracta[3]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[4]  (.CLK(clk),
    .D(n_216),
    .QN(fracta[4]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[5]  (.CLK(clk),
    .D(n_217),
    .QN(fracta[5]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[6]  (.CLK(clk),
    .D(n_209),
    .QN(fracta[6]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[7]  (.CLK(clk),
    .D(n_218),
    .QN(fracta[7]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[8]  (.CLK(clk),
    .D(n_213),
    .QN(fracta[8]));
 DFFHQNx1_ASAP7_75t_R \u1_fracta_out_reg[9]  (.CLK(clk),
    .D(n_219),
    .QN(fracta[9]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[0]  (.CLK(clk),
    .D(n_486),
    .QN(fractb[0]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[10]  (.CLK(clk),
    .D(n_188),
    .QN(fractb[10]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[11]  (.CLK(clk),
    .D(n_189),
    .QN(fractb[11]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[12]  (.CLK(clk),
    .D(n_180),
    .QN(fractb[12]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[13]  (.CLK(clk),
    .D(n_173),
    .QN(fractb[13]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[14]  (.CLK(clk),
    .D(n_171),
    .QN(fractb[14]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[15]  (.CLK(clk),
    .D(n_170),
    .QN(fractb[15]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[16]  (.CLK(clk),
    .D(n_179),
    .QN(fractb[16]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[17]  (.CLK(clk),
    .D(n_178),
    .QN(fractb[17]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[18]  (.CLK(clk),
    .D(n_172),
    .QN(fractb[18]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[19]  (.CLK(clk),
    .D(n_168),
    .QN(fractb[19]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[1]  (.CLK(clk),
    .D(n_295),
    .QN(fractb[1]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[20]  (.CLK(clk),
    .D(n_177),
    .QN(fractb[20]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[21]  (.CLK(clk),
    .D(n_208),
    .QN(fractb[21]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[22]  (.CLK(clk),
    .D(n_212),
    .QN(fractb[22]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[23]  (.CLK(clk),
    .D(n_210),
    .QN(fractb[23]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[24]  (.CLK(clk),
    .D(n_175),
    .QN(fractb[24]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[25]  (.CLK(clk),
    .D(n_174),
    .QN(fractb[25]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[26]  (.CLK(clk),
    .D(u1_fractb_s[26]),
    .QN(fractb[26]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[2]  (.CLK(clk),
    .D(n_349),
    .QN(fractb[2]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[3]  (.CLK(clk),
    .D(n_186),
    .QN(fractb[3]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[4]  (.CLK(clk),
    .D(n_185),
    .QN(fractb[4]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[5]  (.CLK(clk),
    .D(n_181),
    .QN(fractb[5]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[6]  (.CLK(clk),
    .D(n_184),
    .QN(fractb[6]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[7]  (.CLK(clk),
    .D(n_176),
    .QN(fractb[7]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[8]  (.CLK(clk),
    .D(n_183),
    .QN(fractb[8]));
 DFFHQNx1_ASAP7_75t_R \u1_fractb_out_reg[9]  (.CLK(clk),
    .D(n_182),
    .QN(fractb[9]));
 DFFHQNx1_ASAP7_75t_R u1_nan_sign_reg (.CLK(clk),
    .D(n_2582),
    .QN(nan_sign_d));
 DFFHQNx1_ASAP7_75t_R u1_result_zero_sign_reg (.CLK(clk),
    .D(n_2209),
    .QN(result_zero_sign_d));
 DFFHQNx1_ASAP7_75t_R u1_sign_reg (.CLK(clk),
    .D(n_1429),
    .QN(sign_fasu));
 DFFHQNx1_ASAP7_75t_R u1_signa_r_reg (.CLK(clk),
    .D(n_725),
    .QN(u1_signa_r));
 DFFHQNx1_ASAP7_75t_R u1_signb_r_reg (.CLK(clk),
    .D(n_728),
    .QN(u1_signb_r));
 SDFHx1_ASAP7_75t_R \u2_exp_out_reg[0]  (.CLK(clk),
    .QN(exp_mul[0]),
    .D(u2_n_775),
    .SE(u2_exp_tmp1[0]),
    .SI(n_29));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[1]  (.CLK(clk),
    .D(n_390),
    .QN(exp_mul[1]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[2]  (.CLK(clk),
    .D(n_426),
    .QN(exp_mul[2]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[3]  (.CLK(clk),
    .D(n_433),
    .QN(exp_mul[3]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[4]  (.CLK(clk),
    .D(n_424),
    .QN(exp_mul[4]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[5]  (.CLK(clk),
    .D(n_434),
    .QN(exp_mul[5]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[6]  (.CLK(clk),
    .D(n_438),
    .QN(exp_mul[6]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_out_reg[7]  (.CLK(clk),
    .D(n_431),
    .QN(exp_mul[7]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_ovf_reg[0]  (.CLK(clk),
    .D(n_13844),
    .QN(exp_ovf[0]));
 DFFHQNx1_ASAP7_75t_R \u2_exp_ovf_reg[1]  (.CLK(clk),
    .D(n_1272),
    .QN(exp_ovf[1]));
 DFFHQNx1_ASAP7_75t_R u2_inf_reg (.CLK(clk),
    .D(n_2199),
    .QN(inf_mul));
 DFFHQNx1_ASAP7_75t_R u2_sign_exe_reg (.CLK(clk),
    .D(n_1972),
    .QN(sign_exe));
 SDFHx1_ASAP7_75t_R u2_sign_reg (.CLK(clk),
    .QN(sign_mul),
    .D(n_728),
    .SE(opa_r[31]),
    .SI(opb_r[31]));
 DFFHQNx1_ASAP7_75t_R \u2_underflow_reg[0]  (.CLK(clk),
    .D(n_2182),
    .QN(underflow_fmul_d[0]));
 DFFHQNx1_ASAP7_75t_R \u2_underflow_reg[1]  (.CLK(clk),
    .D(n_2489),
    .QN(underflow_fmul_d[1]));
 DFFHQNx1_ASAP7_75t_R \u2_underflow_reg[2]  (.CLK(clk),
    .D(n_2500),
    .QN(underflow_fmul_d[2]));
 INVxp67_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_drc_bufs966 (.A(fasu_op),
    .Y(u3_sub_52_45_Y_add_52_31_n_842));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g835 (.A(u3_sub_52_45_Y_add_52_31_n_633),
    .B(fracta[26]),
    .C(u3_sub_52_45_Y_add_52_31_n_790),
    .Y(u3_sub_52_45_Y_add_52_31_n_630));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g838 (.A(u3_sub_52_45_Y_add_52_31_n_636),
    .B(u3_sub_52_45_Y_add_52_31_n_829),
    .C(u3_sub_52_45_Y_add_52_31_n_771),
    .Y(u3_sub_52_45_Y_add_52_31_n_633));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g840 (.A(u3_sub_52_45_Y_add_52_31_n_639),
    .B(fracta[24]),
    .C(u3_sub_52_45_Y_add_52_31_n_786),
    .Y(u3_sub_52_45_Y_add_52_31_n_636));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g843 (.A(u3_sub_52_45_Y_add_52_31_n_642),
    .B(u3_sub_52_45_Y_add_52_31_n_817),
    .C(u3_sub_52_45_Y_add_52_31_n_773),
    .Y(u3_sub_52_45_Y_add_52_31_n_639));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g845 (.A(u3_sub_52_45_Y_add_52_31_n_645),
    .B(fracta[22]),
    .C(u3_sub_52_45_Y_add_52_31_n_793),
    .Y(u3_sub_52_45_Y_add_52_31_n_642));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g848 (.A(u3_sub_52_45_Y_add_52_31_n_648),
    .B(u3_sub_52_45_Y_add_52_31_n_803),
    .C(u3_sub_52_45_Y_add_52_31_n_789),
    .Y(u3_sub_52_45_Y_add_52_31_n_645));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g850 (.A(u3_sub_52_45_Y_add_52_31_n_651),
    .B(fracta[20]),
    .C(u3_sub_52_45_Y_add_52_31_n_782),
    .Y(u3_sub_52_45_Y_add_52_31_n_648));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g853 (.A(u3_sub_52_45_Y_add_52_31_n_654),
    .B(u3_sub_52_45_Y_add_52_31_n_831),
    .C(u3_sub_52_45_Y_add_52_31_n_775),
    .Y(u3_sub_52_45_Y_add_52_31_n_651));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g855 (.A(u3_sub_52_45_Y_add_52_31_n_657),
    .B(fracta[18]),
    .C(u3_sub_52_45_Y_add_52_31_n_770),
    .Y(u3_sub_52_45_Y_add_52_31_n_654));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g858 (.A(u3_sub_52_45_Y_add_52_31_n_660),
    .B(u3_sub_52_45_Y_add_52_31_n_819),
    .C(u3_sub_52_45_Y_add_52_31_n_774),
    .Y(u3_sub_52_45_Y_add_52_31_n_657));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g860 (.A(u3_sub_52_45_Y_add_52_31_n_663),
    .B(fracta[16]),
    .C(u3_sub_52_45_Y_add_52_31_n_794),
    .Y(u3_sub_52_45_Y_add_52_31_n_660));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g863 (.A(u3_sub_52_45_Y_add_52_31_n_666),
    .B(u3_sub_52_45_Y_add_52_31_n_809),
    .C(u3_sub_52_45_Y_add_52_31_n_791),
    .Y(u3_sub_52_45_Y_add_52_31_n_663));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g865 (.A(u3_sub_52_45_Y_add_52_31_n_669),
    .B(fracta[14]),
    .C(u3_sub_52_45_Y_add_52_31_n_795),
    .Y(u3_sub_52_45_Y_add_52_31_n_666));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g868 (.A(u3_sub_52_45_Y_add_52_31_n_672),
    .B(u3_sub_52_45_Y_add_52_31_n_812),
    .C(u3_sub_52_45_Y_add_52_31_n_778),
    .Y(u3_sub_52_45_Y_add_52_31_n_669));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g870 (.A(u3_sub_52_45_Y_add_52_31_n_675),
    .B(fracta[12]),
    .C(u3_sub_52_45_Y_add_52_31_n_772),
    .Y(u3_sub_52_45_Y_add_52_31_n_672));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g873 (.A(u3_sub_52_45_Y_add_52_31_n_678),
    .B(u3_sub_52_45_Y_add_52_31_n_824),
    .C(u3_sub_52_45_Y_add_52_31_n_781),
    .Y(u3_sub_52_45_Y_add_52_31_n_675));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g875 (.A(u3_sub_52_45_Y_add_52_31_n_681),
    .B(fracta[10]),
    .C(u3_sub_52_45_Y_add_52_31_n_777),
    .Y(u3_sub_52_45_Y_add_52_31_n_678));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g878 (.A(u3_sub_52_45_Y_add_52_31_n_684),
    .B(u3_sub_52_45_Y_add_52_31_n_807),
    .C(u3_sub_52_45_Y_add_52_31_n_779),
    .Y(u3_sub_52_45_Y_add_52_31_n_681));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g880 (.A(u3_sub_52_45_Y_add_52_31_n_687),
    .B(fracta[8]),
    .C(u3_sub_52_45_Y_add_52_31_n_776),
    .Y(u3_sub_52_45_Y_add_52_31_n_684));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g883 (.A(u3_sub_52_45_Y_add_52_31_n_690),
    .B(u3_sub_52_45_Y_add_52_31_n_798),
    .C(u3_sub_52_45_Y_add_52_31_n_780),
    .Y(u3_sub_52_45_Y_add_52_31_n_687));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g885 (.A(u3_sub_52_45_Y_add_52_31_n_693),
    .B(fracta[6]),
    .C(u3_sub_52_45_Y_add_52_31_n_796),
    .Y(u3_sub_52_45_Y_add_52_31_n_690));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g888 (.A(u3_sub_52_45_Y_add_52_31_n_696),
    .B(u3_sub_52_45_Y_add_52_31_n_821),
    .C(u3_sub_52_45_Y_add_52_31_n_787),
    .Y(u3_sub_52_45_Y_add_52_31_n_693));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g890 (.A(u3_sub_52_45_Y_add_52_31_n_698),
    .B(fracta[4]),
    .C(u3_sub_52_45_Y_add_52_31_n_788),
    .Y(u3_sub_52_45_Y_add_52_31_n_696));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g892 (.A(u3_sub_52_45_Y_add_52_31_n_699),
    .Y(u3_sub_52_45_Y_add_52_31_n_698));
 MAJIxp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g893 (.A(u3_sub_52_45_Y_add_52_31_n_702),
    .B(fracta[3]),
    .C(u3_sub_52_45_Y_add_52_31_n_792),
    .Y(u3_sub_52_45_Y_add_52_31_n_699));
 NOR2xp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g907 (.A(u3_sub_52_45_Y_add_52_31_n_784),
    .B(u3_sub_52_45_Y_add_52_31_n_767),
    .Y(u3_sub_52_45_Y_add_52_31_n_702));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g919 (.A(u3_sub_52_45_Y_add_52_31_n_788),
    .B(fracta[4]),
    .Y(u3_sub_52_45_Y_add_52_31_n_762));
 NAND2xp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g921 (.A(u3_sub_52_45_Y_add_52_31_n_797),
    .B(u3_sub_52_45_Y_add_52_31_n_785),
    .Y(u3_sub_52_45_Y_add_52_31_n_767));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g922 (.A(fractb[18]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_770));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g923 (.A(fractb[25]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_771));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g924 (.A(fractb[12]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_772));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g925 (.A(fractb[23]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_773));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g926 (.A(fractb[17]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_774));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g927 (.A(fractb[19]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_775));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g928 (.A(fractb[8]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_776));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g929 (.A(fractb[10]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_777));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g930 (.A(fractb[13]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_778));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g931 (.A(fractb[9]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_779));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g932 (.A(fractb[7]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_780));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g933 (.A(fractb[11]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_781));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g934 (.A(fractb[20]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_782));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g935 (.A(fractb[2]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_784));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g936 (.A(fractb[1]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_785));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g937 (.A(fractb[24]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_786));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g938 (.A(fractb[5]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_787));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g939 (.A(fractb[4]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_788));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g940 (.A(fractb[21]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_789));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g941 (.A(fractb[26]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_790));
 XNOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g942 (.A(fractb[15]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_791));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g943 (.A(fractb[3]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_792));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g944 (.A(fractb[22]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_793));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g945 (.A(fractb[16]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_794));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g946 (.A(fractb[14]),
    .B(u3_sub_52_45_Y_add_52_31_n_841),
    .Y(u3_sub_52_45_Y_add_52_31_n_795));
 XOR2xp5_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g947 (.A(fractb[6]),
    .B(u3_sub_52_45_Y_add_52_31_n_842),
    .Y(u3_sub_52_45_Y_add_52_31_n_796));
 NOR2xp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g948 (.A(fasu_op),
    .B(fractb[0]),
    .Y(u3_sub_52_45_Y_add_52_31_n_797));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g949 (.A(fracta[7]),
    .Y(u3_sub_52_45_Y_add_52_31_n_798));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g950 (.A(fracta[21]),
    .Y(u3_sub_52_45_Y_add_52_31_n_803));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g951 (.A(fracta[9]),
    .Y(u3_sub_52_45_Y_add_52_31_n_807));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g952 (.A(fracta[15]),
    .Y(u3_sub_52_45_Y_add_52_31_n_809));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g953 (.A(fracta[13]),
    .Y(u3_sub_52_45_Y_add_52_31_n_812));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g955 (.A(fracta[23]),
    .Y(u3_sub_52_45_Y_add_52_31_n_817));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g956 (.A(fracta[17]),
    .Y(u3_sub_52_45_Y_add_52_31_n_819));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g957 (.A(fracta[5]),
    .Y(u3_sub_52_45_Y_add_52_31_n_821));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g958 (.A(fracta[11]),
    .Y(u3_sub_52_45_Y_add_52_31_n_824));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g959 (.A(fracta[25]),
    .Y(u3_sub_52_45_Y_add_52_31_n_829));
 INVxp33_ASAP7_75t_R u3_sub_52_45_Y_add_52_31_g960 (.A(fracta[19]),
    .Y(u3_sub_52_45_Y_add_52_31_n_831));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker (.A(u4_fract_out_pl1[23]),
    .Y(u4_n_1792));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker599 (.A(u4_n_1454),
    .Y(u4_n_1793));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker600 (.A(u4_fract_out[11]),
    .Y(u4_n_1794));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker601 (.A(u4_fract_out[12]),
    .Y(u4_n_1795));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker602 (.A(u4_fract_out[13]),
    .Y(u4_n_1796));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker603 (.A(u4_fract_out[14]),
    .Y(u4_n_1797));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker604 (.A(u4_fract_out[15]),
    .Y(u4_n_1798));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker605 (.A(u4_fract_out[16]),
    .Y(u4_n_1799));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker606 (.A(u4_fract_out[17]),
    .Y(u4_n_1800));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker607 (.A(u4_fract_out[18]),
    .Y(u4_n_1801));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker608 (.A(u4_fract_out[19]),
    .Y(u4_n_1802));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker609 (.A(u4_fract_out[20]),
    .Y(u4_n_1803));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker610 (.A(u4_fract_out[21]),
    .Y(u4_n_1804));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker611 (.A(u4_fract_out[22]),
    .Y(u4_n_1805));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker612 (.A(u4_g),
    .Y(u4_n_1806));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker613 (.A(u4_fract_out[1]),
    .Y(u4_n_1807));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker614 (.A(u4_fract_out[2]),
    .Y(u4_n_1808));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker615 (.A(u4_fract_out[3]),
    .Y(u4_n_1809));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker616 (.A(u4_fract_out[4]),
    .Y(u4_n_1810));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker617 (.A(u4_fract_out[5]),
    .Y(u4_n_1811));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker618 (.A(u4_fract_out[6]),
    .Y(u4_n_1812));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker619 (.A(u4_fract_out[7]),
    .Y(u4_n_1813));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker620 (.A(u4_fract_out[8]),
    .Y(u4_n_1814));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker621 (.A(u4_fract_out[9]),
    .Y(u4_n_1815));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker622 (.A(u4_fract_out[10]),
    .Y(u4_n_1816));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker623 (.A(u4_n_1454),
    .Y(u4_n_1817));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker624 (.A(u4_fract_trunc[13]),
    .Y(u4_n_1818));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker625 (.A(u4_fract_trunc[14]),
    .Y(u4_n_1819));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker626 (.A(u4_fract_trunc[15]),
    .Y(u4_n_1820));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker627 (.A(u4_fract_trunc[16]),
    .Y(u4_n_1821));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker628 (.A(u4_fract_trunc[17]),
    .Y(u4_n_1822));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker629 (.A(u4_fract_trunc[18]),
    .Y(u4_n_1823));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker630 (.A(u4_fract_trunc[19]),
    .Y(u4_n_1824));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker631 (.A(u4_fract_trunc[20]),
    .Y(u4_n_1825));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker632 (.A(u4_fract_trunc[21]),
    .Y(u4_n_1826));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker633 (.A(u4_fract_trunc[22]),
    .Y(u4_n_1827));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker634 (.A(u4_fract_trunc[23]),
    .Y(u4_n_1828));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker635 (.A(u4_fract_trunc[24]),
    .Y(u4_n_1829));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker636 (.A(u4_n_1248),
    .Y(u4_n_1830));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker637 (.A(u4_fract_out[7]),
    .Y(u4_n_1831));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker638 (.A(u4_fract_out[8]),
    .Y(u4_n_1832));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker639 (.A(u4_fract_out[9]),
    .Y(u4_n_1833));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker640 (.A(u4_fract_out[10]),
    .Y(u4_n_1834));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker641 (.A(u4_fract_out[11]),
    .Y(u4_n_1835));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker642 (.A(u4_fract_out[12]),
    .Y(u4_n_1836));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker643 (.A(u4_fract_out[13]),
    .Y(u4_n_1837));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker644 (.A(u4_fract_out[14]),
    .Y(u4_n_1838));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker645 (.A(u4_fract_out[15]),
    .Y(u4_n_1839));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker646 (.A(u4_fract_out[16]),
    .Y(u4_n_1840));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker647 (.A(u4_fract_out[17]),
    .Y(u4_n_1841));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker648 (.A(u4_fract_out[18]),
    .Y(u4_n_1842));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker649 (.A(u4_fract_out[19]),
    .Y(u4_n_1843));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker650 (.A(u4_fract_out[20]),
    .Y(u4_n_1844));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker651 (.A(u4_fract_out[21]),
    .Y(u4_n_1845));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker652 (.A(u4_fract_out[22]),
    .Y(u4_n_1846));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker653 (.A(n_3490),
    .Y(u4_n_1847));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker654 (.A(n_3491),
    .Y(u4_n_1848));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker655 (.A(u4_n_1439),
    .Y(u4_n_1849));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker656 (.A(u4_n_1438),
    .Y(u4_n_1850));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker657 (.A(u4_n_1266),
    .Y(u4_n_1851));
 HB1xp67_ASAP7_75t_SL u4_cdn_loop_breaker658 (.A(u4_n_1442),
    .Y(u4_n_1852));
 INVxp33_ASAP7_75t_R u4_sll_315_50_drc_bufs4549 (.A(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_3));
 INVxp33_ASAP7_75t_R u4_sll_315_50_drc_bufs4550 (.A(u4_sll_315_50_n_17),
    .Y(u4_sll_315_50_n_5));
 INVxp33_ASAP7_75t_R u4_sll_315_50_drc_bufs4556 (.A(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_1));
 INVxp33_ASAP7_75t_R u4_sll_315_50_drc_bufs4557 (.A(n_3820),
    .Y(u4_sll_315_50_n_6));
 INVxp33_ASAP7_75t_R u4_sll_315_50_drc_bufs4562 (.A(u4_sll_315_50_n_9),
    .Y(u4_sll_315_50_n_8));
 HB1xp67_ASAP7_75t_R u4_sll_315_50_drc_bufs4570 (.A(n_3819),
    .Y(u4_sll_315_50_n_11));
 HB1xp67_ASAP7_75t_R u4_sll_315_50_drc_bufs4586 (.A(u4_sll_315_50_n_16),
    .Y(u4_sll_315_50_n_0));
 A2O1A1Ixp33_ASAP7_75t_R u4_sll_315_50_g4263 (.A1(u4_sll_315_50_n_176),
    .A2(u4_sll_315_50_n_218),
    .B(n_3753),
    .C(u4_sll_315_50_n_213),
    .Y(n_3744));
 NAND3xp33_ASAP7_75t_R u4_sll_315_50_g4264 (.A(u4_sll_315_50_n_216),
    .B(u4_sll_315_50_n_168),
    .C(u4_sll_315_50_n_103),
    .Y(n_3748));
 NAND3xp33_ASAP7_75t_R u4_sll_315_50_g4265 (.A(u4_sll_315_50_n_214),
    .B(u4_sll_315_50_n_167),
    .C(u4_sll_315_50_n_103),
    .Y(n_3747));
 OAI311xp33_ASAP7_75t_R u4_sll_315_50_g4266 (.A1(u4_sll_315_50_n_68),
    .A2(n_3753),
    .A3(u4_sll_315_50_n_151),
    .B1(u4_sll_315_50_n_169),
    .C1(u4_sll_315_50_n_217),
    .Y(n_3743));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4267 (.A1(n_3753),
    .A2(u4_sll_315_50_n_219),
    .B1(u4_sll_315_50_n_30),
    .B2(u4_sll_315_50_n_205),
    .Y(n_3746));
 OAI311xp33_ASAP7_75t_R u4_sll_315_50_g4268 (.A1(u4_sll_315_50_n_34),
    .A2(n_3752),
    .A3(n_3751),
    .B1(u4_sll_315_50_n_153),
    .C1(u4_sll_315_50_n_215),
    .Y(n_3749));
 OAI322xp33_ASAP7_75t_R u4_sll_315_50_g4269 (.A1(u4_sll_315_50_n_201),
    .A2(n_3753),
    .A3(n_3752),
    .B1(u4_sll_315_50_n_194),
    .B2(u4_sll_315_50_n_31),
    .C1(u4_sll_315_50_n_212),
    .C2(u4_sll_315_50_n_30),
    .Y(n_3750));
 OAI322xp33_ASAP7_75t_R u4_sll_315_50_g4270 (.A1(u4_sll_315_50_n_207),
    .A2(n_3753),
    .A3(n_3752),
    .B1(u4_sll_315_50_n_193),
    .B2(u4_sll_315_50_n_31),
    .C1(u4_sll_315_50_n_204),
    .C2(u4_sll_315_50_n_30),
    .Y(n_3745));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4271 (.A1(u4_sll_315_50_n_160),
    .A2(n_3752),
    .B1(u4_sll_315_50_n_76),
    .B2(u4_sll_315_50_n_138),
    .C(u4_sll_315_50_n_209),
    .Y(u4_sll_315_50_n_219));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4272 (.A1(u4_sll_315_50_n_67),
    .A2(u4_sll_315_50_n_152),
    .B1(u4_sll_315_50_n_70),
    .B2(u4_sll_315_50_n_137),
    .C(u4_sll_315_50_n_208),
    .Y(u4_sll_315_50_n_218));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4273 (.A1(u4_sll_315_50_n_206),
    .A2(n_3753),
    .B1(u4_sll_315_50_n_102),
    .B2(u4_sll_315_50_n_114),
    .C(u4_sll_315_50_n_202),
    .Y(u4_sll_315_50_n_217));
 AOI21xp33_ASAP7_75t_R u4_sll_315_50_g4274 (.A1(u4_sll_315_50_n_102),
    .A2(u4_sll_315_50_n_136),
    .B(u4_sll_315_50_n_210),
    .Y(u4_sll_315_50_n_216));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4275 (.A1(u4_sll_315_50_n_197),
    .A2(n_3753),
    .B1(u4_sll_315_50_n_102),
    .B2(u4_sll_315_50_n_115),
    .C(u4_sll_315_50_n_200),
    .Y(u4_sll_315_50_n_215));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4276 (.A1(u4_sll_315_50_n_198),
    .A2(n_3753),
    .B1(u4_sll_315_50_n_101),
    .B2(u4_sll_315_50_n_150),
    .C(u4_sll_315_50_n_195),
    .Y(u4_sll_315_50_n_214));
 A2O1A1Ixp33_ASAP7_75t_R u4_sll_315_50_g4277 (.A1(u4_sll_315_50_n_127),
    .A2(u4_sll_315_50_n_74),
    .B(u4_sll_315_50_n_196),
    .C(n_3753),
    .Y(u4_sll_315_50_n_213));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4278 (.A(u4_sll_315_50_n_211),
    .Y(u4_sll_315_50_n_212));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4279 (.A1(n_3752),
    .A2(u4_sll_315_50_n_199),
    .B1(u4_sll_315_50_n_13),
    .B2(u4_sll_315_50_n_179),
    .Y(u4_sll_315_50_n_211));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4280 (.A1(u4_sll_315_50_n_30),
    .A2(u4_sll_315_50_n_203),
    .B1(u4_sll_315_50_n_31),
    .B2(u4_sll_315_50_n_191),
    .Y(u4_sll_315_50_n_210));
 A2O1A1Ixp33_ASAP7_75t_R u4_sll_315_50_g4281 (.A1(u4_sll_315_50_n_99),
    .A2(u4_sll_315_50_n_187),
    .B(n_3752),
    .C(u4_sll_315_50_n_157),
    .Y(u4_sll_315_50_n_209));
 AOI21xp33_ASAP7_75t_R u4_sll_315_50_g4282 (.A1(u4_sll_315_50_n_155),
    .A2(u4_sll_315_50_n_188),
    .B(u4_sll_315_50_n_13),
    .Y(u4_sll_315_50_n_208));
 AND2x2_ASAP7_75t_R u4_sll_315_50_g4283 (.A(u4_sll_315_50_n_99),
    .B(u4_sll_315_50_n_189),
    .Y(u4_sll_315_50_n_207));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4284 (.A(u4_sll_315_50_n_175),
    .B(u4_sll_315_50_n_186),
    .Y(u4_sll_315_50_n_206));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4285 (.A1(u4_sll_315_50_n_67),
    .A2(u4_sll_315_50_n_143),
    .B1(u4_sll_315_50_n_74),
    .B2(u4_sll_315_50_n_109),
    .C(u4_sll_315_50_n_185),
    .Y(u4_sll_315_50_n_205));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4286 (.A1(u4_sll_315_50_n_70),
    .A2(u4_sll_315_50_n_142),
    .B1(u4_sll_315_50_n_76),
    .B2(u4_sll_315_50_n_147),
    .C(u4_sll_315_50_n_190),
    .Y(u4_sll_315_50_n_204));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4287 (.A1(u4_sll_315_50_n_76),
    .A2(u4_sll_315_50_n_127),
    .B1(u4_sll_315_50_n_70),
    .B2(u4_sll_315_50_n_128),
    .C(u4_sll_315_50_n_184),
    .Y(u4_sll_315_50_n_203));
 AOI21xp33_ASAP7_75t_R u4_sll_315_50_g4288 (.A1(u4_sll_315_50_n_164),
    .A2(u4_sll_315_50_n_182),
    .B(u4_sll_315_50_n_31),
    .Y(u4_sll_315_50_n_202));
 OAI21xp33_ASAP7_75t_R u4_sll_315_50_g4289 (.A1(fract_denorm[47]),
    .A2(n_3751),
    .B(u4_sll_315_50_n_192),
    .Y(u4_sll_315_50_n_201));
 AOI21xp33_ASAP7_75t_R u4_sll_315_50_g4290 (.A1(u4_sll_315_50_n_161),
    .A2(u4_sll_315_50_n_178),
    .B(u4_sll_315_50_n_31),
    .Y(u4_sll_315_50_n_200));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4291 (.A1(u4_sll_315_50_n_37),
    .A2(u4_sll_315_50_n_133),
    .B1(u4_sll_315_50_n_32),
    .B2(u4_sll_315_50_n_110),
    .C(u4_sll_315_50_n_181),
    .Y(u4_sll_315_50_n_199));
 NAND3xp33_ASAP7_75t_R u4_sll_315_50_g4292 (.A(u4_sll_315_50_n_171),
    .B(u4_sll_315_50_n_158),
    .C(u4_sll_315_50_n_170),
    .Y(u4_sll_315_50_n_198));
 NAND3xp33_ASAP7_75t_R u4_sll_315_50_g4293 (.A(u4_sll_315_50_n_159),
    .B(u4_sll_315_50_n_173),
    .C(u4_sll_315_50_n_174),
    .Y(u4_sll_315_50_n_197));
 OAI311xp33_ASAP7_75t_R u4_sll_315_50_g4294 (.A1(u4_sll_315_50_n_75),
    .A2(u4_sll_315_50_n_17),
    .A3(u4_sll_315_50_n_39),
    .B1(u4_sll_315_50_n_156),
    .C1(u4_sll_315_50_n_177),
    .Y(u4_sll_315_50_n_196));
 AOI21xp33_ASAP7_75t_R u4_sll_315_50_g4295 (.A1(u4_sll_315_50_n_162),
    .A2(u4_sll_315_50_n_180),
    .B(u4_sll_315_50_n_31),
    .Y(u4_sll_315_50_n_195));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4296 (.A1(u4_sll_315_50_n_36),
    .A2(u4_sll_315_50_n_131),
    .B1(u4_sll_315_50_n_33),
    .B2(u4_sll_315_50_n_138),
    .C(u4_sll_315_50_n_165),
    .Y(u4_sll_315_50_n_194));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4297 (.A1(u4_sll_315_50_n_36),
    .A2(u4_sll_315_50_n_104),
    .B1(u4_sll_315_50_n_33),
    .B2(u4_sll_315_50_n_105),
    .C(u4_sll_315_50_n_166),
    .Y(u4_sll_315_50_n_193));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4298 (.A(n_3751),
    .B(u4_sll_315_50_n_183),
    .Y(u4_sll_315_50_n_192));
 AOI221xp5_ASAP7_75t_R u4_sll_315_50_g4299 (.A1(u4_sll_315_50_n_36),
    .A2(u4_sll_315_50_n_129),
    .B1(u4_sll_315_50_n_33),
    .B2(u4_sll_315_50_n_130),
    .C(u4_sll_315_50_n_163),
    .Y(u4_sll_315_50_n_191));
 AO222x2_ASAP7_75t_R u4_sll_315_50_g4300 (.A1(u4_sll_315_50_n_72),
    .A2(u4_sll_315_50_n_144),
    .B1(u4_sll_315_50_n_67),
    .B2(u4_sll_315_50_n_140),
    .C1(u4_sll_315_50_n_74),
    .C2(u4_sll_315_50_n_146),
    .Y(u4_sll_315_50_n_190));
 AOI222xp33_ASAP7_75t_R u4_sll_315_50_g4301 (.A1(u4_sll_315_50_n_33),
    .A2(u4_sll_315_50_n_121),
    .B1(u4_sll_315_50_n_37),
    .B2(u4_sll_315_50_n_148),
    .C1(u4_sll_315_50_n_32),
    .C2(u4_sll_315_50_n_115),
    .Y(u4_sll_315_50_n_189));
 AOI222xp33_ASAP7_75t_R u4_sll_315_50_g4302 (.A1(u4_sll_315_50_n_33),
    .A2(u4_sll_315_50_n_132),
    .B1(u4_sll_315_50_n_32),
    .B2(u4_sll_315_50_n_134),
    .C1(u4_sll_315_50_n_37),
    .C2(u4_sll_315_50_n_124),
    .Y(u4_sll_315_50_n_188));
 AOI222xp33_ASAP7_75t_R u4_sll_315_50_g4303 (.A1(u4_sll_315_50_n_33),
    .A2(u4_sll_315_50_n_118),
    .B1(u4_sll_315_50_n_37),
    .B2(u4_sll_315_50_n_131),
    .C1(u4_sll_315_50_n_32),
    .C2(u4_sll_315_50_n_113),
    .Y(u4_sll_315_50_n_187));
 AOI222xp33_ASAP7_75t_R u4_sll_315_50_g4304 (.A1(u4_sll_315_50_n_70),
    .A2(u4_sll_315_50_n_149),
    .B1(u4_sll_315_50_n_76),
    .B2(u4_sll_315_50_n_98),
    .C1(u4_sll_315_50_n_72),
    .C2(u4_sll_315_50_n_107),
    .Y(u4_sll_315_50_n_186));
 AO222x2_ASAP7_75t_R u4_sll_315_50_g4305 (.A1(u4_sll_315_50_n_72),
    .A2(u4_sll_315_50_n_133),
    .B1(u4_sll_315_50_n_76),
    .B2(u4_sll_315_50_n_122),
    .C1(u4_sll_315_50_n_70),
    .C2(u4_sll_315_50_n_110),
    .Y(u4_sll_315_50_n_185));
 OAI311xp33_ASAP7_75t_R u4_sll_315_50_g4306 (.A1(u4_sll_315_50_n_77),
    .A2(u4_sll_315_50_n_17),
    .A3(u4_sll_315_50_n_39),
    .B1(u4_sll_315_50_n_154),
    .C1(u4_sll_315_50_n_172),
    .Y(u4_sll_315_50_n_184));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4307 (.A1(n_3483),
    .A2(u4_sll_315_50_n_118),
    .B1(n_3824),
    .B2(u4_sll_315_50_n_113),
    .Y(u4_sll_315_50_n_183));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4308 (.A1(u4_sll_315_50_n_116),
    .A2(u4_sll_315_50_n_36),
    .B1(u4_sll_315_50_n_117),
    .B2(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_182));
 AO22x1_ASAP7_75t_R u4_sll_315_50_g4309 (.A1(u4_sll_315_50_n_135),
    .A2(u4_sll_315_50_n_36),
    .B1(u4_sll_315_50_n_143),
    .B2(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_181));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4310 (.A1(u4_sll_315_50_n_114),
    .A2(u4_sll_315_50_n_36),
    .B1(u4_sll_315_50_n_116),
    .B2(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_180));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4311 (.A1(u4_sll_315_50_n_109),
    .A2(u4_sll_315_50_n_36),
    .B1(u4_sll_315_50_n_122),
    .B2(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_179));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4312 (.A1(u4_sll_315_50_n_148),
    .A2(u4_sll_315_50_n_36),
    .B1(u4_sll_315_50_n_104),
    .B2(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_178));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4313 (.A1(u4_sll_315_50_n_128),
    .A2(u4_sll_315_50_n_67),
    .B1(u4_sll_315_50_n_126),
    .B2(u4_sll_315_50_n_70),
    .Y(u4_sll_315_50_n_177));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4314 (.A1(u4_sll_315_50_n_136),
    .A2(u4_sll_315_50_n_72),
    .B1(u4_sll_315_50_n_129),
    .B2(u4_sll_315_50_n_74),
    .Y(u4_sll_315_50_n_176));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4315 (.A1(u4_sll_315_50_n_112),
    .A2(u4_sll_315_50_n_67),
    .B1(u4_sll_315_50_n_108),
    .B2(u4_sll_315_50_n_74),
    .Y(u4_sll_315_50_n_175));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4316 (.A1(u4_sll_315_50_n_142),
    .A2(u4_sll_315_50_n_72),
    .B1(u4_sll_315_50_n_144),
    .B2(u4_sll_315_50_n_74),
    .Y(u4_sll_315_50_n_174));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4317 (.A1(u4_sll_315_50_n_139),
    .A2(u4_sll_315_50_n_67),
    .B1(u4_sll_315_50_n_140),
    .B2(u4_sll_315_50_n_70),
    .Y(u4_sll_315_50_n_173));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4318 (.A1(u4_sll_315_50_n_124),
    .A2(u4_sll_315_50_n_67),
    .B1(u4_sll_315_50_n_125),
    .B2(u4_sll_315_50_n_74),
    .Y(u4_sll_315_50_n_172));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4319 (.A1(u4_sll_315_50_n_111),
    .A2(u4_sll_315_50_n_67),
    .B1(u4_sll_315_50_n_112),
    .B2(u4_sll_315_50_n_70),
    .Y(u4_sll_315_50_n_171));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4320 (.A1(u4_sll_315_50_n_149),
    .A2(u4_sll_315_50_n_72),
    .B1(u4_sll_315_50_n_107),
    .B2(u4_sll_315_50_n_74),
    .Y(u4_sll_315_50_n_170));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4321 (.A1(u4_sll_315_50_n_123),
    .A2(u4_sll_315_50_n_100),
    .B1(u4_sll_315_50_n_120),
    .B2(u4_sll_315_50_n_101),
    .Y(u4_sll_315_50_n_169));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4322 (.A1(u4_sll_315_50_n_137),
    .A2(u4_sll_315_50_n_100),
    .B1(u4_sll_315_50_n_152),
    .B2(u4_sll_315_50_n_101),
    .Y(u4_sll_315_50_n_168));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4323 (.A1(u4_sll_315_50_n_120),
    .A2(u4_sll_315_50_n_100),
    .B1(u4_sll_315_50_n_123),
    .B2(u4_sll_315_50_n_102),
    .Y(u4_sll_315_50_n_167));
 AO22x1_ASAP7_75t_R u4_sll_315_50_g4324 (.A1(u4_sll_315_50_n_106),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_139),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_166));
 AO22x1_ASAP7_75t_R u4_sll_315_50_g4325 (.A1(u4_sll_315_50_n_32),
    .A2(u4_sll_315_50_n_141),
    .B1(u4_sll_315_50_n_145),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_165));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4326 (.A1(u4_sll_315_50_n_119),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_111),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_164));
 AO22x1_ASAP7_75t_R u4_sll_315_50_g4327 (.A1(u4_sll_315_50_n_132),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_134),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_163));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4328 (.A1(u4_sll_315_50_n_117),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_119),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_162));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4329 (.A1(u4_sll_315_50_n_105),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_106),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_161));
 AO22x1_ASAP7_75t_R u4_sll_315_50_g4330 (.A1(u4_sll_315_50_n_145),
    .A2(u4_sll_315_50_n_32),
    .B1(u4_sll_315_50_n_135),
    .B2(u4_sll_315_50_n_37),
    .Y(u4_sll_315_50_n_160));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4331 (.A1(u4_sll_315_50_n_146),
    .A2(u4_sll_315_50_n_76),
    .B1(u4_sll_315_50_n_147),
    .B2(u4_sll_315_50_n_78),
    .Y(u4_sll_315_50_n_159));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4332 (.A1(u4_sll_315_50_n_108),
    .A2(u4_sll_315_50_n_76),
    .B1(u4_sll_315_50_n_98),
    .B2(u4_sll_315_50_n_78),
    .Y(u4_sll_315_50_n_158));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4333 (.A(u4_sll_315_50_n_141),
    .B(u4_sll_315_50_n_78),
    .Y(u4_sll_315_50_n_157));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4334 (.A(u4_sll_315_50_n_125),
    .B(u4_sll_315_50_n_72),
    .Y(u4_sll_315_50_n_156));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4335 (.A(u4_sll_315_50_n_130),
    .B(u4_sll_315_50_n_36),
    .Y(u4_sll_315_50_n_155));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4336 (.A(u4_sll_315_50_n_126),
    .B(u4_sll_315_50_n_72),
    .Y(u4_sll_315_50_n_154));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4337 (.A(u4_sll_315_50_n_121),
    .B(u4_sll_315_50_n_100),
    .Y(u4_sll_315_50_n_153));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4338 (.A(u4_sll_315_50_n_150),
    .Y(u4_sll_315_50_n_151));
 OAI21xp33_ASAP7_75t_R u4_sll_315_50_g4339 (.A1(u4_sll_315_50_n_84),
    .A2(u4_sll_315_50_n_2),
    .B(u4_sll_315_50_n_35),
    .Y(u4_sll_315_50_n_152));
 OAI21xp33_ASAP7_75t_R u4_sll_315_50_g4340 (.A1(u4_sll_315_50_n_91),
    .A2(u4_sll_315_50_n_2),
    .B(u4_sll_315_50_n_35),
    .Y(u4_sll_315_50_n_150));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4341 (.A1(u4_sll_315_50_n_64),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_65),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_149));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4342 (.A1(u4_sll_315_50_n_42),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_81),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_148));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4343 (.A1(u4_sll_315_50_n_88),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_38),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_147));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4344 (.A1(u4_sll_315_50_n_94),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_89),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_146));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4345 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_52),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_93),
    .Y(u4_sll_315_50_n_145));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4346 (.A1(u4_sll_315_50_n_65),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_97),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_144));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4347 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_48),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_80),
    .Y(u4_sll_315_50_n_143));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4348 (.A1(u4_sll_315_50_n_82),
    .A2(u4_sll_315_50_n_0),
    .B1(u4_sll_315_50_n_64),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_142));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4349 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_59),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_61),
    .Y(u4_sll_315_50_n_141));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4350 (.A1(u4_sll_315_50_n_60),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_62),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_140));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4351 (.A1(u4_sll_315_50_n_57),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_58),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_139));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4352 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_56),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_53),
    .Y(u4_sll_315_50_n_138));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4353 (.A1(u4_sll_315_50_n_43),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_54),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_137));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4354 (.A1(u4_sll_315_50_n_92),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_45),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_136));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4355 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_49),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_41),
    .Y(u4_sll_315_50_n_135));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4356 (.A1(u4_sll_315_50_n_93),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_49),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_134));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4357 (.A1(u4_sll_315_50_n_79),
    .A2(u4_sll_315_50_n_1),
    .B1(u4_sll_315_50_n_51),
    .B2(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_133));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4358 (.A1(u4_sll_315_50_n_61),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_52),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_132));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4359 (.A1(u4_sll_315_50_n_45),
    .A2(u4_sll_315_50_n_1),
    .B1(u4_sll_315_50_n_40),
    .B2(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_131));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4360 (.A1(u4_sll_315_50_n_53),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_59),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_130));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4361 (.A1(u4_sll_315_50_n_40),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_56),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_129));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4362 (.A1(u4_sll_315_50_n_80),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_47),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_128));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4363 (.A1(u4_sll_315_50_n_95),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_55),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_127));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4364 (.A1(u4_sll_315_50_n_66),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_79),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_126));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4365 (.A1(u4_sll_315_50_n_51),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_96),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_125));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4366 (.A1(u4_sll_315_50_n_41),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_48),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_124));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4367 (.A1(u4_sll_315_50_n_86),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_42),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_123));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4368 (.A1(u4_sll_315_50_n_55),
    .A2(u4_sll_315_50_n_1),
    .B1(u4_sll_315_50_n_39),
    .B2(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_122));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4369 (.A1(u4_sll_315_50_n_91),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_87),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_121));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4370 (.A1(u4_sll_315_50_n_87),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_44),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_120));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4371 (.A1(u4_sll_315_50_n_85),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_57),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_119));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4372 (.A1(u4_sll_315_50_n_84),
    .A2(u4_sll_315_50_n_1),
    .B1(u4_sll_315_50_n_43),
    .B2(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_118));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4373 (.A1(u4_sll_315_50_n_50),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_90),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_117));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4374 (.A1(u4_sll_315_50_n_46),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_63),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_116));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4375 (.A1(u4_sll_315_50_n_44),
    .A2(u4_sll_315_50_n_17),
    .B1(u4_sll_315_50_n_86),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_115));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4376 (.A1(u4_sll_315_50_n_81),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_83),
    .B2(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_114));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4377 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_54),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_92),
    .Y(u4_sll_315_50_n_113));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4378 (.A1(u4_sll_315_50_n_62),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_82),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_112));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4379 (.A1(u4_sll_315_50_n_58),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_60),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_111));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4380 (.A1(u4_sll_315_50_n_1),
    .A2(u4_sll_315_50_n_47),
    .B1(u4_sll_315_50_n_6),
    .B2(u4_sll_315_50_n_66),
    .Y(u4_sll_315_50_n_110));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4381 (.A1(u4_sll_315_50_n_96),
    .A2(u4_sll_315_50_n_1),
    .B1(u4_sll_315_50_n_95),
    .B2(u4_sll_315_50_n_6),
    .Y(u4_sll_315_50_n_109));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4382 (.A1(u4_sll_315_50_n_89),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_88),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_108));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4383 (.A1(u4_sll_315_50_n_97),
    .A2(u4_sll_315_50_n_16),
    .B1(u4_sll_315_50_n_94),
    .B2(u4_sll_315_50_n_4),
    .Y(u4_sll_315_50_n_107));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4384 (.A1(u4_sll_315_50_n_90),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_85),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_106));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4385 (.A1(u4_sll_315_50_n_63),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_50),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_105));
 OAI22xp33_ASAP7_75t_R u4_sll_315_50_g4386 (.A1(u4_sll_315_50_n_83),
    .A2(u4_sll_315_50_n_3),
    .B1(u4_sll_315_50_n_46),
    .B2(u4_sll_315_50_n_5),
    .Y(u4_sll_315_50_n_104));
 OR2x2_ASAP7_75t_R u4_sll_315_50_g4387 (.A(u4_sll_315_50_n_68),
    .B(u4_sll_315_50_n_34),
    .Y(u4_sll_315_50_n_103));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4388 (.A(n_3753),
    .B(u4_sll_315_50_n_73),
    .Y(u4_sll_315_50_n_102));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4389 (.A(n_3753),
    .B(u4_sll_315_50_n_69),
    .Y(u4_sll_315_50_n_101));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4390 (.A(n_3753),
    .B(u4_sll_315_50_n_71),
    .Y(u4_sll_315_50_n_100));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4391 (.A(u4_sll_315_50_n_77),
    .Y(u4_sll_315_50_n_78));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4392 (.A(u4_sll_315_50_n_75),
    .Y(u4_sll_315_50_n_76));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4393 (.A(u4_sll_315_50_n_73),
    .Y(u4_sll_315_50_n_74));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4394 (.A(u4_sll_315_50_n_71),
    .Y(u4_sll_315_50_n_72));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4395 (.A(u4_sll_315_50_n_69),
    .Y(u4_sll_315_50_n_70));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4396 (.A(u4_sll_315_50_n_68),
    .Y(u4_sll_315_50_n_67));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4397 (.A(fract_denorm[47]),
    .B(u4_sll_315_50_n_36),
    .Y(u4_sll_315_50_n_99));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4398 (.A(u4_sll_315_50_n_38),
    .B(u4_sll_315_50_n_0),
    .Y(u4_sll_315_50_n_98));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4399 (.A1(fract_denorm[8]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[7]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_97));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4400 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[7]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[6]),
    .Y(u4_sll_315_50_n_96));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4401 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[5]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[4]),
    .Y(u4_sll_315_50_n_95));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4402 (.A1(fract_denorm[6]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[5]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_94));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4403 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[25]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[24]),
    .Y(u4_sll_315_50_n_93));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4404 (.A1(u4_sll_315_50_n_7),
    .A2(fract_denorm[41]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[40]),
    .Y(u4_sll_315_50_n_92));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4405 (.A1(fract_denorm[46]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[45]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_91));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4406 (.A1(fract_denorm[26]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[25]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_90));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4407 (.A1(fract_denorm[4]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[3]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_89));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4408 (.A1(fract_denorm[2]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[1]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_88));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4409 (.A1(fract_denorm[44]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[43]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_87));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4410 (.A1(fract_denorm[40]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[39]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_86));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4411 (.A1(fract_denorm[24]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[23]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_85));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4412 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[47]),
    .B1(u4_sll_315_50_n_29),
    .B2(fract_denorm[46]),
    .Y(u4_sll_315_50_n_84));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4413 (.A1(fract_denorm[34]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[33]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_83));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4414 (.A1(fract_denorm[14]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[13]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_82));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4415 (.A1(fract_denorm[36]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[35]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_81));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4416 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[17]),
    .B1(n_3819),
    .B2(fract_denorm[16]),
    .Y(u4_sll_315_50_n_80));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4417 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[11]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[10]),
    .Y(u4_sll_315_50_n_79));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4418 (.A(n_3752),
    .B(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_77));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4419 (.A(n_3752),
    .B(u4_sll_315_50_n_36),
    .Y(u4_sll_315_50_n_75));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4420 (.A(u4_sll_315_50_n_37),
    .B(u4_sll_315_50_n_13),
    .Y(u4_sll_315_50_n_73));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4421 (.A(u4_sll_315_50_n_13),
    .B(u4_sll_315_50_n_32),
    .Y(u4_sll_315_50_n_71));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4422 (.A(u4_sll_315_50_n_13),
    .B(u4_sll_315_50_n_33),
    .Y(u4_sll_315_50_n_69));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4423 (.A(u4_sll_315_50_n_13),
    .B(u4_sll_315_50_n_36),
    .Y(u4_sll_315_50_n_68));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4424 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[13]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[12]),
    .Y(u4_sll_315_50_n_66));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4425 (.A1(fract_denorm[10]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[9]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_65));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4426 (.A1(fract_denorm[12]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[11]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_64));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4427 (.A1(fract_denorm[30]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[29]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_63));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4428 (.A1(fract_denorm[16]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[15]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_62));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4429 (.A1(exp_r[0]),
    .A2(fract_denorm[29]),
    .B1(n_3819),
    .B2(fract_denorm[28]),
    .Y(u4_sll_315_50_n_61));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4430 (.A1(fract_denorm[18]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[17]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_60));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4431 (.A1(exp_r[0]),
    .A2(fract_denorm[31]),
    .B1(n_3819),
    .B2(fract_denorm[30]),
    .Y(u4_sll_315_50_n_59));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4432 (.A1(fract_denorm[20]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[19]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_58));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4433 (.A1(fract_denorm[22]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[21]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_57));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4434 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[35]),
    .B1(n_3819),
    .B2(fract_denorm[34]),
    .Y(u4_sll_315_50_n_56));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4435 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[3]),
    .B1(n_3819),
    .B2(fract_denorm[2]),
    .Y(u4_sll_315_50_n_55));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4436 (.A1(fract_denorm[43]),
    .A2(u4_sll_315_50_n_19),
    .B1(fract_denorm[42]),
    .B2(u4_sll_315_50_n_11),
    .Y(u4_sll_315_50_n_54));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4437 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[33]),
    .B1(n_3819),
    .B2(fract_denorm[32]),
    .Y(u4_sll_315_50_n_53));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4438 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[27]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[26]),
    .Y(u4_sll_315_50_n_52));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4439 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[9]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[8]),
    .Y(u4_sll_315_50_n_51));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4440 (.A1(fract_denorm[28]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[27]),
    .B2(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_50));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4441 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[23]),
    .B1(n_3819),
    .B2(fract_denorm[22]),
    .Y(u4_sll_315_50_n_49));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4442 (.A1(exp_r[0]),
    .A2(fract_denorm[19]),
    .B1(n_3819),
    .B2(fract_denorm[18]),
    .Y(u4_sll_315_50_n_48));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4443 (.A1(fract_denorm[15]),
    .A2(u4_sll_315_50_n_19),
    .B1(fract_denorm[14]),
    .B2(u4_sll_315_50_n_11),
    .Y(u4_sll_315_50_n_47));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4444 (.A1(fract_denorm[32]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[31]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_46));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4445 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[39]),
    .B1(u4_sll_315_50_n_10),
    .B2(fract_denorm[38]),
    .Y(u4_sll_315_50_n_45));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4446 (.A1(fract_denorm[42]),
    .A2(u4_sll_315_50_n_9),
    .B1(fract_denorm[41]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_44));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4447 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[45]),
    .B1(u4_sll_315_50_n_29),
    .B2(fract_denorm[44]),
    .Y(u4_sll_315_50_n_43));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4448 (.A1(fract_denorm[38]),
    .A2(u4_sll_315_50_n_7),
    .B1(fract_denorm[37]),
    .B2(u4_sll_315_50_n_8),
    .Y(u4_sll_315_50_n_42));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4449 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[21]),
    .B1(n_3819),
    .B2(fract_denorm[20]),
    .Y(u4_sll_315_50_n_41));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4450 (.A1(u4_sll_315_50_n_18),
    .A2(fract_denorm[37]),
    .B1(u4_sll_315_50_n_10),
    .B2(fract_denorm[36]),
    .Y(u4_sll_315_50_n_40));
 AOI22xp33_ASAP7_75t_R u4_sll_315_50_g4451 (.A1(u4_sll_315_50_n_19),
    .A2(fract_denorm[1]),
    .B1(u4_sll_315_50_n_11),
    .B2(fract_denorm[0]),
    .Y(u4_sll_315_50_n_39));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4452 (.A(fract_denorm[0]),
    .B(u4_sll_315_50_n_7),
    .Y(u4_sll_315_50_n_38));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4453 (.A(u4_sll_315_50_n_14),
    .B(n_3824),
    .Y(u4_sll_315_50_n_37));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4454 (.A(n_3751),
    .B(n_3483),
    .Y(u4_sll_315_50_n_36));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4455 (.A(fract_denorm[47]),
    .B(u4_sll_315_50_n_2),
    .Y(u4_sll_315_50_n_35));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4456 (.A(fract_denorm[47]),
    .B(u4_sll_315_50_n_30),
    .Y(u4_sll_315_50_n_34));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4457 (.A(n_3751),
    .B(n_3824),
    .Y(u4_sll_315_50_n_33));
 NOR2xp33_ASAP7_75t_R u4_sll_315_50_g4458 (.A(n_3483),
    .B(u4_sll_315_50_n_14),
    .Y(u4_sll_315_50_n_32));
 NAND2xp33_ASAP7_75t_R u4_sll_315_50_g4459 (.A(n_3752),
    .B(u4_sll_315_50_n_30),
    .Y(u4_sll_315_50_n_31));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4460 (.A(n_3753),
    .Y(u4_sll_315_50_n_30));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4466 (.A(n_3819),
    .Y(u4_sll_315_50_n_19));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4473 (.A(u4_sll_315_50_n_11),
    .Y(u4_sll_315_50_n_18));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4482 (.A(u4_sll_315_50_n_10),
    .Y(u4_sll_315_50_n_9));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4485 (.A(u4_sll_315_50_n_7),
    .Y(u4_sll_315_50_n_10));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4486 (.A(n_3819),
    .Y(u4_sll_315_50_n_7));
 HB1xp67_ASAP7_75t_R u4_sll_315_50_g4490 (.A(u4_sll_315_50_n_17),
    .Y(u4_sll_315_50_n_16));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4500 (.A(u4_sll_315_50_n_3),
    .Y(u4_sll_315_50_n_4));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4519 (.A(u4_sll_315_50_n_17),
    .Y(u4_sll_315_50_n_2));
 HB1xp67_ASAP7_75t_R u4_sll_315_50_g4530 (.A(u4_sll_315_50_n_1),
    .Y(u4_sll_315_50_n_17));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4542 (.A(n_3751),
    .Y(u4_sll_315_50_n_14));
 INVxp33_ASAP7_75t_R u4_sll_315_50_g4543 (.A(n_3752),
    .Y(u4_sll_315_50_n_13));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29153 (.A(u5_mul_69_18_n_41),
    .Y(u5_mul_69_18_n_39));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29154 (.A(u5_mul_69_18_n_74),
    .Y(u5_mul_69_18_n_41));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29161 (.A(u5_mul_69_18_n_139),
    .Y(u5_mul_69_18_n_65));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29167 (.A(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_38));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29168 (.A(u5_mul_69_18_n_87),
    .Y(u5_mul_69_18_n_47));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29174 (.A(u5_mul_69_18_n_62),
    .Y(u5_mul_69_18_n_37));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29175 (.A(u5_mul_69_18_n_134),
    .Y(u5_mul_69_18_n_62));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29181 (.A(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_36));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29182 (.A(u5_mul_69_18_n_79),
    .Y(u5_mul_69_18_n_43));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29189 (.A(u5_mul_69_18_n_129),
    .Y(u5_mul_69_18_n_60));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29196 (.A(u5_mul_69_18_n_123),
    .Y(u5_mul_69_18_n_57));
 INVxp33_ASAP7_75t_R u5_mul_69_18_drc_bufs29203 (.A(u5_mul_69_18_n_99),
    .Y(u5_mul_69_18_n_52));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29226 (.A(u5_mul_69_18_n_151),
    .Y(u5_mul_69_18_n_35));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29244 (.A(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_34));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29297 (.A(u5_mul_69_18_n_149),
    .Y(u5_mul_69_18_n_33));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29315 (.A(u5_mul_69_18_n_633),
    .Y(u5_mul_69_18_n_32));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29363 (.A(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_31));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29369 (.A(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_30));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29375 (.A(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_29));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_drc_bufs29411 (.A(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_28));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g2 (.A(u5_mul_69_18_n_1854),
    .B(n_14301),
    .Y(u5_mul_69_18_n_27));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26791 (.A1(u5_mul_69_18_n_1577),
    .A2(u5_mul_69_18_n_2034),
    .B(u5_mul_69_18_n_1599),
    .Y(u5_mul_69_18_n_2036));
 OA21x2_ASAP7_75t_R u5_mul_69_18_g26793 (.A1(u5_mul_69_18_n_1626),
    .A2(u5_mul_69_18_n_2032),
    .B(u5_mul_69_18_n_1643),
    .Y(u5_mul_69_18_n_2034));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26795 (.A1(u5_mul_69_18_n_2030),
    .A2(u5_mul_69_18_n_1679),
    .B(u5_mul_69_18_n_1686),
    .Y(u5_mul_69_18_n_2032));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26797 (.A1(u5_mul_69_18_n_1714),
    .A2(u5_mul_69_18_n_2028),
    .B(u5_mul_69_18_n_1735),
    .Y(u5_mul_69_18_n_2030));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26799 (.A1(u5_mul_69_18_n_1760),
    .A2(u5_mul_69_18_n_2026),
    .B(u5_mul_69_18_n_1770),
    .Y(u5_mul_69_18_n_2028));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26801 (.A1(u5_mul_69_18_n_1798),
    .A2(u5_mul_69_18_n_2024),
    .B(u5_mul_69_18_n_1812),
    .Y(u5_mul_69_18_n_2026));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26803 (.A1(u5_mul_69_18_n_1797),
    .A2(u5_mul_69_18_n_2022),
    .B(u5_mul_69_18_n_1810),
    .Y(u5_mul_69_18_n_2024));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26805 (.A1(u5_mul_69_18_n_1832),
    .A2(u5_mul_69_18_n_2020),
    .B(u5_mul_69_18_n_1839),
    .Y(u5_mul_69_18_n_2022));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26807 (.A1(u5_mul_69_18_n_2018),
    .A2(u5_mul_69_18_n_1836),
    .B(u5_mul_69_18_n_23),
    .Y(u5_mul_69_18_n_2020));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26809 (.A1(u5_mul_69_18_n_1857),
    .A2(u5_mul_69_18_n_2016),
    .B(u5_mul_69_18_n_1869),
    .Y(u5_mul_69_18_n_2018));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26811 (.A1(u5_mul_69_18_n_2014),
    .A2(u5_mul_69_18_n_1888),
    .B(u5_mul_69_18_n_25),
    .Y(u5_mul_69_18_n_2016));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26813 (.A1(u5_mul_69_18_n_1912),
    .A2(u5_mul_69_18_n_2012),
    .B(u5_mul_69_18_n_1919),
    .Y(u5_mul_69_18_n_2014));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26815 (.A1(u5_mul_69_18_n_2010),
    .A2(u5_mul_69_18_n_1917),
    .B(u5_mul_69_18_n_26),
    .Y(u5_mul_69_18_n_2012));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26817 (.A1(u5_mul_69_18_n_1934),
    .A2(u5_mul_69_18_n_2008),
    .B(u5_mul_69_18_n_1943),
    .Y(u5_mul_69_18_n_2010));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26819 (.A1(u5_mul_69_18_n_1921),
    .A2(u5_mul_69_18_n_2006),
    .B(u5_mul_69_18_n_1929),
    .Y(u5_mul_69_18_n_2008));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26821 (.A1(u5_mul_69_18_n_1940),
    .A2(u5_mul_69_18_n_2004),
    .B(u5_mul_69_18_n_1938),
    .Y(u5_mul_69_18_n_2006));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26823 (.A1(u5_mul_69_18_n_2002),
    .A2(u5_mul_69_18_n_1932),
    .B(u5_mul_69_18_n_1941),
    .Y(u5_mul_69_18_n_2004));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26825 (.A1(u5_mul_69_18_n_1944),
    .A2(u5_mul_69_18_n_2000),
    .B(u5_mul_69_18_n_1958),
    .Y(u5_mul_69_18_n_2002));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26827 (.A1(u5_mul_69_18_n_1945),
    .A2(u5_mul_69_18_n_1998),
    .B(u5_mul_69_18_n_1950),
    .Y(u5_mul_69_18_n_2000));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26829 (.A1(u5_mul_69_18_n_1996),
    .A2(u5_mul_69_18_n_1961),
    .B(u5_mul_69_18_n_1962),
    .Y(u5_mul_69_18_n_1998));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26831 (.A1(u5_mul_69_18_n_1956),
    .A2(u5_mul_69_18_n_1994),
    .B(u5_mul_69_18_n_1957),
    .Y(u5_mul_69_18_n_1996));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26833 (.A1(u5_mul_69_18_n_1922),
    .A2(u5_mul_69_18_n_1992),
    .B(u5_mul_69_18_n_1930),
    .Y(u5_mul_69_18_n_1994));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26835 (.A1(u5_mul_69_18_n_1936),
    .A2(u5_mul_69_18_n_1990),
    .B(u5_mul_69_18_n_1942),
    .Y(u5_mul_69_18_n_1992));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26837 (.A1(u5_mul_69_18_n_1988),
    .A2(u5_mul_69_18_n_1915),
    .B(u5_mul_69_18_n_27),
    .Y(u5_mul_69_18_n_1990));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26839 (.A1(u5_mul_69_18_n_1907),
    .A2(u5_mul_69_18_n_1986),
    .B(u5_mul_69_18_n_1913),
    .Y(u5_mul_69_18_n_1988));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26841 (.A1(u5_mul_69_18_n_1911),
    .A2(u5_mul_69_18_n_1984),
    .B(u5_mul_69_18_n_1918),
    .Y(u5_mul_69_18_n_1986));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26843 (.A1(u5_mul_69_18_n_1884),
    .A2(u5_mul_69_18_n_1982),
    .B(u5_mul_69_18_n_1889),
    .Y(u5_mul_69_18_n_1984));
 AO21x1_ASAP7_75t_R u5_mul_69_18_g26845 (.A1(u5_mul_69_18_n_1885),
    .A2(u5_mul_69_18_n_1980),
    .B(u5_mul_69_18_n_1890),
    .Y(u5_mul_69_18_n_1982));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26847 (.A1(u5_mul_69_18_n_1867),
    .A2(u5_mul_69_18_n_1978),
    .B(u5_mul_69_18_n_24),
    .Y(u5_mul_69_18_n_1980));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26849 (.A1(u5_mul_69_18_n_1976),
    .A2(u5_mul_69_18_n_1860),
    .B(u5_mul_69_18_n_1868),
    .Y(u5_mul_69_18_n_1978));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26851 (.A1(u5_mul_69_18_n_1838),
    .A2(u5_mul_69_18_n_1974),
    .B(u5_mul_69_18_n_22),
    .Y(u5_mul_69_18_n_1976));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26853 (.A1(u5_mul_69_18_n_1972),
    .A2(u5_mul_69_18_n_1804),
    .B(u5_mul_69_18_n_1811),
    .Y(u5_mul_69_18_n_1974));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26855 (.A1(u5_mul_69_18_n_1799),
    .A2(u5_mul_69_18_n_1970),
    .B(u5_mul_69_18_n_1809),
    .Y(u5_mul_69_18_n_1972));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26857 (.A1(u5_mul_69_18_n_1968),
    .A2(u5_mul_69_18_n_1774),
    .B(u5_mul_69_18_n_20),
    .Y(u5_mul_69_18_n_1970));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26859 (.A1(u5_mul_69_18_n_1759),
    .A2(u5_mul_69_18_n_1965),
    .B(u5_mul_69_18_n_1775),
    .Y(u5_mul_69_18_n_1968));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26861 (.A1(u5_mul_69_18_n_1951),
    .A2(u5_mul_69_18_n_1925),
    .B(u5_mul_69_18_n_1962),
    .Y(u5_mul_69_18_n_1966));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26862 (.A1(u5_mul_69_18_n_1772),
    .A2(u5_mul_69_18_n_1949),
    .B(u5_mul_69_18_n_19),
    .Y(u5_mul_69_18_n_1965));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26864 (.A1(u5_mul_69_18_n_1926),
    .A2(u5_mul_69_18_n_1931),
    .B(u5_mul_69_18_n_1957),
    .Y(u5_mul_69_18_n_1963));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26865 (.A(u5_mul_69_18_n_1925),
    .B(u5_mul_69_18_n_1951),
    .Y(u5_mul_69_18_n_1962));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26866 (.A(u5_mul_69_18_n_1925),
    .B(u5_mul_69_18_n_1951),
    .Y(u5_mul_69_18_n_1961));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26867 (.A1(n_14298),
    .A2(u5_mul_69_18_n_1895),
    .B(u5_mul_69_18_n_1958),
    .Y(u5_mul_69_18_n_1960));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26868 (.A1(u5_mul_69_18_n_1924),
    .A2(n_14299),
    .B(u5_mul_69_18_n_1950),
    .Y(u5_mul_69_18_n_1959));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26869 (.A(u5_mul_69_18_n_1895),
    .B(n_14298),
    .Y(u5_mul_69_18_n_1958));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26870 (.A(u5_mul_69_18_n_1931),
    .B(u5_mul_69_18_n_1926),
    .Y(u5_mul_69_18_n_1956));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26871 (.A1(u5_mul_69_18_n_1876),
    .A2(n_14300),
    .B(u5_mul_69_18_n_1943),
    .Y(u5_mul_69_18_n_1955));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26872 (.A1(u5_mul_69_18_n_1899),
    .A2(u5_mul_69_18_n_1900),
    .B(u5_mul_69_18_n_1942),
    .Y(u5_mul_69_18_n_1954));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26873 (.A1(u5_mul_69_18_n_1898),
    .A2(u5_mul_69_18_n_1903),
    .B(u5_mul_69_18_n_1941),
    .Y(u5_mul_69_18_n_1953));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26874 (.A1(u5_mul_69_18_n_1902),
    .A2(u5_mul_69_18_n_1874),
    .B(u5_mul_69_18_n_1930),
    .Y(u5_mul_69_18_n_1952));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26875 (.A(u5_mul_69_18_n_1931),
    .B(u5_mul_69_18_n_1926),
    .Y(u5_mul_69_18_n_1957));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26877 (.A1(u5_mul_69_18_n_1901),
    .A2(u5_mul_69_18_n_1873),
    .B(u5_mul_69_18_n_1929),
    .Y(u5_mul_69_18_n_1947));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26878 (.A(u5_mul_69_18_n_1939),
    .B(u5_mul_69_18_n_1938),
    .Y(u5_mul_69_18_n_1946));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26879 (.A(u5_mul_69_18_n_1924),
    .B(n_14299),
    .Y(u5_mul_69_18_n_1945));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26880 (.A(u5_mul_69_18_n_1895),
    .B(n_14298),
    .Y(u5_mul_69_18_n_1944));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26881 (.A(u5_mul_69_18_n_1891),
    .B(u5_mul_69_18_n_1820),
    .Y(u5_mul_69_18_n_1951));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26882 (.A(u5_mul_69_18_n_1924),
    .B(n_14299),
    .Y(u5_mul_69_18_n_1950));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26883 (.A1(u5_mul_69_18_n_1687),
    .A2(u5_mul_69_18_n_1894),
    .B(u5_mul_69_18_n_1673),
    .Y(u5_mul_69_18_n_1949));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26884 (.A(u5_mul_69_18_n_1939),
    .Y(u5_mul_69_18_n_1940));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26885 (.A1(n_14305),
    .A2(u5_mul_69_18_n_1848),
    .B(u5_mul_69_18_n_1918),
    .Y(u5_mul_69_18_n_1937));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26886 (.A(u5_mul_69_18_n_1876),
    .B(n_14300),
    .Y(u5_mul_69_18_n_1943));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26887 (.A(u5_mul_69_18_n_1899),
    .B(u5_mul_69_18_n_1900),
    .Y(u5_mul_69_18_n_1936));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26888 (.A(u5_mul_69_18_n_1899),
    .B(u5_mul_69_18_n_1900),
    .Y(u5_mul_69_18_n_1942));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26889 (.A1(u5_mul_69_18_n_1852),
    .A2(n_14304),
    .B(u5_mul_69_18_n_1919),
    .Y(u5_mul_69_18_n_1935));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26890 (.A(u5_mul_69_18_n_1876),
    .B(n_14300),
    .Y(u5_mul_69_18_n_1934));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26891 (.A(u5_mul_69_18_n_1916),
    .B(u5_mul_69_18_n_26),
    .Y(u5_mul_69_18_n_1933));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26892 (.A(u5_mul_69_18_n_1903),
    .B(u5_mul_69_18_n_1898),
    .Y(u5_mul_69_18_n_1941));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26893 (.A(u5_mul_69_18_n_1903),
    .B(u5_mul_69_18_n_1898),
    .Y(u5_mul_69_18_n_1932));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26894 (.A(u5_mul_69_18_n_1905),
    .B(u5_mul_69_18_n_1897),
    .Y(u5_mul_69_18_n_1939));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26895 (.A(u5_mul_69_18_n_1896),
    .B(u5_mul_69_18_n_1906),
    .Y(u5_mul_69_18_n_1938));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26896 (.A(u5_mul_69_18_n_1872),
    .B(n_14308),
    .Y(u5_mul_69_18_n_1931));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26897 (.A1(u5_mul_69_18_n_1847),
    .A2(n_14302),
    .B(u5_mul_69_18_n_1913),
    .Y(u5_mul_69_18_n_1923));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26898 (.A(u5_mul_69_18_n_1874),
    .B(u5_mul_69_18_n_1902),
    .Y(u5_mul_69_18_n_1930));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26899 (.A(u5_mul_69_18_n_1874),
    .B(u5_mul_69_18_n_1902),
    .Y(u5_mul_69_18_n_1922));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26900 (.A(u5_mul_69_18_n_1873),
    .B(u5_mul_69_18_n_1901),
    .Y(u5_mul_69_18_n_1929));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26901 (.A(u5_mul_69_18_n_1873),
    .B(u5_mul_69_18_n_1901),
    .Y(u5_mul_69_18_n_1921));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26902 (.A(u5_mul_69_18_n_1914),
    .B(u5_mul_69_18_n_27),
    .Y(u5_mul_69_18_n_1920));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26905 (.A(n_14307),
    .B(n_14323),
    .C(u5_mul_69_18_n_1787),
    .Y(u5_mul_69_18_n_1926));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26906 (.A(n_14308),
    .B(u5_mul_69_18_n_1743),
    .C(u5_mul_69_18_n_1819),
    .Y(u5_mul_69_18_n_1925));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26907 (.A(n_14310),
    .B(n_14322),
    .C(u5_mul_69_18_n_1820),
    .Y(u5_mul_69_18_n_1924));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26908 (.A(u5_mul_69_18_n_1916),
    .Y(u5_mul_69_18_n_1917));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26909 (.A(u5_mul_69_18_n_1914),
    .Y(u5_mul_69_18_n_1915));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26910 (.A(u5_mul_69_18_n_1852),
    .B(n_14304),
    .Y(u5_mul_69_18_n_1912));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26911 (.A(u5_mul_69_18_n_1852),
    .B(n_14304),
    .Y(u5_mul_69_18_n_1919));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26912 (.A(u5_mul_69_18_n_1848),
    .B(n_14305),
    .Y(u5_mul_69_18_n_1911));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26913 (.A(u5_mul_69_18_n_1848),
    .B(n_14305),
    .Y(u5_mul_69_18_n_1918));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26914 (.A(u5_mul_69_18_n_1887),
    .B(u5_mul_69_18_n_25),
    .Y(u5_mul_69_18_n_1910));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26915 (.A1(u5_mul_69_18_n_1850),
    .A2(n_14461),
    .B(u5_mul_69_18_n_1889),
    .Y(u5_mul_69_18_n_1909));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26916 (.A1(u5_mul_69_18_n_1851),
    .A2(n_14309),
    .B(u5_mul_69_18_n_1890),
    .Y(u5_mul_69_18_n_1908));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26917 (.A(n_14303),
    .B(u5_mul_69_18_n_1875),
    .Y(u5_mul_69_18_n_1916));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26919 (.A(u5_mul_69_18_n_1854),
    .B(n_14301),
    .Y(u5_mul_69_18_n_1914));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26921 (.A(u5_mul_69_18_n_1847),
    .B(n_14302),
    .Y(u5_mul_69_18_n_1907));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26922 (.A(u5_mul_69_18_n_1847),
    .B(n_14302),
    .Y(u5_mul_69_18_n_1913));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26923 (.A(u5_mul_69_18_n_1905),
    .Y(u5_mul_69_18_n_1906));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26924 (.A(u5_mul_69_18_n_1896),
    .Y(u5_mul_69_18_n_1897));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26925 (.A(u5_mul_69_18_n_1893),
    .Y(u5_mul_69_18_n_1894));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g26927 (.A(u5_mul_69_18_n_1840),
    .B(u5_mul_69_18_n_1784),
    .Y(u5_mul_69_18_n_1905));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26929 (.A(u5_mul_69_18_n_1843),
    .B(u5_mul_69_18_n_1846),
    .Y(u5_mul_69_18_n_1903));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26930 (.A(n_14310),
    .B(n_14322),
    .Y(u5_mul_69_18_n_1891));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26931 (.A(n_14307),
    .B(u5_mul_69_18_n_1844),
    .Y(u5_mul_69_18_n_1902));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26932 (.A(u5_mul_69_18_n_1842),
    .B(u5_mul_69_18_n_1786),
    .Y(u5_mul_69_18_n_1901));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26933 (.A(u5_mul_69_18_n_1841),
    .B(u5_mul_69_18_n_1785),
    .Y(u5_mul_69_18_n_1900));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26934 (.A(u5_mul_69_18_n_1833),
    .B(n_14341),
    .C(u5_mul_69_18_n_1748),
    .Y(u5_mul_69_18_n_1899));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26935 (.A(u5_mul_69_18_n_1817),
    .B(u5_mul_69_18_n_1694),
    .C(u5_mul_69_18_n_1788),
    .Y(u5_mul_69_18_n_1898));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26936 (.A(u5_mul_69_18_n_1846),
    .B(u5_mul_69_18_n_1691),
    .C(n_14462),
    .Y(u5_mul_69_18_n_1896));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g26937 (.A(u5_mul_69_18_n_1821),
    .B(n_14325),
    .C(u5_mul_69_18_n_1818),
    .Y(u5_mul_69_18_n_1895));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26938 (.A1(u5_mul_69_18_n_1632),
    .A2(u5_mul_69_18_n_1864),
    .B(u5_mul_69_18_n_1642),
    .Y(u5_mul_69_18_n_1893));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26939 (.A(u5_mul_69_18_n_1887),
    .Y(u5_mul_69_18_n_1888));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26941 (.A(n_14309),
    .B(u5_mul_69_18_n_1851),
    .Y(u5_mul_69_18_n_1890));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26942 (.A(u5_mul_69_18_n_1851),
    .B(n_14309),
    .Y(u5_mul_69_18_n_1885));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26943 (.A(u5_mul_69_18_n_1850),
    .B(n_14461),
    .Y(u5_mul_69_18_n_1884));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26944 (.A(n_14461),
    .B(u5_mul_69_18_n_1850),
    .Y(u5_mul_69_18_n_1889));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26945 (.A1(n_14313),
    .A2(u5_mul_69_18_n_1823),
    .B(u5_mul_69_18_n_1869),
    .Y(u5_mul_69_18_n_1883));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26947 (.A(u5_mul_69_18_n_1849),
    .B(n_14306),
    .Y(u5_mul_69_18_n_1887));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26948 (.A1(u5_mul_69_18_n_1822),
    .A2(n_14311),
    .B(u5_mul_69_18_n_1868),
    .Y(u5_mul_69_18_n_1882));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26949 (.A(u5_mul_69_18_n_1866),
    .B(u5_mul_69_18_n_24),
    .Y(u5_mul_69_18_n_1881));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26953 (.A(u5_mul_69_18_n_1819),
    .B(u5_mul_69_18_n_1743),
    .Y(u5_mul_69_18_n_1872));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26960 (.A(u5_mul_69_18_n_1786),
    .B(n_14339),
    .C(u5_mul_69_18_n_1782),
    .Y(u5_mul_69_18_n_1876));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26961 (.A(u5_mul_69_18_n_1806),
    .B(n_14340),
    .C(u5_mul_69_18_n_1790),
    .Y(u5_mul_69_18_n_1875));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26962 (.A(u5_mul_69_18_n_1780),
    .B(n_14324),
    .C(u5_mul_69_18_n_1785),
    .Y(u5_mul_69_18_n_1874));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g26963 (.A(u5_mul_69_18_n_1784),
    .B(n_14331),
    .C(n_14317),
    .Y(u5_mul_69_18_n_1873));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26964 (.A(u5_mul_69_18_n_1866),
    .Y(u5_mul_69_18_n_1867));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26967 (.A(n_14313),
    .B(u5_mul_69_18_n_1823),
    .Y(u5_mul_69_18_n_1869));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26968 (.A(n_14311),
    .B(u5_mul_69_18_n_1822),
    .Y(u5_mul_69_18_n_1860));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26969 (.A(n_14311),
    .B(u5_mul_69_18_n_1822),
    .Y(u5_mul_69_18_n_1868));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g26970 (.A1(u5_mul_69_18_n_1752),
    .A2(n_14314),
    .B(u5_mul_69_18_n_1839),
    .Y(u5_mul_69_18_n_1859));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26971 (.A(u5_mul_69_18_n_1837),
    .B(u5_mul_69_18_n_22),
    .Y(u5_mul_69_18_n_1858));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26973 (.A(n_14313),
    .B(u5_mul_69_18_n_1823),
    .Y(u5_mul_69_18_n_1857));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g26974 (.A(u5_mul_69_18_n_1835),
    .B(u5_mul_69_18_n_23),
    .Y(u5_mul_69_18_n_1856));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g26975 (.A(u5_mul_69_18_n_1826),
    .B(n_14312),
    .Y(u5_mul_69_18_n_1866));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g26978 (.A1(u5_mul_69_18_n_1808),
    .A2(u5_mul_69_18_n_1601),
    .B(u5_mul_69_18_n_1578),
    .Y(u5_mul_69_18_n_1864));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26983 (.A(n_14330),
    .B(n_14334),
    .C(u5_mul_69_18_n_1749),
    .Y(u5_mul_69_18_n_1854));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26984 (.A(u5_mul_69_18_n_1787),
    .B(n_14323),
    .Y(u5_mul_69_18_n_1844));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26987 (.A(n_14462),
    .B(u5_mul_69_18_n_1691),
    .Y(u5_mul_69_18_n_1843));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26988 (.A(u5_mul_69_18_n_1782),
    .B(n_14339),
    .Y(u5_mul_69_18_n_1842));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g26989 (.A(u5_mul_69_18_n_1780),
    .B(n_14324),
    .Y(u5_mul_69_18_n_1841));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g26990 (.A(n_14317),
    .B(n_14331),
    .Y(u5_mul_69_18_n_1840));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26991 (.A(u5_mul_69_18_n_1789),
    .B(u5_mul_69_18_n_1688),
    .C(n_14320),
    .Y(u5_mul_69_18_n_1852));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26992 (.A(u5_mul_69_18_n_1746),
    .B(n_14365),
    .C(u5_mul_69_18_n_1657),
    .Y(u5_mul_69_18_n_1851));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26993 (.A(n_14329),
    .B(n_14345),
    .C(u5_mul_69_18_n_1703),
    .Y(u5_mul_69_18_n_1850));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26994 (.A(u5_mul_69_18_n_1750),
    .B(u5_mul_69_18_n_1639),
    .C(n_14319),
    .Y(u5_mul_69_18_n_1849));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26995 (.A(n_14328),
    .B(u5_mul_69_18_n_1616),
    .C(u5_mul_69_18_n_1705),
    .Y(u5_mul_69_18_n_1848));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g26996 (.A(u5_mul_69_18_n_1783),
    .B(n_14338),
    .C(u5_mul_69_18_n_1745),
    .Y(u5_mul_69_18_n_1847));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g26997 (.A(n_14321),
    .B(u5_mul_69_18_n_1617),
    .C(n_14463),
    .Y(u5_mul_69_18_n_1846));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g26999 (.A(u5_mul_69_18_n_1837),
    .Y(u5_mul_69_18_n_1838));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27000 (.A(u5_mul_69_18_n_1835),
    .Y(u5_mul_69_18_n_1836));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27001 (.A(u5_mul_69_18_n_1752),
    .B(n_14314),
    .Y(u5_mul_69_18_n_1839));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27002 (.A(u5_mul_69_18_n_1752),
    .B(n_14314),
    .Y(u5_mul_69_18_n_1832));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27003 (.A1(n_14326),
    .A2(u5_mul_69_18_n_1710),
    .B(u5_mul_69_18_n_1812),
    .Y(u5_mul_69_18_n_1831));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27004 (.A1(n_14327),
    .A2(u5_mul_69_18_n_1709),
    .B(u5_mul_69_18_n_1811),
    .Y(u5_mul_69_18_n_1830));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27006 (.A(u5_mul_69_18_n_1753),
    .B(n_14315),
    .Y(u5_mul_69_18_n_1837));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27008 (.A(u5_mul_69_18_n_1794),
    .B(n_14316),
    .Y(u5_mul_69_18_n_1835));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27009 (.A1(u5_mul_69_18_n_1712),
    .A2(u5_mul_69_18_n_1756),
    .B(u5_mul_69_18_n_1809),
    .Y(u5_mul_69_18_n_1829));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27010 (.A1(u5_mul_69_18_n_1754),
    .A2(n_14318),
    .B(u5_mul_69_18_n_1810),
    .Y(u5_mul_69_18_n_1828));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27013 (.A(u5_mul_69_18_n_1738),
    .B(u5_mul_69_18_n_1662),
    .Y(u5_mul_69_18_n_1833));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27016 (.A(n_14337),
    .B(n_14366),
    .C(u5_mul_69_18_n_1659),
    .Y(u5_mul_69_18_n_1826));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27022 (.A(n_14336),
    .B(n_14358),
    .C(u5_mul_69_18_n_1707),
    .Y(u5_mul_69_18_n_1823));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27023 (.A(u5_mul_69_18_n_1695),
    .B(u5_mul_69_18_n_1566),
    .C(u5_mul_69_18_n_1554),
    .Y(u5_mul_69_18_n_1822));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27025 (.A(u5_mul_69_18_n_1689),
    .B(u5_mul_69_18_n_1652),
    .C(u5_mul_69_18_n_1696),
    .Y(u5_mul_69_18_n_1821));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27026 (.A(u5_mul_69_18_n_1693),
    .B(u5_mul_69_18_n_1660),
    .C(u5_mul_69_18_n_1731),
    .Y(u5_mul_69_18_n_1820));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27027 (.A(n_14335),
    .B(u5_mul_69_18_n_1581),
    .C(u5_mul_69_18_n_1697),
    .Y(u5_mul_69_18_n_1819));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27028 (.A(u5_mul_69_18_n_1739),
    .B(u5_mul_69_18_n_1706),
    .Y(u5_mul_69_18_n_1818));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27029 (.A(n_14321),
    .B(u5_mul_69_18_n_1716),
    .Y(u5_mul_69_18_n_1817));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27030 (.A(u5_mul_69_18_n_1807),
    .Y(u5_mul_69_18_n_1808));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27032 (.A(u5_mul_69_18_n_1710),
    .B(n_14326),
    .Y(u5_mul_69_18_n_1812));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27033 (.A(u5_mul_69_18_n_1709),
    .B(n_14327),
    .Y(u5_mul_69_18_n_1811));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27034 (.A(u5_mul_69_18_n_1709),
    .B(n_14327),
    .Y(u5_mul_69_18_n_1804));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27035 (.A1(u5_mul_69_18_n_1711),
    .A2(n_14333),
    .B(u5_mul_69_18_n_1770),
    .Y(u5_mul_69_18_n_1803));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27036 (.A1(u5_mul_69_18_n_1665),
    .A2(u5_mul_69_18_n_1713),
    .B(u5_mul_69_18_n_1775),
    .Y(u5_mul_69_18_n_1802));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27037 (.A(u5_mul_69_18_n_1773),
    .B(u5_mul_69_18_n_20),
    .Y(u5_mul_69_18_n_1801));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27038 (.A(u5_mul_69_18_n_1771),
    .B(u5_mul_69_18_n_19),
    .Y(u5_mul_69_18_n_1800));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27039 (.A(u5_mul_69_18_n_1712),
    .B(u5_mul_69_18_n_1756),
    .Y(u5_mul_69_18_n_1799));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27040 (.A(n_14326),
    .B(u5_mul_69_18_n_1710),
    .Y(u5_mul_69_18_n_1798));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27041 (.A(n_14318),
    .B(u5_mul_69_18_n_1754),
    .Y(u5_mul_69_18_n_1797));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27042 (.A(n_14318),
    .B(u5_mul_69_18_n_1754),
    .Y(u5_mul_69_18_n_1810));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27045 (.A(u5_mul_69_18_n_1712),
    .B(u5_mul_69_18_n_1756),
    .Y(u5_mul_69_18_n_1809));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27046 (.A1(u5_mul_69_18_n_1733),
    .A2(u5_mul_69_18_n_1538),
    .B(u5_mul_69_18_n_1503),
    .Y(u5_mul_69_18_n_1807));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27048 (.A(u5_mul_69_18_n_1701),
    .B(u5_mul_69_18_n_1624),
    .Y(u5_mul_69_18_n_1806));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27053 (.A(u5_mul_69_18_n_1658),
    .B(n_14353),
    .C(n_14343),
    .Y(u5_mul_69_18_n_1794));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27060 (.A(u5_mul_69_18_n_1699),
    .B(n_14355),
    .C(u5_mul_69_18_n_1561),
    .Y(u5_mul_69_18_n_1790));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27061 (.A(u5_mul_69_18_n_1702),
    .B(u5_mul_69_18_n_1517),
    .C(n_14386),
    .Y(u5_mul_69_18_n_1789));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27062 (.A(u5_mul_69_18_n_1706),
    .B(u5_mul_69_18_n_1653),
    .C(u5_mul_69_18_n_1655),
    .Y(u5_mul_69_18_n_1788));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27063 (.A(u5_mul_69_18_n_1704),
    .B(u5_mul_69_18_n_1612),
    .C(n_14349),
    .Y(u5_mul_69_18_n_1787));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27064 (.A(u5_mul_69_18_n_1654),
    .B(u5_mul_69_18_n_1594),
    .C(u5_mul_69_18_n_1620),
    .Y(u5_mul_69_18_n_1786));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27065 (.A(u5_mul_69_18_n_1682),
    .B(u5_mul_69_18_n_1472),
    .C(u5_mul_69_18_n_1662),
    .Y(u5_mul_69_18_n_1785));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27066 (.A(u5_mul_69_18_n_1700),
    .B(u5_mul_69_18_n_1614),
    .C(n_14347),
    .Y(u5_mul_69_18_n_1784));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27067 (.A(u5_mul_69_18_n_1684),
    .B(u5_mul_69_18_n_1485),
    .C(u5_mul_69_18_n_1560),
    .Y(u5_mul_69_18_n_1783));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27068 (.A(u5_mul_69_18_n_1698),
    .B(u5_mul_69_18_n_1669),
    .Y(u5_mul_69_18_n_1782));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27070 (.A(u5_mul_69_18_n_1704),
    .B(u5_mul_69_18_n_1719),
    .Y(u5_mul_69_18_n_1780));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27071 (.A(u5_mul_69_18_n_1773),
    .Y(u5_mul_69_18_n_1774));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27072 (.A(u5_mul_69_18_n_1771),
    .Y(u5_mul_69_18_n_1772));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27074 (.A(u5_mul_69_18_n_1711),
    .B(n_14333),
    .Y(u5_mul_69_18_n_1760));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27075 (.A(u5_mul_69_18_n_1665),
    .B(u5_mul_69_18_n_1713),
    .Y(u5_mul_69_18_n_1775));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27076 (.A(u5_mul_69_18_n_1665),
    .B(u5_mul_69_18_n_1713),
    .Y(u5_mul_69_18_n_1759));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27077 (.A1(u5_mul_69_18_n_1663),
    .A2(n_14342),
    .B(u5_mul_69_18_n_1735),
    .Y(u5_mul_69_18_n_1758));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27078 (.A(u5_mul_69_18_n_1708),
    .B(u5_mul_69_18_n_1737),
    .Y(u5_mul_69_18_n_1773));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27080 (.A(u5_mul_69_18_n_1664),
    .B(n_14332),
    .Y(u5_mul_69_18_n_1771));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27082 (.A(n_14333),
    .B(u5_mul_69_18_n_1711),
    .Y(u5_mul_69_18_n_1770));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27094 (.A(u5_mul_69_18_n_1677),
    .B(u5_mul_69_18_n_1480),
    .Y(u5_mul_69_18_n_1756));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27097 (.A(u5_mul_69_18_n_1638),
    .B(u5_mul_69_18_n_1473),
    .C(u5_mul_69_18_n_1618),
    .Y(u5_mul_69_18_n_1754));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27098 (.A(u5_mul_69_18_n_1655),
    .B(u5_mul_69_18_n_1653),
    .Y(u5_mul_69_18_n_1739));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27099 (.A(n_14346),
    .B(u5_mul_69_18_n_1567),
    .C(n_14367),
    .Y(u5_mul_69_18_n_1753));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27100 (.A(u5_mul_69_18_n_1621),
    .B(n_14378),
    .C(n_14344),
    .Y(u5_mul_69_18_n_1752));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27102 (.A(u5_mul_69_18_n_1682),
    .B(u5_mul_69_18_n_1472),
    .Y(u5_mul_69_18_n_1738));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27103 (.A(n_14350),
    .B(u5_mul_69_18_n_1494),
    .C(n_14354),
    .Y(u5_mul_69_18_n_1750));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27104 (.A(u5_mul_69_18_n_1661),
    .B(u5_mul_69_18_n_1469),
    .C(n_14356),
    .Y(u5_mul_69_18_n_1749));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27105 (.A(u5_mul_69_18_n_1656),
    .B(n_14370),
    .C(n_14364),
    .Y(u5_mul_69_18_n_1748));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27107 (.A(u5_mul_69_18_n_1649),
    .B(u5_mul_69_18_n_1492),
    .Y(u5_mul_69_18_n_1746));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27108 (.A(u5_mul_69_18_n_1661),
    .B(u5_mul_69_18_n_1668),
    .Y(u5_mul_69_18_n_1745));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27110 (.A(u5_mul_69_18_n_1647),
    .B(u5_mul_69_18_n_1597),
    .Y(u5_mul_69_18_n_1743));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27115 (.A(u5_mul_69_18_n_1732),
    .Y(u5_mul_69_18_n_1733));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27117 (.A1(n_14348),
    .A2(u5_mul_69_18_n_1570),
    .B(u5_mul_69_18_n_1687),
    .Y(u5_mul_69_18_n_1722));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27118 (.A1(u5_mul_69_18_n_1622),
    .A2(u5_mul_69_18_n_1572),
    .B(u5_mul_69_18_n_1686),
    .Y(u5_mul_69_18_n_1721));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27119 (.A(u5_mul_69_18_n_1604),
    .B(n_14360),
    .Y(u5_mul_69_18_n_1737));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27122 (.A(n_14342),
    .B(u5_mul_69_18_n_1663),
    .Y(u5_mul_69_18_n_1735));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27123 (.A(n_14349),
    .B(u5_mul_69_18_n_1612),
    .Y(u5_mul_69_18_n_1719));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27127 (.A(u5_mul_69_18_n_1617),
    .B(n_14463),
    .Y(u5_mul_69_18_n_1716));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27129 (.A(n_14342),
    .B(u5_mul_69_18_n_1663),
    .Y(u5_mul_69_18_n_1714));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27130 (.A1(u5_mul_69_18_n_1641),
    .A2(u5_mul_69_18_n_1452),
    .B(u5_mul_69_18_n_1460),
    .Y(u5_mul_69_18_n_1732));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27131 (.A(u5_mul_69_18_n_1625),
    .B(u5_mul_69_18_n_1471),
    .Y(u5_mul_69_18_n_1731));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27140 (.A(u5_mul_69_18_n_1701),
    .Y(u5_mul_69_18_n_1702));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27142 (.A(u5_mul_69_18_n_1698),
    .Y(u5_mul_69_18_n_1699));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27143 (.A(u5_mul_69_18_n_1692),
    .Y(u5_mul_69_18_n_1693));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27144 (.A(u5_mul_69_18_n_1627),
    .B(u5_mul_69_18_n_1549),
    .Y(u5_mul_69_18_n_1713));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27145 (.A(n_14360),
    .B(u5_mul_69_18_n_1500),
    .C(u5_mul_69_18_n_1527),
    .Y(u5_mul_69_18_n_1712));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27146 (.A(u5_mul_69_18_n_1563),
    .B(u5_mul_69_18_n_1359),
    .C(n_14352),
    .Y(u5_mul_69_18_n_1711));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27147 (.A(u5_mul_69_18_n_1619),
    .B(u5_mul_69_18_n_1467),
    .C(u5_mul_69_18_n_1587),
    .Y(u5_mul_69_18_n_1710));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27148 (.A(n_14359),
    .B(u5_mul_69_18_n_1518),
    .C(u5_mul_69_18_n_1480),
    .Y(u5_mul_69_18_n_1709));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27149 (.A(u5_mul_69_18_n_1550),
    .B(n_14394),
    .C(u5_mul_69_18_n_1489),
    .Y(u5_mul_69_18_n_1708));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27150 (.A(u5_mul_69_18_n_1568),
    .B(u5_mul_69_18_n_1462),
    .C(n_14371),
    .Y(u5_mul_69_18_n_1707));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27151 (.A(n_14464),
    .B(u5_mul_69_18_n_1463),
    .C(n_14363),
    .Y(u5_mul_69_18_n_1706));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27152 (.A(u5_mul_69_18_n_1558),
    .B(n_14384),
    .C(u5_mul_69_18_n_1491),
    .Y(u5_mul_69_18_n_1705));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27153 (.A(u5_mul_69_18_n_1552),
    .B(n_14379),
    .C(u5_mul_69_18_n_1482),
    .Y(u5_mul_69_18_n_1704));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27154 (.A(n_14357),
    .B(u5_mul_69_18_n_1413),
    .C(u5_mul_69_18_n_1493),
    .Y(u5_mul_69_18_n_1703));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27155 (.A(u5_mul_69_18_n_1546),
    .B(u5_mul_69_18_n_1360),
    .C(u5_mul_69_18_n_1486),
    .Y(u5_mul_69_18_n_1701));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27156 (.A(n_14369),
    .B(u5_mul_69_18_n_1497),
    .C(n_14372),
    .Y(u5_mul_69_18_n_1700));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27157 (.A(u5_mul_69_18_n_1591),
    .B(u5_mul_69_18_n_1490),
    .C(u5_mul_69_18_n_1470),
    .Y(u5_mul_69_18_n_1698));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27158 (.A(n_14361),
    .B(u5_mul_69_18_n_1474),
    .C(u5_mul_69_18_n_1598),
    .Y(u5_mul_69_18_n_1697));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27159 (.A(n_14368),
    .B(u5_mul_69_18_n_1468),
    .C(u5_mul_69_18_n_1597),
    .Y(u5_mul_69_18_n_1696));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27160 (.A(u5_mul_69_18_n_1606),
    .B(u5_mul_69_18_n_1496),
    .Y(u5_mul_69_18_n_1695));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27161 (.A(u5_mul_69_18_n_1548),
    .B(u5_mul_69_18_n_1565),
    .C(n_14351),
    .Y(u5_mul_69_18_n_1694));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27162 (.A(u5_mul_69_18_n_1564),
    .B(u5_mul_69_18_n_1461),
    .C(u5_mul_69_18_n_1583),
    .Y(u5_mul_69_18_n_1692));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27163 (.A(u5_mul_69_18_n_1602),
    .B(u5_mul_69_18_n_1520),
    .Y(u5_mul_69_18_n_1691));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27165 (.A(u5_mul_69_18_n_1628),
    .B(u5_mul_69_18_n_1523),
    .Y(u5_mul_69_18_n_1689));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27166 (.A(n_14373),
    .B(n_14414),
    .C(u5_mul_69_18_n_1477),
    .Y(u5_mul_69_18_n_1688));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27168 (.A(u5_mul_69_18_n_1570),
    .B(n_14348),
    .Y(u5_mul_69_18_n_1687));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27169 (.A1(n_14362),
    .A2(u5_mul_69_18_n_1569),
    .B(u5_mul_69_18_n_1643),
    .Y(u5_mul_69_18_n_1680));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27170 (.A(u5_mul_69_18_n_1572),
    .B(u5_mul_69_18_n_1622),
    .Y(u5_mul_69_18_n_1686));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27171 (.A(u5_mul_69_18_n_1572),
    .B(u5_mul_69_18_n_1622),
    .Y(u5_mul_69_18_n_1679));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27172 (.A1(u5_mul_69_18_n_1501),
    .A2(u5_mul_69_18_n_1600),
    .B(u5_mul_69_18_n_1642),
    .Y(u5_mul_69_18_n_1678));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27173 (.A(n_14359),
    .B(u5_mul_69_18_n_1518),
    .Y(u5_mul_69_18_n_1677));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27178 (.A(u5_mul_69_18_n_1570),
    .B(n_14348),
    .Y(u5_mul_69_18_n_1673));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27182 (.A(u5_mul_69_18_n_1561),
    .B(n_14355),
    .Y(u5_mul_69_18_n_1669));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27183 (.A(n_14356),
    .B(u5_mul_69_18_n_1469),
    .Y(u5_mul_69_18_n_1668));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27186 (.A(u5_mul_69_18_n_1575),
    .B(u5_mul_69_18_n_1532),
    .Y(u5_mul_69_18_n_1684));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27188 (.A(u5_mul_69_18_n_1574),
    .B(n_14389),
    .Y(u5_mul_69_18_n_1682));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27190 (.A(u5_mul_69_18_n_1534),
    .B(u5_mul_69_18_n_1305),
    .C(n_14377),
    .Y(u5_mul_69_18_n_1665));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27192 (.A(n_14381),
    .B(n_14415),
    .C(u5_mul_69_18_n_1362),
    .Y(u5_mul_69_18_n_1664));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27194 (.A(n_14357),
    .B(u5_mul_69_18_n_1413),
    .Y(u5_mul_69_18_n_1649));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27196 (.A(n_14380),
    .B(u5_mul_69_18_n_1316),
    .C(u5_mul_69_18_n_1499),
    .Y(u5_mul_69_18_n_1663));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27197 (.A(n_14368),
    .B(u5_mul_69_18_n_1468),
    .Y(u5_mul_69_18_n_1647));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27201 (.A(u5_mul_69_18_n_1524),
    .B(u5_mul_69_18_n_1488),
    .C(u5_mul_69_18_n_1464),
    .Y(u5_mul_69_18_n_1662));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27202 (.A(u5_mul_69_18_n_1532),
    .B(n_14404),
    .C(u5_mul_69_18_n_1425),
    .Y(u5_mul_69_18_n_1661));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27203 (.A(u5_mul_69_18_n_1475),
    .B(u5_mul_69_18_n_1365),
    .C(n_14385),
    .Y(u5_mul_69_18_n_1660));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27204 (.A(n_14387),
    .B(u5_mul_69_18_n_1234),
    .C(u5_mul_69_18_n_1496),
    .Y(u5_mul_69_18_n_1659));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27205 (.A(u5_mul_69_18_n_1466),
    .B(n_14383),
    .C(u5_mul_69_18_n_1476),
    .Y(u5_mul_69_18_n_1658));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27206 (.A(u5_mul_69_18_n_1465),
    .B(u5_mul_69_18_n_1423),
    .C(u5_mul_69_18_n_1531),
    .Y(u5_mul_69_18_n_1657));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27207 (.A(u5_mul_69_18_n_1528),
    .B(n_14390),
    .C(u5_mul_69_18_n_1484),
    .Y(u5_mul_69_18_n_1656));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27208 (.A(u5_mul_69_18_n_1541),
    .B(u5_mul_69_18_n_1479),
    .Y(u5_mul_69_18_n_1655));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27209 (.A(u5_mul_69_18_n_1520),
    .B(n_14382),
    .C(u5_mul_69_18_n_1478),
    .Y(u5_mul_69_18_n_1654));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27210 (.A(u5_mul_69_18_n_1523),
    .B(u5_mul_69_18_n_1323),
    .C(u5_mul_69_18_n_1495),
    .Y(u5_mul_69_18_n_1653));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27211 (.A(u5_mul_69_18_n_1471),
    .B(u5_mul_69_18_n_1422),
    .C(u5_mul_69_18_n_1514),
    .Y(u5_mul_69_18_n_1652));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27213 (.A(n_14362),
    .B(u5_mul_69_18_n_1569),
    .Y(u5_mul_69_18_n_1643));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27214 (.A1(u5_mul_69_18_n_1389),
    .A2(u5_mul_69_18_n_1540),
    .B(u5_mul_69_18_n_1599),
    .Y(u5_mul_69_18_n_1634));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27215 (.A1(u5_mul_69_18_n_1426),
    .A2(n_14375),
    .B(u5_mul_69_18_n_1601),
    .Y(u5_mul_69_18_n_1633));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27216 (.A(u5_mul_69_18_n_1600),
    .B(u5_mul_69_18_n_1501),
    .Y(u5_mul_69_18_n_1642));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27217 (.A(u5_mul_69_18_n_1501),
    .B(u5_mul_69_18_n_1600),
    .Y(u5_mul_69_18_n_1632));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27221 (.A(u5_mul_69_18_n_1495),
    .B(u5_mul_69_18_n_1323),
    .Y(u5_mul_69_18_n_1628));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27222 (.A(u5_mul_69_18_n_1489),
    .B(n_14394),
    .Y(u5_mul_69_18_n_1627));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27223 (.A(n_14362),
    .B(u5_mul_69_18_n_1569),
    .Y(u5_mul_69_18_n_1626));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27224 (.A(u5_mul_69_18_n_1514),
    .B(u5_mul_69_18_n_1422),
    .Y(u5_mul_69_18_n_1625));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27225 (.A(n_14386),
    .B(u5_mul_69_18_n_1517),
    .Y(u5_mul_69_18_n_1624));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27226 (.A1(u5_mul_69_18_n_1391),
    .A2(u5_mul_69_18_n_1535),
    .B(u5_mul_69_18_n_1379),
    .Y(u5_mul_69_18_n_1641));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27228 (.A(u5_mul_69_18_n_1510),
    .B(n_14405),
    .Y(u5_mul_69_18_n_1639));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27229 (.A(n_14376),
    .B(u5_mul_69_18_n_1449),
    .Y(u5_mul_69_18_n_1638));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27240 (.A(n_14387),
    .B(u5_mul_69_18_n_1234),
    .Y(u5_mul_69_18_n_1606));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27242 (.A(u5_mul_69_18_n_1418),
    .B(u5_mul_69_18_n_1197),
    .C(u5_mul_69_18_n_1455),
    .Y(u5_mul_69_18_n_1622));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27243 (.A(u5_mul_69_18_n_1527),
    .B(u5_mul_69_18_n_1500),
    .Y(u5_mul_69_18_n_1604));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27245 (.A(u5_mul_69_18_n_1478),
    .B(n_14382),
    .Y(u5_mul_69_18_n_1602));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27246 (.A(u5_mul_69_18_n_1498),
    .B(u5_mul_69_18_n_1384),
    .C(u5_mul_69_18_n_1411),
    .Y(u5_mul_69_18_n_1621));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27247 (.A(u5_mul_69_18_n_1481),
    .B(u5_mul_69_18_n_1188),
    .C(n_14402),
    .Y(u5_mul_69_18_n_1620));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27248 (.A(n_14376),
    .B(u5_mul_69_18_n_1195),
    .C(u5_mul_69_18_n_1322),
    .Y(u5_mul_69_18_n_1619));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27249 (.A(u5_mul_69_18_n_1537),
    .B(n_14408),
    .C(u5_mul_69_18_n_1354),
    .Y(u5_mul_69_18_n_1618));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27250 (.A(u5_mul_69_18_n_1479),
    .B(u5_mul_69_18_n_1386),
    .C(u5_mul_69_18_n_1412),
    .Y(u5_mul_69_18_n_1617));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27251 (.A(u5_mul_69_18_n_1483),
    .B(n_14442),
    .C(u5_mul_69_18_n_1357),
    .Y(u5_mul_69_18_n_1616));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27253 (.A(u5_mul_69_18_n_1487),
    .B(u5_mul_69_18_n_1326),
    .C(u5_mul_69_18_n_1361),
    .Y(u5_mul_69_18_n_1614));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27255 (.A(u5_mul_69_18_n_1424),
    .B(n_14417),
    .C(n_14389),
    .Y(u5_mul_69_18_n_1612));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27257 (.A1(u5_mul_69_18_n_1367),
    .A2(n_14388),
    .B(u5_mul_69_18_n_1538),
    .Y(u5_mul_69_18_n_1579));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27258 (.A(u5_mul_69_18_n_1426),
    .B(n_14375),
    .Y(u5_mul_69_18_n_1601));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27259 (.A(u5_mul_69_18_n_1426),
    .B(n_14375),
    .Y(u5_mul_69_18_n_1578));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27260 (.A(u5_mul_69_18_n_1457),
    .B(u5_mul_69_18_n_1447),
    .Y(u5_mul_69_18_n_1600));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27261 (.A(u5_mul_69_18_n_1389),
    .B(u5_mul_69_18_n_1540),
    .Y(u5_mul_69_18_n_1577));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27263 (.A(u5_mul_69_18_n_1389),
    .B(u5_mul_69_18_n_1540),
    .Y(u5_mul_69_18_n_1599));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27264 (.A(u5_mul_69_18_n_1425),
    .B(n_14404),
    .Y(u5_mul_69_18_n_1575));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27265 (.A(u5_mul_69_18_n_1424),
    .B(n_14417),
    .Y(u5_mul_69_18_n_1574));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27267 (.A(u5_mul_69_18_n_1405),
    .B(u5_mul_69_18_n_1279),
    .Y(u5_mul_69_18_n_1598));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27268 (.A(u5_mul_69_18_n_1446),
    .B(u5_mul_69_18_n_1319),
    .Y(u5_mul_69_18_n_1597));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27271 (.A(u5_mul_69_18_n_1444),
    .B(u5_mul_69_18_n_1382),
    .Y(u5_mul_69_18_n_1594));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27274 (.A(u5_mul_69_18_n_1429),
    .B(u5_mul_69_18_n_1330),
    .Y(u5_mul_69_18_n_1591));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27278 (.A(u5_mul_69_18_n_1437),
    .B(n_14396),
    .Y(u5_mul_69_18_n_1587));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27283 (.A(u5_mul_69_18_n_1445),
    .B(u5_mul_69_18_n_705),
    .Y(u5_mul_69_18_n_1583));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27285 (.A(u5_mul_69_18_n_1407),
    .B(u5_mul_69_18_n_1313),
    .Y(u5_mul_69_18_n_1581));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27286 (.A(u5_mul_69_18_n_1551),
    .Y(u5_mul_69_18_n_1552));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27287 (.A(u5_mul_69_18_n_1549),
    .Y(u5_mul_69_18_n_1550));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27288 (.A(u5_mul_69_18_n_1416),
    .B(u5_mul_69_18_n_1427),
    .Y(u5_mul_69_18_n_1572));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27289 (.A(u5_mul_69_18_n_1412),
    .B(u5_mul_69_18_n_1386),
    .Y(u5_mul_69_18_n_1541));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27291 (.A(u5_mul_69_18_n_1458),
    .B(u5_mul_69_18_n_1199),
    .C(u5_mul_69_18_n_1301),
    .Y(u5_mul_69_18_n_1570));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27292 (.A(u5_mul_69_18_n_1416),
    .B(u5_mul_69_18_n_1190),
    .C(n_14423),
    .Y(u5_mul_69_18_n_1569));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27293 (.A(u5_mul_69_18_n_1417),
    .B(n_14451),
    .C(u5_mul_69_18_n_1358),
    .Y(u5_mul_69_18_n_1568));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27294 (.A(u5_mul_69_18_n_1415),
    .B(n_14407),
    .C(u5_mul_69_18_n_1239),
    .Y(u5_mul_69_18_n_1567));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27295 (.A(u5_mul_69_18_n_1421),
    .B(u5_mul_69_18_n_1200),
    .C(n_14393),
    .Y(u5_mul_69_18_n_1566));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27296 (.A(u5_mul_69_18_n_1420),
    .B(u5_mul_69_18_n_1196),
    .C(u5_mul_69_18_n_1236),
    .Y(u5_mul_69_18_n_1565));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27297 (.A(u5_mul_69_18_n_1419),
    .B(n_14410),
    .C(n_14395),
    .Y(u5_mul_69_18_n_1564));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27298 (.A(u5_mul_69_18_n_1356),
    .B(u5_mul_69_18_n_1218),
    .C(n_14403),
    .Y(u5_mul_69_18_n_1563));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27300 (.A(u5_mul_69_18_n_1383),
    .B(u5_mul_69_18_n_1226),
    .C(u5_mul_69_18_n_1268),
    .Y(u5_mul_69_18_n_1561));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27301 (.A(u5_mul_69_18_n_1402),
    .B(u5_mul_69_18_n_1149),
    .Y(u5_mul_69_18_n_1560));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27303 (.A(u5_mul_69_18_n_1441),
    .B(n_14441),
    .Y(u5_mul_69_18_n_1558));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27307 (.A(u5_mul_69_18_n_1410),
    .B(n_14426),
    .Y(u5_mul_69_18_n_1554));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27309 (.A(u5_mul_69_18_n_1404),
    .B(u5_mul_69_18_n_1265),
    .Y(u5_mul_69_18_n_1551));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27310 (.A(u5_mul_69_18_n_1409),
    .B(u5_mul_69_18_n_1277),
    .Y(u5_mul_69_18_n_1549));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27311 (.A(u5_mul_69_18_n_1395),
    .B(u5_mul_69_18_n_1140),
    .Y(u5_mul_69_18_n_1548));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27313 (.A(u5_mul_69_18_n_1448),
    .B(u5_mul_69_18_n_1134),
    .Y(u5_mul_69_18_n_1546));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27320 (.A1(n_14391),
    .A2(u5_mul_69_18_n_1284),
    .B(u5_mul_69_18_n_1460),
    .Y(u5_mul_69_18_n_1511));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27321 (.A(u5_mul_69_18_n_1366),
    .B(u5_mul_69_18_n_1186),
    .Y(u5_mul_69_18_n_1510));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27324 (.A(u5_mul_69_18_n_1303),
    .B(u5_mul_69_18_n_845),
    .C(u5_mul_69_18_n_1210),
    .Y(u5_mul_69_18_n_1540));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27330 (.A(u5_mul_69_18_n_1367),
    .B(n_14388),
    .Y(u5_mul_69_18_n_1503));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27332 (.A(u5_mul_69_18_n_1367),
    .B(n_14388),
    .Y(u5_mul_69_18_n_1538));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27333 (.A(u5_mul_69_18_n_1311),
    .B(u5_mul_69_18_n_1225),
    .C(u5_mul_69_18_n_1267),
    .Y(u5_mul_69_18_n_1537));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27335 (.A1(u5_mul_69_18_n_1393),
    .A2(u5_mul_69_18_n_1335),
    .B(u5_mul_69_18_n_14),
    .Y(u5_mul_69_18_n_1535));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27336 (.A(n_14455),
    .B(u5_mul_69_18_n_1000),
    .C(u5_mul_69_18_n_1215),
    .Y(u5_mul_69_18_n_1534));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27338 (.A(u5_mul_69_18_n_1372),
    .B(n_14440),
    .Y(u5_mul_69_18_n_1532));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27339 (.A(u5_mul_69_18_n_1375),
    .B(u5_mul_69_18_n_1165),
    .Y(u5_mul_69_18_n_1531));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27342 (.A(u5_mul_69_18_n_1378),
    .B(n_14418),
    .Y(u5_mul_69_18_n_1528));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27343 (.A(u5_mul_69_18_n_1368),
    .B(u5_mul_69_18_n_1194),
    .Y(u5_mul_69_18_n_1527));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27346 (.A(u5_mul_69_18_n_1346),
    .B(u5_mul_69_18_n_1142),
    .Y(u5_mul_69_18_n_1524));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27347 (.A(u5_mul_69_18_n_1353),
    .B(u5_mul_69_18_n_1124),
    .Y(u5_mul_69_18_n_1523));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27350 (.A(u5_mul_69_18_n_1343),
    .B(u5_mul_69_18_n_1249),
    .Y(u5_mul_69_18_n_1520));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27352 (.A(u5_mul_69_18_n_1344),
    .B(n_14458),
    .Y(u5_mul_69_18_n_1518));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27353 (.A(n_14450),
    .B(u5_mul_69_18_n_1224),
    .C(u5_mul_69_18_n_1327),
    .Y(u5_mul_69_18_n_1517));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27356 (.A(u5_mul_69_18_n_1371),
    .B(u5_mul_69_18_n_1169),
    .Y(u5_mul_69_18_n_1514));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27358 (.A(u5_mul_69_18_n_1492),
    .Y(u5_mul_69_18_n_1493));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27360 (.A(u5_mul_69_18_n_1329),
    .B(u5_mul_69_18_n_1158),
    .C(n_14460),
    .Y(u5_mul_69_18_n_1501));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27361 (.A(u5_mul_69_18_n_1277),
    .B(n_14422),
    .C(n_14430),
    .Y(u5_mul_69_18_n_1500));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27362 (.A(u5_mul_69_18_n_1312),
    .B(u5_mul_69_18_n_1221),
    .C(n_14421),
    .Y(u5_mul_69_18_n_1499));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27363 (.A(u5_mul_69_18_n_1246),
    .B(u5_mul_69_18_n_1219),
    .C(u5_mul_69_18_n_1332),
    .Y(u5_mul_69_18_n_1498));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27364 (.A(n_14425),
    .B(u5_mul_69_18_n_1202),
    .C(u5_mul_69_18_n_1291),
    .Y(u5_mul_69_18_n_1497));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27365 (.A(n_14448),
    .B(u5_mul_69_18_n_1171),
    .C(n_14449),
    .Y(u5_mul_69_18_n_1496));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27366 (.A(n_14447),
    .B(u5_mul_69_18_n_1130),
    .C(u5_mul_69_18_n_1278),
    .Y(u5_mul_69_18_n_1495));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27367 (.A(n_14431),
    .B(u5_mul_69_18_n_1217),
    .C(u5_mul_69_18_n_1189),
    .Y(u5_mul_69_18_n_1494));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27368 (.A(u5_mul_69_18_n_1324),
    .B(u5_mul_69_18_n_1339),
    .C(n_14446),
    .Y(u5_mul_69_18_n_1492));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27369 (.A(n_14392),
    .B(n_14420),
    .C(u5_mul_69_18_n_1232),
    .Y(u5_mul_69_18_n_1491));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27370 (.A(u5_mul_69_18_n_1266),
    .B(u5_mul_69_18_n_207),
    .C(u5_mul_69_18_n_1206),
    .Y(u5_mul_69_18_n_1490));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27371 (.A(n_14416),
    .B(u5_mul_69_18_n_1216),
    .C(u5_mul_69_18_n_1133),
    .Y(u5_mul_69_18_n_1489));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27372 (.A(n_14418),
    .B(u5_mul_69_18_n_1208),
    .C(u5_mul_69_18_n_1135),
    .Y(u5_mul_69_18_n_1488));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27373 (.A(n_14443),
    .B(u5_mul_69_18_n_1157),
    .C(u5_mul_69_18_n_1140),
    .Y(u5_mul_69_18_n_1487));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27374 (.A(u5_mul_69_18_n_1330),
    .B(u5_mul_69_18_n_1172),
    .C(n_14412),
    .Y(u5_mul_69_18_n_1486));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27375 (.A(u5_mul_69_18_n_1295),
    .B(u5_mul_69_18_n_1152),
    .C(n_14441),
    .Y(u5_mul_69_18_n_1485));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27376 (.A(n_14428),
    .B(u5_mul_69_18_n_1149),
    .C(n_14419),
    .Y(u5_mul_69_18_n_1484));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27377 (.A(n_14444),
    .B(u5_mul_69_18_n_1211),
    .C(n_14429),
    .Y(u5_mul_69_18_n_1483));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27378 (.A(u5_mul_69_18_n_1298),
    .B(u5_mul_69_18_n_1147),
    .C(n_14437),
    .Y(u5_mul_69_18_n_1482));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27379 (.A(n_14439),
    .B(u5_mul_69_18_n_1148),
    .C(n_14411),
    .Y(u5_mul_69_18_n_1481));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27380 (.A(u5_mul_69_18_n_1364),
    .B(n_14452),
    .C(n_14453),
    .Y(u5_mul_69_18_n_1480));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27381 (.A(u5_mul_69_18_n_1241),
    .B(u5_mul_69_18_n_1128),
    .C(n_14399),
    .Y(u5_mul_69_18_n_1479));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27382 (.A(n_14436),
    .B(u5_mul_69_18_n_1222),
    .C(u5_mul_69_18_n_1144),
    .Y(u5_mul_69_18_n_1478));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27383 (.A(u5_mul_69_18_n_1256),
    .B(u5_mul_69_18_n_1173),
    .C(u5_mul_69_18_n_1134),
    .Y(u5_mul_69_18_n_1477));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27384 (.A(n_14445),
    .B(u5_mul_69_18_n_1164),
    .C(u5_mul_69_18_n_1306),
    .Y(u5_mul_69_18_n_1476));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27385 (.A(u5_mul_69_18_n_1257),
    .B(u5_mul_69_18_n_1203),
    .C(u5_mul_69_18_n_1137),
    .Y(u5_mul_69_18_n_1475));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27386 (.A(n_14435),
    .B(u5_mul_69_18_n_1153),
    .C(u5_mul_69_18_n_1265),
    .Y(u5_mul_69_18_n_1474));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27387 (.A(n_14433),
    .B(u5_mul_69_18_n_1161),
    .C(u5_mul_69_18_n_1125),
    .Y(u5_mul_69_18_n_1473));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27388 (.A(u5_mul_69_18_n_1363),
    .B(n_14456),
    .C(u5_mul_69_18_n_1260),
    .Y(u5_mul_69_18_n_1472));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27389 (.A(n_14409),
    .B(u5_mul_69_18_n_704),
    .C(u5_mul_69_18_n_1160),
    .Y(u5_mul_69_18_n_1471));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27390 (.A(u5_mul_69_18_n_1249),
    .B(u5_mul_69_18_n_1150),
    .C(u5_mul_69_18_n_1139),
    .Y(u5_mul_69_18_n_1470));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27391 (.A(n_14440),
    .B(u5_mul_69_18_n_1209),
    .C(u5_mul_69_18_n_1143),
    .Y(u5_mul_69_18_n_1469));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27392 (.A(u5_mul_69_18_n_1313),
    .B(n_14424),
    .C(n_14438),
    .Y(u5_mul_69_18_n_1468));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27393 (.A(n_14413),
    .B(u5_mul_69_18_n_695),
    .C(u5_mul_69_18_n_1229),
    .Y(u5_mul_69_18_n_1467));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27394 (.A(u5_mul_69_18_n_1366),
    .B(u5_mul_69_18_n_1187),
    .C(n_14405),
    .Y(u5_mul_69_18_n_1466));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27395 (.A(u5_mul_69_18_n_1247),
    .B(n_14459),
    .C(n_14426),
    .Y(u5_mul_69_18_n_1465));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27396 (.A(n_14432),
    .B(u5_mul_69_18_n_1258),
    .C(u5_mul_69_18_n_1205),
    .Y(u5_mul_69_18_n_1464));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27397 (.A(u5_mul_69_18_n_1320),
    .B(u5_mul_69_18_n_1212),
    .C(n_14454),
    .Y(u5_mul_69_18_n_1463));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27398 (.A(n_14406),
    .B(u5_mul_69_18_n_1131),
    .C(u5_mul_69_18_n_1213),
    .Y(u5_mul_69_18_n_1462));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27399 (.A(u5_mul_69_18_n_1270),
    .B(n_14434),
    .C(u5_mul_69_18_n_1279),
    .Y(u5_mul_69_18_n_1461));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27400 (.A(u5_mul_69_18_n_1457),
    .Y(u5_mul_69_18_n_1458));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27402 (.A1(n_14398),
    .A2(u5_mul_69_18_n_1063),
    .B(u5_mul_69_18_n_1391),
    .Y(u5_mul_69_18_n_1453));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27403 (.A(u5_mul_69_18_n_1284),
    .B(n_14391),
    .Y(u5_mul_69_18_n_1452));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27404 (.A(u5_mul_69_18_n_1284),
    .B(n_14391),
    .Y(u5_mul_69_18_n_1460));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27407 (.A(u5_mul_69_18_n_1322),
    .B(u5_mul_69_18_n_1195),
    .Y(u5_mul_69_18_n_1449));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27408 (.A(u5_mul_69_18_n_1256),
    .B(u5_mul_69_18_n_1173),
    .Y(u5_mul_69_18_n_1448));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27409 (.A(u5_mul_69_18_n_1301),
    .B(u5_mul_69_18_n_1199),
    .Y(u5_mul_69_18_n_1447));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27410 (.A(n_14454),
    .B(u5_mul_69_18_n_1212),
    .Y(u5_mul_69_18_n_1446));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27411 (.A(n_14409),
    .B(u5_mul_69_18_n_1160),
    .Y(u5_mul_69_18_n_1445));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27412 (.A(u5_mul_69_18_n_1268),
    .B(u5_mul_69_18_n_1226),
    .Y(u5_mul_69_18_n_1444));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27415 (.A(u5_mul_69_18_n_1295),
    .B(u5_mul_69_18_n_1152),
    .Y(u5_mul_69_18_n_1441));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27417 (.A(u5_mul_69_18_n_1392),
    .B(u5_mul_69_18_n_14),
    .Y(u5_mul_69_18_n_1439));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27419 (.A(n_14403),
    .B(u5_mul_69_18_n_1218),
    .Y(u5_mul_69_18_n_1437));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27428 (.A(n_14412),
    .B(u5_mul_69_18_n_1172),
    .Y(u5_mul_69_18_n_1429));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27430 (.A(n_14423),
    .B(u5_mul_69_18_n_1190),
    .Y(u5_mul_69_18_n_1427));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27431 (.A(u5_mul_69_18_n_1285),
    .B(u5_mul_69_18_n_1061),
    .Y(u5_mul_69_18_n_1457));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27433 (.A(n_14401),
    .B(u5_mul_69_18_n_1097),
    .Y(u5_mul_69_18_n_1455));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27435 (.A(u5_mul_69_18_n_1247),
    .B(n_14459),
    .Y(u5_mul_69_18_n_1410));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27436 (.A(n_14430),
    .B(n_14422),
    .Y(u5_mul_69_18_n_1409));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27438 (.A(n_14438),
    .B(n_14424),
    .Y(u5_mul_69_18_n_1407));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27440 (.A(u5_mul_69_18_n_1270),
    .B(n_14434),
    .Y(u5_mul_69_18_n_1405));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27441 (.A(n_14435),
    .B(u5_mul_69_18_n_1153),
    .Y(u5_mul_69_18_n_1404));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27442 (.A(n_14427),
    .B(u5_mul_69_18_n_992),
    .C(u5_mul_69_18_n_1060),
    .Y(u5_mul_69_18_n_1426));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27444 (.A(n_14428),
    .B(n_14419),
    .Y(u5_mul_69_18_n_1402));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27451 (.A(n_14443),
    .B(u5_mul_69_18_n_1157),
    .Y(u5_mul_69_18_n_1395));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27453 (.A(u5_mul_69_18_n_1163),
    .B(u5_mul_69_18_n_1198),
    .C(u5_mul_69_18_n_1116),
    .Y(u5_mul_69_18_n_1425));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27454 (.A(u5_mul_69_18_n_1142),
    .B(u5_mul_69_18_n_999),
    .C(u5_mul_69_18_n_1207),
    .Y(u5_mul_69_18_n_1424));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27455 (.A(u5_mul_69_18_n_1145),
    .B(u5_mul_69_18_n_872),
    .C(u5_mul_69_18_n_1168),
    .Y(u5_mul_69_18_n_1423));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27456 (.A(u5_mul_69_18_n_1191),
    .B(u5_mul_69_18_n_1159),
    .C(u5_mul_69_18_n_1201),
    .Y(u5_mul_69_18_n_1422));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27457 (.A(u5_mul_69_18_n_1129),
    .B(n_14458),
    .C(u5_mul_69_18_n_1151),
    .Y(u5_mul_69_18_n_1421));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27458 (.A(u5_mul_69_18_n_1169),
    .B(u5_mul_69_18_n_704),
    .C(u5_mul_69_18_n_1193),
    .Y(u5_mul_69_18_n_1420));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27459 (.A(u5_mul_69_18_n_1132),
    .B(u5_mul_69_18_n_1204),
    .C(u5_mul_69_18_n_1138),
    .Y(u5_mul_69_18_n_1419));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27460 (.A(u5_mul_69_18_n_1123),
    .B(u5_mul_69_18_n_699),
    .C(u5_mul_69_18_n_1214),
    .Y(u5_mul_69_18_n_1418));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27461 (.A(n_14400),
    .B(u5_mul_69_18_n_703),
    .C(u5_mul_69_18_n_1127),
    .Y(u5_mul_69_18_n_1417));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27462 (.A(n_14401),
    .B(u5_mul_69_18_n_887),
    .C(u5_mul_69_18_n_699),
    .Y(u5_mul_69_18_n_1416));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27463 (.A(u5_mul_69_18_n_1162),
    .B(u5_mul_69_18_n_991),
    .C(u5_mul_69_18_n_1194),
    .Y(u5_mul_69_18_n_1415));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27465 (.A(u5_mul_69_18_n_1165),
    .B(u5_mul_69_18_n_1059),
    .C(u5_mul_69_18_n_1136),
    .Y(u5_mul_69_18_n_1413));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27466 (.A(u5_mul_69_18_n_1124),
    .B(u5_mul_69_18_n_698),
    .C(u5_mul_69_18_n_1166),
    .Y(u5_mul_69_18_n_1412));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27467 (.A(u5_mul_69_18_n_1141),
    .B(u5_mul_69_18_n_173),
    .C(u5_mul_69_18_n_1175),
    .Y(u5_mul_69_18_n_1411));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27468 (.A(u5_mul_69_18_n_1392),
    .Y(u5_mul_69_18_n_1393));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27469 (.A(u5_mul_69_18_n_1382),
    .Y(u5_mul_69_18_n_1383));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27471 (.A(u5_mul_69_18_n_984),
    .B(n_14397),
    .Y(u5_mul_69_18_n_1392));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27472 (.A(u5_mul_69_18_n_1063),
    .B(n_14398),
    .Y(u5_mul_69_18_n_1391));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27473 (.A(u5_mul_69_18_n_1063),
    .B(n_14398),
    .Y(u5_mul_69_18_n_1379));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27474 (.A(u5_mul_69_18_n_1135),
    .B(u5_mul_69_18_n_1208),
    .Y(u5_mul_69_18_n_1378));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27478 (.A(u5_mul_69_18_n_1136),
    .B(u5_mul_69_18_n_1059),
    .Y(u5_mul_69_18_n_1375));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27481 (.A(u5_mul_69_18_n_1209),
    .B(u5_mul_69_18_n_1143),
    .Y(u5_mul_69_18_n_1372));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27483 (.A1(u5_mul_69_18_n_704),
    .A2(u5_mul_69_18_n_1192),
    .B1(u5_mul_69_18_n_705),
    .B2(u5_mul_69_18_n_1193),
    .Y(u5_mul_69_18_n_1371));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27486 (.A(u5_mul_69_18_n_1223),
    .B(u5_mul_69_18_n_1078),
    .Y(u5_mul_69_18_n_1389));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27487 (.A(u5_mul_69_18_n_1162),
    .B(u5_mul_69_18_n_991),
    .Y(u5_mul_69_18_n_1368));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27490 (.A(u5_mul_69_18_n_1227),
    .B(u5_mul_69_18_n_1085),
    .Y(u5_mul_69_18_n_1386));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27492 (.A(u5_mul_69_18_n_1174),
    .B(u5_mul_69_18_n_1103),
    .Y(u5_mul_69_18_n_1384));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27493 (.A(u5_mul_69_18_n_1156),
    .B(u5_mul_69_18_n_1109),
    .Y(u5_mul_69_18_n_1382));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27495 (.A(n_14396),
    .Y(u5_mul_69_18_n_1356));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27496 (.A(u5_mul_69_18_n_1166),
    .B(u5_mul_69_18_n_698),
    .Y(u5_mul_69_18_n_1353));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27497 (.A(u5_mul_69_18_n_1223),
    .B(u5_mul_69_18_n_166),
    .C(u5_mul_69_18_n_884),
    .Y(u5_mul_69_18_n_1352));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27499 (.A(n_14457),
    .B(u5_mul_69_18_n_905),
    .C(u5_mul_69_18_n_855),
    .Y(u5_mul_69_18_n_1367));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27504 (.A(u5_mul_69_18_n_1207),
    .B(u5_mul_69_18_n_999),
    .Y(u5_mul_69_18_n_1346));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27506 (.A(u5_mul_69_18_n_1129),
    .B(u5_mul_69_18_n_1151),
    .Y(u5_mul_69_18_n_1344));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27507 (.A(u5_mul_69_18_n_1139),
    .B(u5_mul_69_18_n_1150),
    .Y(u5_mul_69_18_n_1343));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27509 (.A(u5_mul_69_18_n_1170),
    .B(u5_mul_69_18_n_174),
    .C(u5_mul_69_18_n_696),
    .Y(u5_mul_69_18_n_1366));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27510 (.A(u5_mul_69_18_n_1154),
    .B(u5_mul_69_18_n_874),
    .C(u5_mul_69_18_n_1001),
    .Y(u5_mul_69_18_n_1365));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27511 (.A(u5_mul_69_18_n_1220),
    .B(u5_mul_69_18_n_784),
    .C(u5_mul_69_18_n_1002),
    .Y(u5_mul_69_18_n_1364));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27512 (.A(u5_mul_69_18_n_1146),
    .B(u5_mul_69_18_n_851),
    .C(u5_mul_69_18_n_1117),
    .Y(u5_mul_69_18_n_1363));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27513 (.A(u5_mul_69_18_n_1118),
    .B(u5_mul_69_18_n_890),
    .C(u5_mul_69_18_n_1061),
    .Y(u5_mul_69_18_n_1362));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27514 (.A(u5_mul_69_18_n_1228),
    .B(u5_mul_69_18_n_214),
    .C(u5_mul_69_18_n_907),
    .Y(u5_mul_69_18_n_1361));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27515 (.A(u5_mul_69_18_n_1156),
    .B(u5_mul_69_18_n_184),
    .C(u5_mul_69_18_n_847),
    .Y(u5_mul_69_18_n_1360));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27516 (.A(u5_mul_69_18_n_1176),
    .B(u5_mul_69_18_n_210),
    .C(u5_mul_69_18_n_706),
    .Y(u5_mul_69_18_n_1359));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27517 (.A(u5_mul_69_18_n_1170),
    .B(u5_mul_69_18_n_1084),
    .Y(u5_mul_69_18_n_1358));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27518 (.A(u5_mul_69_18_n_1155),
    .B(u5_mul_69_18_n_773),
    .C(u5_mul_69_18_n_998),
    .Y(u5_mul_69_18_n_1357));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27520 (.A(u5_mul_69_18_n_1174),
    .B(u5_mul_69_18_n_169),
    .C(u5_mul_69_18_n_863),
    .Y(u5_mul_69_18_n_1354));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27522 (.A(u5_mul_69_18_n_1331),
    .Y(u5_mul_69_18_n_1332));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27523 (.A(u5_mul_69_18_n_1319),
    .Y(u5_mul_69_18_n_1320));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27524 (.A(u5_mul_69_18_n_1310),
    .Y(u5_mul_69_18_n_1311));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27531 (.A(u5_mul_69_18_n_1118),
    .B(u5_mul_69_18_n_890),
    .Y(u5_mul_69_18_n_1285));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27532 (.A(u5_mul_69_18_n_1014),
    .B(u5_mul_69_18_n_667),
    .Y(u5_mul_69_18_n_1339));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27536 (.A1(u5_mul_69_18_n_1121),
    .A2(u5_mul_69_18_n_1114),
    .B(u5_mul_69_18_n_1122),
    .Y(u5_mul_69_18_n_1335));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27539 (.A(u5_mul_69_18_n_1057),
    .B(u5_mul_69_18_n_976),
    .Y(u5_mul_69_18_n_1331));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27540 (.A(u5_mul_69_18_n_1023),
    .B(u5_mul_69_18_n_974),
    .Y(u5_mul_69_18_n_1330));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27541 (.A(u5_mul_69_18_n_1050),
    .B(u5_mul_69_18_n_956),
    .Y(u5_mul_69_18_n_1329));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27543 (.A(u5_mul_69_18_n_1094),
    .B(u5_mul_69_18_n_703),
    .Y(u5_mul_69_18_n_1327));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27544 (.A(u5_mul_69_18_n_1093),
    .B(u5_mul_69_18_n_700),
    .Y(u5_mul_69_18_n_1326));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27546 (.A(u5_mul_69_18_n_1120),
    .B(u5_mul_69_18_n_1012),
    .Y(u5_mul_69_18_n_1324));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27547 (.A(u5_mul_69_18_n_1088),
    .B(u5_mul_69_18_n_972),
    .Y(u5_mul_69_18_n_1323));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27548 (.A(u5_mul_69_18_n_1115),
    .B(u5_mul_69_18_n_216),
    .Y(u5_mul_69_18_n_1322));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27550 (.A(u5_mul_69_18_n_1089),
    .B(u5_mul_69_18_n_981),
    .Y(u5_mul_69_18_n_1319));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27553 (.A(u5_mul_69_18_n_1079),
    .B(u5_mul_69_18_n_978),
    .Y(u5_mul_69_18_n_1316));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27556 (.A(u5_mul_69_18_n_1096),
    .B(u5_mul_69_18_n_968),
    .Y(u5_mul_69_18_n_1313));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27557 (.A(u5_mul_69_18_n_1071),
    .B(u5_mul_69_18_n_815),
    .Y(u5_mul_69_18_n_1312));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27558 (.A(u5_mul_69_18_n_1067),
    .B(u5_mul_69_18_n_835),
    .Y(u5_mul_69_18_n_1310));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27562 (.A(u5_mul_69_18_n_1065),
    .B(u5_mul_69_18_n_820),
    .Y(u5_mul_69_18_n_1306));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27563 (.A(u5_mul_69_18_n_13),
    .B(u5_mul_69_18_n_1042),
    .Y(u5_mul_69_18_n_1305));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27565 (.A(u5_mul_69_18_n_1080),
    .B(u5_mul_69_18_n_179),
    .Y(u5_mul_69_18_n_1303));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27567 (.A(u5_mul_69_18_n_1051),
    .B(u5_mul_69_18_n_676),
    .Y(u5_mul_69_18_n_1301));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27570 (.A(u5_mul_69_18_n_1032),
    .B(u5_mul_69_18_n_658),
    .Y(u5_mul_69_18_n_1298));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27573 (.A(u5_mul_69_18_n_1020),
    .B(u5_mul_69_18_n_666),
    .Y(u5_mul_69_18_n_1295));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27577 (.A(u5_mul_69_18_n_1095),
    .B(u5_mul_69_18_n_701),
    .Y(u5_mul_69_18_n_1291));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27579 (.A(u5_mul_69_18_n_993),
    .B(u5_mul_69_18_n_961),
    .C(u5_mul_69_18_n_785),
    .Y(u5_mul_69_18_n_1284));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27584 (.A(u5_mul_69_18_n_1119),
    .B(u5_mul_69_18_n_868),
    .C(u5_mul_69_18_n_897),
    .Y(u5_mul_69_18_n_1279));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27585 (.A(u5_mul_69_18_n_1009),
    .B(u5_mul_69_18_n_842),
    .Y(u5_mul_69_18_n_1278));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27586 (.A(u5_mul_69_18_n_13),
    .B(u5_mul_69_18_n_927),
    .C(u5_mul_69_18_n_744),
    .Y(u5_mul_69_18_n_1277));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27593 (.A(u5_mul_69_18_n_1044),
    .B(u5_mul_69_18_n_938),
    .Y(u5_mul_69_18_n_1270));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27595 (.A(u5_mul_69_18_n_1040),
    .B(u5_mul_69_18_n_786),
    .Y(u5_mul_69_18_n_1268));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27596 (.A(u5_mul_69_18_n_1041),
    .B(u5_mul_69_18_n_846),
    .Y(u5_mul_69_18_n_1267));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27597 (.A(u5_mul_69_18_n_1037),
    .B(u5_mul_69_18_n_824),
    .Y(u5_mul_69_18_n_1266));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27598 (.A(u5_mul_69_18_n_1034),
    .B(u5_mul_69_18_n_939),
    .Y(u5_mul_69_18_n_1265));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27603 (.A(u5_mul_69_18_n_1029),
    .B(u5_mul_69_18_n_933),
    .Y(u5_mul_69_18_n_1260));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27605 (.A(u5_mul_69_18_n_1026),
    .B(u5_mul_69_18_n_717),
    .Y(u5_mul_69_18_n_1258));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27606 (.A(u5_mul_69_18_n_1106),
    .B(u5_mul_69_18_n_940),
    .Y(u5_mul_69_18_n_1257));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27607 (.A(u5_mul_69_18_n_1024),
    .B(u5_mul_69_18_n_764),
    .Y(u5_mul_69_18_n_1256));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27614 (.A(u5_mul_69_18_n_1100),
    .B(u5_mul_69_18_n_934),
    .Y(u5_mul_69_18_n_1249));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27616 (.A(u5_mul_69_18_n_1036),
    .B(u5_mul_69_18_n_951),
    .Y(u5_mul_69_18_n_1247));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27617 (.A(u5_mul_69_18_n_1027),
    .B(u5_mul_69_18_n_875),
    .Y(u5_mul_69_18_n_1246));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27622 (.A(u5_mul_69_18_n_1008),
    .B(u5_mul_69_18_n_795),
    .Y(u5_mul_69_18_n_1241));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27624 (.A(u5_mul_69_18_n_1035),
    .B(u5_mul_69_18_n_829),
    .Y(u5_mul_69_18_n_1239));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27627 (.A(u5_mul_69_18_n_1048),
    .B(u5_mul_69_18_n_766),
    .Y(u5_mul_69_18_n_1236));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27629 (.A(u5_mul_69_18_n_1062),
    .B(u5_mul_69_18_n_731),
    .C(u5_mul_69_18_n_994),
    .Y(u5_mul_69_18_n_1234));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27631 (.A(u5_mul_69_18_n_1120),
    .B(u5_mul_69_18_n_745),
    .C(u5_mul_69_18_n_929),
    .Y(u5_mul_69_18_n_1232));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27633 (.A(u5_mul_69_18_n_1227),
    .Y(u5_mul_69_18_n_1228));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27634 (.A(u5_mul_69_18_n_1192),
    .Y(u5_mul_69_18_n_1193));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27635 (.A(u5_mul_69_18_n_1186),
    .Y(u5_mul_69_18_n_1187));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27637 (.A1(u5_mul_69_18_n_985),
    .A2(u5_mul_69_18_n_995),
    .B(u5_mul_69_18_n_1122),
    .Y(u5_mul_69_18_n_1181));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27643 (.A(u5_mul_69_18_n_780),
    .B(u5_mul_69_18_n_963),
    .C(u5_mul_69_18_n_757),
    .Y(u5_mul_69_18_n_1229));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27644 (.A(u5_mul_69_18_n_775),
    .B(u5_mul_69_18_n_707),
    .C(u5_mul_69_18_n_930),
    .Y(u5_mul_69_18_n_1227));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27645 (.A(u5_mul_69_18_n_848),
    .B(u5_mul_69_18_n_967),
    .C(u5_mul_69_18_n_893),
    .Y(u5_mul_69_18_n_1226));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27646 (.A(u5_mul_69_18_n_846),
    .B(u5_mul_69_18_n_976),
    .C(u5_mul_69_18_n_886),
    .Y(u5_mul_69_18_n_1225));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27647 (.A(u5_mul_69_18_n_725),
    .B(u5_mul_69_18_n_974),
    .C(u5_mul_69_18_n_779),
    .Y(u5_mul_69_18_n_1224));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27648 (.A(u5_mul_69_18_n_983),
    .B(u5_mul_69_18_n_178),
    .C(u5_mul_69_18_n_918),
    .Y(u5_mul_69_18_n_1223));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27649 (.A(u5_mul_69_18_n_964),
    .B(u5_mul_69_18_n_710),
    .C(u5_mul_69_18_n_701),
    .Y(u5_mul_69_18_n_1222));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27650 (.A(u5_mul_69_18_n_880),
    .B(u5_mul_69_18_n_980),
    .C(u5_mul_69_18_n_899),
    .Y(u5_mul_69_18_n_1221));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27651 (.A(u5_mul_69_18_n_737),
    .B(u5_mul_69_18_n_665),
    .C(u5_mul_69_18_n_790),
    .Y(u5_mul_69_18_n_1220));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27652 (.A(u5_mul_69_18_n_696),
    .B(u5_mul_69_18_n_188),
    .C(u5_mul_69_18_n_977),
    .Y(u5_mul_69_18_n_1219));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27653 (.A(u5_mul_69_18_n_760),
    .B(u5_mul_69_18_n_215),
    .C(u5_mul_69_18_n_975),
    .Y(u5_mul_69_18_n_1218));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27654 (.A(u5_mul_69_18_n_702),
    .B(u5_mul_69_18_n_176),
    .C(u5_mul_69_18_n_982),
    .Y(u5_mul_69_18_n_1217));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27655 (.A(u5_mul_69_18_n_957),
    .B(u5_mul_69_18_n_661),
    .C(u5_mul_69_18_n_889),
    .Y(u5_mul_69_18_n_1216));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27656 (.A(u5_mul_69_18_n_916),
    .B(u5_mul_69_18_n_676),
    .C(u5_mul_69_18_n_962),
    .Y(u5_mul_69_18_n_1215));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27657 (.A(u5_mul_69_18_n_706),
    .B(u5_mul_69_18_n_187),
    .C(u5_mul_69_18_n_971),
    .Y(u5_mul_69_18_n_1214));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27658 (.A(u5_mul_69_18_n_723),
    .B(u5_mul_69_18_n_208),
    .C(u5_mul_69_18_n_969),
    .Y(u5_mul_69_18_n_1213));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27659 (.A(u5_mul_69_18_n_716),
    .B(u5_mul_69_18_n_181),
    .C(u5_mul_69_18_n_968),
    .Y(u5_mul_69_18_n_1212));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27660 (.A(u5_mul_69_18_n_763),
    .B(u5_mul_69_18_n_667),
    .C(u5_mul_69_18_n_808),
    .Y(u5_mul_69_18_n_1211));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27661 (.A(u5_mul_69_18_n_845),
    .B(u5_mul_69_18_n_205),
    .C(u5_mul_69_18_n_966),
    .Y(u5_mul_69_18_n_1210));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27662 (.A(u5_mul_69_18_n_783),
    .B(u5_mul_69_18_n_666),
    .C(u5_mul_69_18_n_793),
    .Y(u5_mul_69_18_n_1209));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27663 (.A(u5_mul_69_18_n_806),
    .B(u5_mul_69_18_n_664),
    .C(u5_mul_69_18_n_762),
    .Y(u5_mul_69_18_n_1208));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27664 (.A(u5_mul_69_18_n_752),
    .B(u5_mul_69_18_n_668),
    .C(u5_mul_69_18_n_836),
    .Y(u5_mul_69_18_n_1207));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27665 (.A(u5_mul_69_18_n_925),
    .B(u5_mul_69_18_n_946),
    .C(u5_mul_69_18_n_879),
    .Y(u5_mul_69_18_n_1206));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27666 (.A(u5_mul_69_18_n_1003),
    .B(u5_mul_69_18_n_748),
    .C(u5_mul_69_18_n_906),
    .Y(u5_mul_69_18_n_1205));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27667 (.A(u5_mul_69_18_n_945),
    .B(u5_mul_69_18_n_658),
    .C(u5_mul_69_18_n_881),
    .Y(u5_mul_69_18_n_1204));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27668 (.A(u5_mul_69_18_n_937),
    .B(u5_mul_69_18_n_656),
    .C(u5_mul_69_18_n_864),
    .Y(u5_mul_69_18_n_1203));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27669 (.A(u5_mul_69_18_n_754),
    .B(u5_mul_69_18_n_191),
    .C(u5_mul_69_18_n_972),
    .Y(u5_mul_69_18_n_1202));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27670 (.A(u5_mul_69_18_n_910),
    .B(u5_mul_69_18_n_674),
    .C(u5_mul_69_18_n_810),
    .Y(u5_mul_69_18_n_1201));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27671 (.A(u5_mul_69_18_n_928),
    .B(u5_mul_69_18_n_797),
    .C(u5_mul_69_18_n_718),
    .Y(u5_mul_69_18_n_1200));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27672 (.A(u5_mul_69_18_n_911),
    .B(u5_mul_69_18_n_912),
    .C(u5_mul_69_18_n_956),
    .Y(u5_mul_69_18_n_1199));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27673 (.A(u5_mul_69_18_n_792),
    .B(u5_mul_69_18_n_657),
    .C(u5_mul_69_18_n_782),
    .Y(u5_mul_69_18_n_1198));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27674 (.A(u5_mul_69_18_n_871),
    .B(u5_mul_69_18_n_183),
    .C(u5_mul_69_18_n_978),
    .Y(u5_mul_69_18_n_1197));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27675 (.A(u5_mul_69_18_n_697),
    .B(u5_mul_69_18_n_217),
    .C(u5_mul_69_18_n_981),
    .Y(u5_mul_69_18_n_1196));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27676 (.A(u5_mul_69_18_n_694),
    .B(u5_mul_69_18_n_212),
    .C(u5_mul_69_18_n_970),
    .Y(u5_mul_69_18_n_1195));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27677 (.A(u5_mul_69_18_n_711),
    .B(u5_mul_69_18_n_663),
    .C(u5_mul_69_18_n_830),
    .Y(u5_mul_69_18_n_1194));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27678 (.A(u5_mul_69_18_n_802),
    .B(u5_mul_69_18_n_631),
    .C(u5_mul_69_18_n_709),
    .Y(u5_mul_69_18_n_1192));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27679 (.A(u5_mul_69_18_n_913),
    .B(u5_mul_69_18_n_177),
    .C(u5_mul_69_18_n_940),
    .Y(u5_mul_69_18_n_1191));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27680 (.A(u5_mul_69_18_n_900),
    .B(u5_mul_69_18_n_170),
    .C(u5_mul_69_18_n_841),
    .Y(u5_mul_69_18_n_1190));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27681 (.A(u5_mul_69_18_n_914),
    .B(u5_mul_69_18_n_755),
    .C(u5_mul_69_18_n_965),
    .Y(u5_mul_69_18_n_1189));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27682 (.A(u5_mul_69_18_n_701),
    .B(u5_mul_69_18_n_172),
    .C(u5_mul_69_18_n_979),
    .Y(u5_mul_69_18_n_1188));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27683 (.A(u5_mul_69_18_n_787),
    .B(u5_mul_69_18_n_973),
    .C(u5_mul_69_18_n_869),
    .Y(u5_mul_69_18_n_1186));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27687 (.A(u5_mul_69_18_n_1167),
    .Y(u5_mul_69_18_n_1168));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27688 (.A(u5_mul_69_18_n_1126),
    .Y(u5_mul_69_18_n_1127));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27689 (.A(u5_mul_69_18_n_876),
    .B(u5_mul_69_18_n_840),
    .C(u5_mul_69_18_n_923),
    .Y(u5_mul_69_18_n_1176));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27690 (.A(u5_mul_69_18_n_917),
    .B(u5_mul_69_18_n_820),
    .C(u5_mul_69_18_n_728),
    .Y(u5_mul_69_18_n_1175));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27691 (.A(u5_mul_69_18_n_950),
    .B(u5_mul_69_18_n_719),
    .C(u5_mul_69_18_n_875),
    .Y(u5_mul_69_18_n_1174));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27692 (.A(u5_mul_69_18_n_908),
    .B(u5_mul_69_18_n_805),
    .C(u5_mul_69_18_n_758),
    .Y(u5_mul_69_18_n_1173));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27693 (.A(u5_mul_69_18_n_934),
    .B(u5_mul_69_18_n_860),
    .C(u5_mul_69_18_n_873),
    .Y(u5_mul_69_18_n_1172));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27694 (.A(u5_mul_69_18_n_829),
    .B(u5_mul_69_18_n_724),
    .C(u5_mul_69_18_n_727),
    .Y(u5_mul_69_18_n_1171));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27695 (.A(u5_mul_69_18_n_896),
    .B(u5_mul_69_18_n_807),
    .C(u5_mul_69_18_n_768),
    .Y(u5_mul_69_18_n_1170));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27696 (.A(u5_mul_69_18_n_776),
    .B(u5_mul_69_18_n_838),
    .C(u5_mul_69_18_n_712),
    .Y(u5_mul_69_18_n_1169));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27697 (.A(u5_mul_69_18_n_736),
    .B(u5_mul_69_18_n_822),
    .C(u5_mul_69_18_n_904),
    .Y(u5_mul_69_18_n_1167));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27698 (.A(u5_mul_69_18_n_738),
    .B(u5_mul_69_18_n_842),
    .C(u5_mul_69_18_n_740),
    .Y(u5_mul_69_18_n_1166));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27699 (.A(u5_mul_69_18_n_747),
    .B(u5_mul_69_18_n_951),
    .C(u5_mul_69_18_n_730),
    .Y(u5_mul_69_18_n_1165));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27700 (.A(u5_mul_69_18_n_750),
    .B(u5_mul_69_18_n_960),
    .C(u5_mul_69_18_n_903),
    .Y(u5_mul_69_18_n_1164));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27701 (.A(u5_mul_69_18_n_794),
    .B(u5_mul_69_18_n_650),
    .C(u5_mul_69_18_n_714),
    .Y(u5_mul_69_18_n_1163));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27702 (.A(u5_mul_69_18_n_919),
    .B(u5_mul_69_18_n_652),
    .C(u5_mul_69_18_n_831),
    .Y(u5_mul_69_18_n_1162));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27703 (.A(u5_mul_69_18_n_772),
    .B(u5_mul_69_18_n_823),
    .C(u5_mul_69_18_n_846),
    .Y(u5_mul_69_18_n_1161));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27704 (.A(u5_mul_69_18_n_915),
    .B(u5_mul_69_18_n_938),
    .C(u5_mul_69_18_n_894),
    .Y(u5_mul_69_18_n_1160));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27705 (.A(u5_mul_69_18_n_866),
    .B(u5_mul_69_18_n_955),
    .C(u5_mul_69_18_n_870),
    .Y(u5_mul_69_18_n_1159));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27706 (.A(u5_mul_69_18_n_909),
    .B(u5_mul_69_18_n_858),
    .C(u5_mul_69_18_n_954),
    .Y(u5_mul_69_18_n_1158));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27707 (.A(u5_mul_69_18_n_759),
    .B(u5_mul_69_18_n_795),
    .C(u5_mul_69_18_n_761),
    .Y(u5_mul_69_18_n_1157));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27708 (.A(u5_mul_69_18_n_898),
    .B(u5_mul_69_18_n_824),
    .C(u5_mul_69_18_n_767),
    .Y(u5_mul_69_18_n_1156));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27709 (.A(u5_mul_69_18_n_771),
    .B(u5_mul_69_18_n_803),
    .C(u5_mul_69_18_n_769),
    .Y(u5_mul_69_18_n_1155));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27710 (.A(u5_mul_69_18_n_922),
    .B(u5_mul_69_18_n_862),
    .C(u5_mul_69_18_n_939),
    .Y(u5_mul_69_18_n_1154));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27711 (.A(u5_mul_69_18_n_859),
    .B(u5_mul_69_18_n_933),
    .C(u5_mul_69_18_n_861),
    .Y(u5_mul_69_18_n_1153));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27712 (.A(u5_mul_69_18_n_781),
    .B(u5_mul_69_18_n_799),
    .C(u5_mul_69_18_n_892),
    .Y(u5_mul_69_18_n_1152));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27713 (.A(u5_mul_69_18_n_12),
    .B(u5_mul_69_18_n_941),
    .C(u5_mul_69_18_n_720),
    .Y(u5_mul_69_18_n_1151));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27714 (.A(u5_mul_69_18_n_852),
    .B(u5_mul_69_18_n_953),
    .C(u5_mul_69_18_n_854),
    .Y(u5_mul_69_18_n_1150));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27715 (.A(u5_mul_69_18_n_798),
    .B(u5_mul_69_18_n_850),
    .C(u5_mul_69_18_n_778),
    .Y(u5_mul_69_18_n_1149));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27716 (.A(u5_mul_69_18_n_902),
    .B(u5_mul_69_18_n_814),
    .C(u5_mul_69_18_n_746),
    .Y(u5_mul_69_18_n_1148));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27717 (.A(u5_mul_69_18_n_717),
    .B(u5_mul_69_18_n_828),
    .C(u5_mul_69_18_n_713),
    .Y(u5_mul_69_18_n_1147));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27718 (.A(u5_mul_69_18_n_739),
    .B(u5_mul_69_18_n_821),
    .C(u5_mul_69_18_n_734),
    .Y(u5_mul_69_18_n_1146));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27719 (.A(u5_mul_69_18_n_741),
    .B(u5_mul_69_18_n_926),
    .C(u5_mul_69_18_n_819),
    .Y(u5_mul_69_18_n_1145));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27720 (.A(u5_mul_69_18_n_834),
    .B(u5_mul_69_18_n_789),
    .C(u5_mul_69_18_n_742),
    .Y(u5_mul_69_18_n_1144));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27721 (.A(u5_mul_69_18_n_788),
    .B(u5_mul_69_18_n_791),
    .C(u5_mul_69_18_n_743),
    .Y(u5_mul_69_18_n_1143));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27722 (.A(u5_mul_69_18_n_921),
    .B(u5_mul_69_18_n_839),
    .C(u5_mul_69_18_n_882),
    .Y(u5_mul_69_18_n_1142));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27723 (.A(u5_mul_69_18_n_837),
    .B(u5_mul_69_18_n_853),
    .C(u5_mul_69_18_n_849),
    .Y(u5_mul_69_18_n_1141));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27724 (.A(u5_mul_69_18_n_766),
    .B(u5_mul_69_18_n_804),
    .C(u5_mul_69_18_n_770),
    .Y(u5_mul_69_18_n_1140));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27725 (.A(u5_mul_69_18_n_857),
    .B(u5_mul_69_18_n_932),
    .C(u5_mul_69_18_n_856),
    .Y(u5_mul_69_18_n_1139));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27726 (.A(u5_mul_69_18_n_888),
    .B(u5_mul_69_18_n_809),
    .C(u5_mul_69_18_n_729),
    .Y(u5_mul_69_18_n_1138));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27727 (.A(u5_mul_69_18_n_877),
    .B(u5_mul_69_18_n_885),
    .C(u5_mul_69_18_n_817),
    .Y(u5_mul_69_18_n_1137));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27728 (.A(u5_mul_69_18_n_749),
    .B(u5_mul_69_18_n_751),
    .C(u5_mul_69_18_n_816),
    .Y(u5_mul_69_18_n_1136));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27729 (.A(u5_mul_69_18_n_753),
    .B(u5_mul_69_18_n_645),
    .C(u5_mul_69_18_n_796),
    .Y(u5_mul_69_18_n_1135));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27730 (.A(u5_mul_69_18_n_878),
    .B(u5_mul_69_18_n_786),
    .C(u5_mul_69_18_n_942),
    .Y(u5_mul_69_18_n_1134));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27731 (.A(u5_mul_69_18_n_958),
    .B(u5_mul_69_18_n_648),
    .C(u5_mul_69_18_n_924),
    .Y(u5_mul_69_18_n_1133));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27732 (.A(u5_mul_69_18_n_765),
    .B(u5_mul_69_18_n_646),
    .C(u5_mul_69_18_n_943),
    .Y(u5_mul_69_18_n_1132));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27733 (.A(u5_mul_69_18_n_944),
    .B(u5_mul_69_18_n_735),
    .C(u5_mul_69_18_n_733),
    .Y(u5_mul_69_18_n_1131));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27734 (.A(u5_mul_69_18_n_825),
    .B(u5_mul_69_18_n_920),
    .C(u5_mul_69_18_n_732),
    .Y(u5_mul_69_18_n_1130));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27735 (.A(u5_mul_69_18_n_721),
    .B(u5_mul_69_18_n_959),
    .C(u5_mul_69_18_n_722),
    .Y(u5_mul_69_18_n_1129));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27736 (.A(u5_mul_69_18_n_756),
    .B(u5_mul_69_18_n_818),
    .C(u5_mul_69_18_n_726),
    .Y(u5_mul_69_18_n_1128));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27737 (.A(u5_mul_69_18_n_708),
    .B(u5_mul_69_18_n_764),
    .C(u5_mul_69_18_n_832),
    .Y(u5_mul_69_18_n_1126));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27738 (.A(u5_mul_69_18_n_835),
    .B(u5_mul_69_18_n_895),
    .C(u5_mul_69_18_n_774),
    .Y(u5_mul_69_18_n_1125));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27739 (.A(u5_mul_69_18_n_865),
    .B(u5_mul_69_18_n_777),
    .C(u5_mul_69_18_n_949),
    .Y(u5_mul_69_18_n_1124));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27740 (.A(u5_mul_69_18_n_901),
    .B(u5_mul_69_18_n_815),
    .C(u5_mul_69_18_n_715),
    .Y(u5_mul_69_18_n_1123));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27741 (.A(u5_mul_69_18_n_760),
    .B(u5_mul_69_18_n_975),
    .Y(u5_mul_69_18_n_1115));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27742 (.A(u5_mul_69_18_n_985),
    .B(u5_mul_69_18_n_995),
    .Y(u5_mul_69_18_n_1114));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27747 (.A1(u5_mul_69_18_n_184),
    .A2(u5_mul_69_18_n_848),
    .B1(u5_mul_69_18_n_185),
    .B2(u5_mul_69_18_n_847),
    .Y(u5_mul_69_18_n_1109));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27750 (.A(u5_mul_69_18_n_913),
    .B(u5_mul_69_18_n_177),
    .Y(u5_mul_69_18_n_1106));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27752 (.A(u5_mul_69_18_n_844),
    .B(u5_mul_69_18_n_192),
    .Y(u5_mul_69_18_n_1104));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27753 (.A(u5_mul_69_18_n_863),
    .B(u5_mul_69_18_n_169),
    .Y(u5_mul_69_18_n_1103));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27756 (.A(u5_mul_69_18_n_873),
    .B(u5_mul_69_18_n_860),
    .Y(u5_mul_69_18_n_1100));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27759 (.A(u5_mul_69_18_n_699),
    .B(u5_mul_69_18_n_887),
    .Y(u5_mul_69_18_n_1097));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27760 (.A(u5_mul_69_18_n_716),
    .B(u5_mul_69_18_n_181),
    .Y(u5_mul_69_18_n_1096));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27761 (.A(u5_mul_69_18_n_964),
    .B(u5_mul_69_18_n_710),
    .Y(u5_mul_69_18_n_1095));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27762 (.A(u5_mul_69_18_n_982),
    .B(u5_mul_69_18_n_176),
    .Y(u5_mul_69_18_n_1094));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27763 (.A(u5_mul_69_18_n_979),
    .B(u5_mul_69_18_n_172),
    .Y(u5_mul_69_18_n_1093));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27767 (.A1(u5_mul_69_18_n_697),
    .A2(u5_mul_69_18_n_218),
    .B1(u5_mul_69_18_n_698),
    .B2(u5_mul_69_18_n_217),
    .Y(u5_mul_69_18_n_1089));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27768 (.A(u5_mul_69_18_n_754),
    .B(u5_mul_69_18_n_191),
    .Y(u5_mul_69_18_n_1088));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g27771 (.A(u5_mul_69_18_n_985),
    .B(u5_mul_69_18_n_995),
    .Y(u5_mul_69_18_n_1122));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27772 (.A(u5_mul_69_18_n_907),
    .B(u5_mul_69_18_n_214),
    .Y(u5_mul_69_18_n_1085));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27773 (.A(u5_mul_69_18_n_696),
    .B(u5_mul_69_18_n_174),
    .Y(u5_mul_69_18_n_1084));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27777 (.A(u5_mul_69_18_n_983),
    .B(u5_mul_69_18_n_918),
    .Y(u5_mul_69_18_n_1080));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27778 (.A(u5_mul_69_18_n_871),
    .B(u5_mul_69_18_n_183),
    .Y(u5_mul_69_18_n_1079));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27779 (.A1(u5_mul_69_18_n_166),
    .A2(u5_mul_69_18_n_883),
    .B1(u5_mul_69_18_n_167),
    .B2(u5_mul_69_18_n_884),
    .Y(u5_mul_69_18_n_1078));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27786 (.A(u5_mul_69_18_n_901),
    .B(u5_mul_69_18_n_715),
    .Y(u5_mul_69_18_n_1071));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27790 (.A(u5_mul_69_18_n_774),
    .B(u5_mul_69_18_n_895),
    .Y(u5_mul_69_18_n_1067));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27792 (.A(u5_mul_69_18_n_917),
    .B(u5_mul_69_18_n_728),
    .Y(u5_mul_69_18_n_1065));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27794 (.A1(u5_mul_69_18_n_891),
    .A2(u5_mul_69_18_n_843),
    .B(u5_mul_69_18_n_986),
    .Y(u5_mul_69_18_n_1121));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27795 (.A(u5_mul_69_18_n_801),
    .B(u5_mul_69_18_n_682),
    .Y(u5_mul_69_18_n_1120));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27797 (.A(u5_mul_69_18_n_826),
    .B(u5_mul_69_18_n_678),
    .Y(u5_mul_69_18_n_1119));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27798 (.A(u5_mul_69_18_n_947),
    .B(u5_mul_69_18_n_681),
    .Y(u5_mul_69_18_n_1118));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27799 (.A(u5_mul_69_18_n_931),
    .B(u5_mul_69_18_n_685),
    .Y(u5_mul_69_18_n_1117));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27800 (.A(u5_mul_69_18_n_812),
    .B(u5_mul_69_18_n_684),
    .Y(u5_mul_69_18_n_1116));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27802 (.A(u5_mul_69_18_n_846),
    .B(u5_mul_69_18_n_886),
    .Y(u5_mul_69_18_n_1057));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27808 (.A(u5_mul_69_18_n_916),
    .B(u5_mul_69_18_n_962),
    .Y(u5_mul_69_18_n_1051));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27809 (.A(u5_mul_69_18_n_912),
    .B(u5_mul_69_18_n_911),
    .Y(u5_mul_69_18_n_1050));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27811 (.A(u5_mul_69_18_n_804),
    .B(u5_mul_69_18_n_770),
    .Y(u5_mul_69_18_n_1048));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27815 (.A(u5_mul_69_18_n_915),
    .B(u5_mul_69_18_n_894),
    .Y(u5_mul_69_18_n_1044));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27817 (.A(u5_mul_69_18_n_744),
    .B(u5_mul_69_18_n_927),
    .Y(u5_mul_69_18_n_1042));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27818 (.A(u5_mul_69_18_n_772),
    .B(u5_mul_69_18_n_823),
    .Y(u5_mul_69_18_n_1041));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27819 (.A(u5_mul_69_18_n_942),
    .B(u5_mul_69_18_n_878),
    .Y(u5_mul_69_18_n_1040));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27822 (.A(u5_mul_69_18_n_898),
    .B(u5_mul_69_18_n_767),
    .Y(u5_mul_69_18_n_1037));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27823 (.A(u5_mul_69_18_n_747),
    .B(u5_mul_69_18_n_730),
    .Y(u5_mul_69_18_n_1036));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27824 (.A(u5_mul_69_18_n_727),
    .B(u5_mul_69_18_n_724),
    .Y(u5_mul_69_18_n_1035));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27825 (.A(u5_mul_69_18_n_922),
    .B(u5_mul_69_18_n_862),
    .Y(u5_mul_69_18_n_1034));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27827 (.A(u5_mul_69_18_n_945),
    .B(u5_mul_69_18_n_881),
    .Y(u5_mul_69_18_n_1032));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27830 (.A(u5_mul_69_18_n_859),
    .B(u5_mul_69_18_n_861),
    .Y(u5_mul_69_18_n_1029));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27832 (.A(u5_mul_69_18_n_950),
    .B(u5_mul_69_18_n_719),
    .Y(u5_mul_69_18_n_1027));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27833 (.A(u5_mul_69_18_n_713),
    .B(u5_mul_69_18_n_828),
    .Y(u5_mul_69_18_n_1026));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27835 (.A(u5_mul_69_18_n_832),
    .B(u5_mul_69_18_n_708),
    .Y(u5_mul_69_18_n_1024));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27836 (.A(u5_mul_69_18_n_725),
    .B(u5_mul_69_18_n_779),
    .Y(u5_mul_69_18_n_1023));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27839 (.A(u5_mul_69_18_n_783),
    .B(u5_mul_69_18_n_793),
    .Y(u5_mul_69_18_n_1020));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27845 (.A(u5_mul_69_18_n_763),
    .B(u5_mul_69_18_n_808),
    .Y(u5_mul_69_18_n_1014));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27847 (.A(u5_mul_69_18_n_745),
    .B(u5_mul_69_18_n_929),
    .Y(u5_mul_69_18_n_1012));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27850 (.A(u5_mul_69_18_n_738),
    .B(u5_mul_69_18_n_740),
    .Y(u5_mul_69_18_n_1009));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27851 (.A(u5_mul_69_18_n_759),
    .B(u5_mul_69_18_n_761),
    .Y(u5_mul_69_18_n_1008));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27856 (.A(u5_mul_69_18_n_952),
    .B(u5_mul_69_18_n_653),
    .C(u5_mul_69_18_n_660),
    .Y(u5_mul_69_18_n_1063));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27857 (.A(u5_mul_69_18_n_936),
    .B(u5_mul_69_18_n_649),
    .C(u5_mul_69_18_n_659),
    .Y(u5_mul_69_18_n_1062));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27858 (.A(u5_mul_69_18_n_935),
    .B(u5_mul_69_18_n_647),
    .C(u5_mul_69_18_n_675),
    .Y(u5_mul_69_18_n_1061));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g27859 (.A(u5_mul_69_18_n_800),
    .B(u5_mul_69_18_n_651),
    .C(u5_mul_69_18_n_677),
    .Y(u5_mul_69_18_n_1060));
 MAJx2_ASAP7_75t_R u5_mul_69_18_g27860 (.A(u5_mul_69_18_n_811),
    .B(u5_mul_69_18_n_654),
    .C(u5_mul_69_18_n_662),
    .Y(u5_mul_69_18_n_1059));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27862 (.A1(u5_mul_69_18_n_673),
    .A2(u5_mul_69_18_n_655),
    .B(u5_mul_69_18_n_986),
    .Y(u5_mul_69_18_n_996));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27863 (.A(u5_mul_69_18_n_684),
    .B(u5_mul_69_18_n_813),
    .Y(u5_mul_69_18_n_1003));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27864 (.A(u5_mul_69_18_n_680),
    .B(u5_mul_69_18_n_833),
    .Y(u5_mul_69_18_n_1002));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27865 (.A(u5_mul_69_18_n_678),
    .B(u5_mul_69_18_n_827),
    .Y(u5_mul_69_18_n_1001));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27866 (.A(u5_mul_69_18_n_681),
    .B(u5_mul_69_18_n_948),
    .Y(u5_mul_69_18_n_1000));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27867 (.A(u5_mul_69_18_n_685),
    .B(u5_mul_69_18_n_931),
    .Y(u5_mul_69_18_n_999));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27868 (.A(u5_mul_69_18_n_682),
    .B(u5_mul_69_18_n_801),
    .Y(u5_mul_69_18_n_998));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27872 (.A(u5_mul_69_18_n_671),
    .B(u5_mul_69_18_n_686),
    .Y(u5_mul_69_18_n_995));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27874 (.A(u5_mul_69_18_n_670),
    .B(u5_mul_69_18_n_689),
    .Y(u5_mul_69_18_n_994));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g27875 (.A(u5_mul_69_18_n_672),
    .B(u5_mul_69_18_n_688),
    .Y(u5_mul_69_18_n_993));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27876 (.A(u5_mul_69_18_n_679),
    .B(u5_mul_69_18_n_683),
    .Y(u5_mul_69_18_n_992));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g27877 (.A(u5_mul_69_18_n_669),
    .B(u5_mul_69_18_n_687),
    .Y(u5_mul_69_18_n_991));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27879 (.A(u5_mul_69_18_n_947),
    .Y(u5_mul_69_18_n_948));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27880 (.A(u5_mul_69_18_n_883),
    .Y(u5_mul_69_18_n_884));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27881 (.A(u5_mul_69_18_n_867),
    .Y(u5_mul_69_18_n_868));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g27882 (.A(u5_mul_69_18_n_848),
    .Y(u5_mul_69_18_n_847));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27883 (.A1(u5_mul_69_18_n_423),
    .A2(u5_mul_69_18_n_634),
    .B(u5_mul_69_18_n_149),
    .Y(u5_mul_69_18_n_844));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27884 (.A(u5_mul_69_18_n_655),
    .B(u5_mul_69_18_n_673),
    .Y(u5_mul_69_18_n_986));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27886 (.A1(u5_mul_69_18_n_221),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_509),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_985));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27887 (.A(u5_mul_69_18_n_686),
    .B(u5_mul_69_18_n_671),
    .Y(u5_mul_69_18_n_984));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27888 (.A1(u5_mul_69_18_n_585),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_607),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_983));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27889 (.A1(u5_mul_69_18_n_592),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_594),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_982));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27890 (.A1(u5_mul_69_18_n_599),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_603),
    .B2(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_981));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27891 (.A1(u5_mul_69_18_n_593),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_590),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_980));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27892 (.A1(u5_mul_69_18_n_600),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_605),
    .B2(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_979));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27893 (.A1(u5_mul_69_18_n_597),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_589),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_978));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27894 (.A1(u5_mul_69_18_n_602),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_604),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_977));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27895 (.A1(u5_mul_69_18_n_604),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_591),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_976));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27896 (.A1(u5_mul_69_18_n_595),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_593),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_975));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27897 (.A1(u5_mul_69_18_n_606),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_592),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_974));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27898 (.A1(u5_mul_69_18_n_586),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_602),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_973));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27899 (.A1(u5_mul_69_18_n_603),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_588),
    .B2(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_972));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27900 (.A1(u5_mul_69_18_n_590),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_597),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_971));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27901 (.A1(u5_mul_69_18_n_587),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_595),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_970));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27902 (.A1(u5_mul_69_18_n_594),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_586),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_969));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27903 (.A1(u5_mul_69_18_n_601),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_5),
    .B2(u5_mul_69_18_n_599),
    .Y(u5_mul_69_18_n_968));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27904 (.A1(u5_mul_69_18_n_605),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_606),
    .B2(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_967));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27905 (.A1(u5_mul_69_18_n_598),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_585),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_966));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27906 (.A1(u5_mul_69_18_n_379),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_47),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_965));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27907 (.A1(u5_mul_69_18_n_274),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_83),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_964));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27908 (.A1(u5_mul_69_18_n_639),
    .A2(u5_mul_69_18_n_343),
    .B1(u5_mul_69_18_n_431),
    .B2(u5_mul_69_18_n_78),
    .Y(u5_mul_69_18_n_963));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27909 (.A1(u5_mul_69_18_n_223),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_503),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_962));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27910 (.A1(u5_mul_69_18_n_227),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_435),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_961));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27911 (.A1(u5_mul_69_18_n_495),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_479),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_960));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27912 (.A1(u5_mul_69_18_n_219),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_297),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_959));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27913 (.A1(u5_mul_69_18_n_369),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_271),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_958));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27914 (.A1(u5_mul_69_18_n_237),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_424),
    .B2(u5_mul_69_18_n_541),
    .Y(u5_mul_69_18_n_957));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27915 (.A(u5_mul_69_18_n_683),
    .B(u5_mul_69_18_n_679),
    .Y(u5_mul_69_18_n_956));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27916 (.A1(u5_mul_69_18_n_565),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_459),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_955));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27917 (.A1(u5_mul_69_18_n_514),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_535),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_954));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27918 (.A1(u5_mul_69_18_n_644),
    .A2(u5_mul_69_18_n_374),
    .B1(u5_mul_69_18_n_2),
    .B2(u5_mul_69_18_n_440),
    .Y(u5_mul_69_18_n_953));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27919 (.A1(u5_mul_69_18_n_508),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_7),
    .B2(u5_mul_69_18_n_347),
    .Y(u5_mul_69_18_n_952));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27920 (.A1(u5_mul_69_18_n_524),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_532),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_951));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27921 (.A1(u5_mul_69_18_n_624),
    .A2(u5_mul_69_18_n_515),
    .B1(u5_mul_69_18_n_6),
    .B2(u5_mul_69_18_n_490),
    .Y(u5_mul_69_18_n_950));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27922 (.A1(u5_mul_69_18_n_419),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_485),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_949));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27923 (.A1(u5_mul_69_18_n_463),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_368),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_947));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27924 (.A1(u5_mul_69_18_n_464),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_316),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_946));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27925 (.A1(u5_mul_69_18_n_322),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_282),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_945));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27926 (.A1(u5_mul_69_18_n_234),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_292),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_944));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27927 (.A1(u5_mul_69_18_n_478),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_510),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_943));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27928 (.A1(u5_mul_69_18_n_544),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_378),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_942));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27929 (.A1(u5_mul_69_18_n_314),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_520),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_941));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27930 (.A1(u5_mul_69_18_n_547),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_567),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_940));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27931 (.A1(u5_mul_69_18_n_283),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_494),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_939));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27932 (.A1(u5_mul_69_18_n_549),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_563),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_938));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27933 (.A1(u5_mul_69_18_n_530),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_534),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_937));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27934 (.A1(u5_mul_69_18_n_318),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_493),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_936));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27935 (.A1(u5_mul_69_18_n_458),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_550),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_935));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27936 (.A1(u5_mul_69_18_n_457),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_338),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_934));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27937 (.A1(u5_mul_69_18_n_450),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_522),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_933));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27938 (.A1(u5_mul_69_18_n_442),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_359),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_932));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27939 (.A1(u5_mul_69_18_n_284),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_477),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_931));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27940 (.A1(u5_mul_69_18_n_7),
    .A2(u5_mul_69_18_n_622),
    .B(u5_mul_69_18_n_91),
    .Y(u5_mul_69_18_n_930));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27941 (.A1(u5_mul_69_18_n_220),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_489),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_929));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27942 (.A(u5_mul_69_18_n_687),
    .B(u5_mul_69_18_n_669),
    .Y(u5_mul_69_18_n_928));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27943 (.A1(u5_mul_69_18_n_222),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_517),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_927));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27944 (.A1(u5_mul_69_18_n_226),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_11),
    .B2(u5_mul_69_18_n_443),
    .Y(u5_mul_69_18_n_926));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27945 (.A1(u5_mul_69_18_n_625),
    .A2(u5_mul_69_18_n_424),
    .B(u5_mul_69_18_n_45),
    .Y(u5_mul_69_18_n_925));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27946 (.A1(u5_mul_69_18_n_447),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_277),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_924));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27947 (.A1(u5_mul_69_18_n_640),
    .A2(u5_mul_69_18_n_11),
    .B(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_923));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27948 (.A1(u5_mul_69_18_n_562),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_551),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_922));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27949 (.A1(u5_mul_69_18_n_406),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_235),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_921));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27950 (.A1(u5_mul_69_18_n_498),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_242),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_920));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27951 (.A1(u5_mul_69_18_n_564),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_413),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_919));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27952 (.A1(u5_mul_69_18_n_427),
    .A2(u5_mul_69_18_n_641),
    .B(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_918));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27953 (.A1(u5_mul_69_18_n_421),
    .A2(u5_mul_69_18_n_637),
    .B(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_917));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27954 (.A1(u5_mul_69_18_n_550),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_447),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_916));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27955 (.A1(u5_mul_69_18_n_351),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_559),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_915));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27956 (.A1(u5_mul_69_18_n_488),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_371),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_914));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27957 (.A1(u5_mul_69_18_n_494),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_470),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_913));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27958 (.A1(u5_mul_69_18_n_536),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_396),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_912));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27959 (.A1(u5_mul_69_18_n_484),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_463),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_911));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27960 (.A1(u5_mul_69_18_n_534),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_302),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_910));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27961 (.A1(u5_mul_69_18_n_561),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_483),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_909));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27962 (.A1(u5_mul_69_18_n_70),
    .A2(u5_mul_69_18_n_71),
    .B(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_908));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27963 (.A1(u5_mul_69_18_n_588),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_600),
    .B2(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_907));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27964 (.A1(u5_mul_69_18_n_352),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_583),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_906));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27965 (.A1(u5_mul_69_18_n_436),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_513),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_905));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27966 (.A1(u5_mul_69_18_n_572),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_380),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_904));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27967 (.A1(u5_mul_69_18_n_348),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_358),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_903));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27968 (.A1(u5_mul_69_18_n_287),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_434),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_902));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27969 (.A1(u5_mul_69_18_n_425),
    .A2(u5_mul_69_18_n_623),
    .B(u5_mul_69_18_n_61),
    .Y(u5_mul_69_18_n_901));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27970 (.A1(u5_mul_69_18_n_420),
    .A2(u5_mul_69_18_n_643),
    .B(u5_mul_69_18_n_63),
    .Y(u5_mul_69_18_n_900));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27971 (.A1(u5_mul_69_18_n_480),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_344),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_899));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27972 (.A1(u5_mul_69_18_n_438),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_545),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_898));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27973 (.A1(u5_mul_69_18_n_281),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_320),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_897));
 AOI21xp33_ASAP7_75t_R u5_mul_69_18_g27974 (.A1(u5_mul_69_18_n_429),
    .A2(u5_mul_69_18_n_627),
    .B(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_896));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g27975 (.A1(u5_mul_69_18_n_430),
    .A2(u5_mul_69_18_n_629),
    .B(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_895));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27976 (.A1(u5_mul_69_18_n_552),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_386),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_894));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27977 (.A1(u5_mul_69_18_n_441),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_448),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_893));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27978 (.A1(u5_mul_69_18_n_439),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_384),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_892));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27979 (.A(u5_mul_69_18_n_584),
    .B(u5_mul_69_18_n_690),
    .Y(u5_mul_69_18_n_891));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27980 (.A1(u5_mul_69_18_n_396),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_424),
    .B2(u5_mul_69_18_n_237),
    .Y(u5_mul_69_18_n_890));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27981 (.A1(u5_mul_69_18_n_504),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_414),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_889));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27982 (.A1(u5_mul_69_18_n_298),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_562),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_888));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27983 (.A1(u5_mul_69_18_n_589),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_598),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_887));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27984 (.A1(u5_mul_69_18_n_303),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_335),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_886));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27985 (.A1(u5_mul_69_18_n_468),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_546),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_885));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27986 (.A1(u5_mul_69_18_n_607),
    .A2(u5_mul_69_18_n_32),
    .B1(u5_mul_69_18_n_150),
    .B2(u5_mul_69_18_n_30),
    .Y(u5_mul_69_18_n_883));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27987 (.A1(u5_mul_69_18_n_278),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_321),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_882));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27988 (.A1(u5_mul_69_18_n_399),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_361),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_881));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27989 (.A1(u5_mul_69_18_n_497),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_61),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_880));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27990 (.A1(u5_mul_69_18_n_317),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_500),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_879));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27991 (.A1(u5_mul_69_18_n_499),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_349),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_878));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27992 (.A1(u5_mul_69_18_n_405),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_351),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_877));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27993 (.A1(u5_mul_69_18_n_624),
    .A2(u5_mul_69_18_n_569),
    .B1(u5_mul_69_18_n_6),
    .B2(u5_mul_69_18_n_496),
    .Y(u5_mul_69_18_n_876));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27994 (.A1(u5_mul_69_18_n_629),
    .A2(u5_mul_69_18_n_528),
    .B1(u5_mul_69_18_n_430),
    .B2(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_875));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27995 (.A1(u5_mul_69_18_n_596),
    .A2(u5_mul_69_18_n_632),
    .B1(u5_mul_69_18_n_5),
    .B2(u5_mul_69_18_n_601),
    .Y(u5_mul_69_18_n_874));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g27996 (.A1(u5_mul_69_18_n_324),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_73),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_873));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g27997 (.A(u5_mul_69_18_n_689),
    .B(u5_mul_69_18_n_670),
    .Y(u5_mul_69_18_n_872));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27998 (.A1(u5_mul_69_18_n_367),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_63),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_871));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g27999 (.A1(u5_mul_69_18_n_581),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_279),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_870));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28000 (.A1(u5_mul_69_18_n_292),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_58),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_869));
 OAI32xp33_ASAP7_75t_R u5_mul_69_18_g28001 (.A1(u5_mul_69_18_n_632),
    .A2(u5_mul_69_18_n_177),
    .A3(u5_mul_69_18_n_163),
    .B1(u5_mul_69_18_n_5),
    .B2(u5_mul_69_18_n_596),
    .Y(u5_mul_69_18_n_867));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28002 (.A1(u5_mul_69_18_n_525),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_304),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_866));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28003 (.A1(u5_mul_69_18_n_521),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_50),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_865));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28004 (.A1(u5_mul_69_18_n_523),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_3),
    .B2(u5_mul_69_18_n_548),
    .Y(u5_mul_69_18_n_864));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28005 (.A1(u5_mul_69_18_n_591),
    .A2(u5_mul_69_18_n_633),
    .B1(u5_mul_69_18_n_587),
    .B2(u5_mul_69_18_n_422),
    .Y(u5_mul_69_18_n_863));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28006 (.A1(u5_mul_69_18_n_487),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_565),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_862));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28008 (.A1(u5_mul_69_18_n_452),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_281),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_861));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28009 (.A1(u5_mul_69_18_n_359),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_240),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_860));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28010 (.A1(u5_mul_69_18_n_451),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_529),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_859));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28011 (.A1(u5_mul_69_18_n_225),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_458),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_858));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28012 (.A1(u5_mul_69_18_n_402),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_457),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_857));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28013 (.A1(u5_mul_69_18_n_636),
    .A2(u5_mul_69_18_n_445),
    .B1(u5_mul_69_18_n_428),
    .B2(u5_mul_69_18_n_324),
    .Y(u5_mul_69_18_n_856));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28014 (.A(u5_mul_69_18_n_688),
    .B(u5_mul_69_18_n_672),
    .Y(u5_mul_69_18_n_855));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28015 (.A1(u5_mul_69_18_n_556),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_306),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_854));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28016 (.A1(u5_mul_69_18_n_479),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_397),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_853));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28017 (.A1(u5_mul_69_18_n_434),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_437),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_852));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28018 (.A1(u5_mul_69_18_n_228),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_3),
    .B2(u5_mul_69_18_n_449),
    .Y(u5_mul_69_18_n_851));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28019 (.A1(u5_mul_69_18_n_229),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_420),
    .B2(u5_mul_69_18_n_516),
    .Y(u5_mul_69_18_n_850));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28020 (.A1(u5_mul_69_18_n_334),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_527),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_849));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28021 (.A1(u5_mul_69_18_n_316),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_531),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_848));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28022 (.A1(u5_mul_69_18_n_403),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_512),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_846));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28023 (.A1(u5_mul_69_18_n_557),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_142),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_845));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28025 (.A(u5_mul_69_18_n_826),
    .Y(u5_mul_69_18_n_827));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28026 (.A(u5_mul_69_18_n_693),
    .Y(u5_mul_69_18_n_825));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28027 (.A(u5_mul_69_18_n_692),
    .Y(u5_mul_69_18_n_820));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28028 (.A(u5_mul_69_18_n_812),
    .Y(u5_mul_69_18_n_813));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28029 (.A(u5_mul_69_18_n_691),
    .Y(u5_mul_69_18_n_724));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28030 (.A(u5_mul_69_18_n_705),
    .Y(u5_mul_69_18_n_704));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28031 (.A(u5_mul_69_18_n_703),
    .Y(u5_mul_69_18_n_702));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28032 (.A(u5_mul_69_18_n_700),
    .Y(u5_mul_69_18_n_701));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28033 (.A(u5_mul_69_18_n_698),
    .Y(u5_mul_69_18_n_697));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28034 (.A(u5_mul_69_18_n_694),
    .Y(u5_mul_69_18_n_695));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28035 (.A1(u5_mul_69_18_n_446),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_539),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_842));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28036 (.A1(u5_mul_69_18_n_641),
    .A2(u5_mul_69_18_n_395),
    .B1(u5_mul_69_18_n_427),
    .B2(u5_mul_69_18_n_557),
    .Y(u5_mul_69_18_n_841));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28037 (.A1(u5_mul_69_18_n_578),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_481),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_840));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28038 (.A1(u5_mul_69_18_n_432),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_399),
    .B2(u5_mul_69_18_n_29),
    .Y(u5_mul_69_18_n_839));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28039 (.A1(u5_mul_69_18_n_568),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_446),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_838));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28040 (.A1(u5_mul_69_18_n_575),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_515),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_837));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28041 (.A1(u5_mul_69_18_n_411),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_474),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_836));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28042 (.A1(u5_mul_69_18_n_490),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_511),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_835));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28043 (.A1(u5_mul_69_18_n_580),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_402),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_834));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28044 (.A1(u5_mul_69_18_n_271),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_564),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_833));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28045 (.A1(u5_mul_69_18_n_276),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_363),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_832));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28046 (.A1(u5_mul_69_18_n_462),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_288),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_831));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28047 (.A1(u5_mul_69_18_n_517),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_286),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_830));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28048 (.A1(u5_mul_69_18_n_626),
    .A2(u5_mul_69_18_n_296),
    .B1(u5_mul_69_18_n_1),
    .B2(u5_mul_69_18_n_577),
    .Y(u5_mul_69_18_n_829));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28049 (.A1(u5_mul_69_18_n_307),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_2),
    .B2(u5_mul_69_18_n_452),
    .Y(u5_mul_69_18_n_828));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28050 (.A1(u5_mul_69_18_n_510),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_581),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_826));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28051 (.A1(u5_mul_69_18_n_302),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_419),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_693));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28052 (.A1(u5_mul_69_18_n_500),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_499),
    .B2(u5_mul_69_18_n_31),
    .Y(u5_mul_69_18_n_824));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28053 (.A1(u5_mul_69_18_n_387),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_370),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_823));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28054 (.A1(u5_mul_69_18_n_486),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_543),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_822));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28055 (.A1(u5_mul_69_18_n_236),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_284),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_821));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28056 (.A1(u5_mul_69_18_n_358),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_303),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_692));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28057 (.A1(u5_mul_69_18_n_326),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_289),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_819));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28058 (.A1(u5_mul_69_18_n_401),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_356),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_818));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28059 (.A1(u5_mul_69_18_n_628),
    .A2(u5_mul_69_18_n_361),
    .B1(u5_mul_69_18_n_0),
    .B2(u5_mul_69_18_n_526),
    .Y(u5_mul_69_18_n_817));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28060 (.A1(u5_mul_69_18_n_381),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_315),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_816));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28061 (.A1(u5_mul_69_18_n_641),
    .A2(u5_mul_69_18_n_345),
    .B1(u5_mul_69_18_n_427),
    .B2(u5_mul_69_18_n_409),
    .Y(u5_mul_69_18_n_815));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28062 (.A1(u5_mul_69_18_n_385),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_464),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_814));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28063 (.A1(u5_mul_69_18_n_476),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_346),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_812));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28064 (.A1(u5_mul_69_18_n_453),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_354),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_811));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28065 (.A1(u5_mul_69_18_n_320),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_498),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_810));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28066 (.A1(u5_mul_69_18_n_469),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_468),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_809));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28067 (.A1(u5_mul_69_18_n_461),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_388),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_808));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28068 (.A1(u5_mul_69_18_n_629),
    .A2(u5_mul_69_18_n_364),
    .B1(u5_mul_69_18_n_430),
    .B2(u5_mul_69_18_n_342),
    .Y(u5_mul_69_18_n_807));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28069 (.A1(u5_mul_69_18_n_460),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_406),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_806));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28070 (.A1(u5_mul_69_18_n_531),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_329),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_805));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28071 (.A1(u5_mul_69_18_n_241),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_473),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_804));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28072 (.A1(u5_mul_69_18_n_233),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_439),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_803));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28073 (.A1(u5_mul_69_18_n_386),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_560),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_802));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28074 (.A1(u5_mul_69_18_n_315),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_465),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_801));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28075 (.A1(u5_mul_69_18_n_553),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_561),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_800));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28076 (.A1(u5_mul_69_18_n_482),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_506),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_799));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28077 (.A1(u5_mul_69_18_n_537),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_352),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_798));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28078 (.A1(u5_mul_69_18_n_297),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_8),
    .B2(u5_mul_69_18_n_554),
    .Y(u5_mul_69_18_n_797));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28079 (.A1(u5_mul_69_18_n_346),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_433),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_796));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28080 (.A1(u5_mul_69_18_n_301),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_385),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_795));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28081 (.A1(u5_mul_69_18_n_340),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_393),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_794));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28082 (.A1(u5_mul_69_18_n_466),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_416),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_793));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28083 (.A1(u5_mul_69_18_n_375),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_571),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_792));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28084 (.A1(u5_mul_69_18_n_384),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_236),
    .B2(u5_mul_69_18_n_31),
    .Y(u5_mul_69_18_n_791));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28085 (.A1(u5_mul_69_18_n_415),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_291),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_790));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28086 (.A1(u5_mul_69_18_n_473),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_374),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_789));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28087 (.A1(u5_mul_69_18_n_391),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_460),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_788));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28088 (.A1(u5_mul_69_18_n_505),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_574),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_787));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28089 (.A1(u5_mul_69_18_n_240),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_472),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_786));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28090 (.A1(u5_mul_69_18_n_347),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_553),
    .B2(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_785));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28091 (.A1(u5_mul_69_18_n_273),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_491),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_784));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28092 (.A1(u5_mul_69_18_n_622),
    .A2(u5_mul_69_18_n_570),
    .B1(u5_mul_69_18_n_7),
    .B2(u5_mul_69_18_n_331),
    .Y(u5_mul_69_18_n_783));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28093 (.A1(u5_mul_69_18_n_389),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_467),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_782));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28094 (.A1(u5_mul_69_18_n_383),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_390),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_781));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28095 (.A1(u5_mul_69_18_n_299),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_578),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_780));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28096 (.A1(u5_mul_69_18_n_448),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_412),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_779));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28097 (.A1(u5_mul_69_18_n_507),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_8),
    .B2(u5_mul_69_18_n_418),
    .Y(u5_mul_69_18_n_778));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28098 (.A1(u5_mul_69_18_n_242),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_241),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_777));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28099 (.A1(u5_mul_69_18_n_305),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_501),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_776));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28100 (.A1(u5_mul_69_18_n_293),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_287),
    .B2(u5_mul_69_18_n_29),
    .Y(u5_mul_69_18_n_775));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28101 (.A1(u5_mul_69_18_n_512),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_343),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_774));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28102 (.A1(u5_mul_69_18_n_489),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_538),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_773));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28103 (.A1(u5_mul_69_18_n_336),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_299),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_772));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28104 (.A1(u5_mul_69_18_n_337),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_382),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_771));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28105 (.A1(u5_mul_69_18_n_357),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_231),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_770));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28106 (.A1(u5_mul_69_18_n_355),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_375),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_769));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28107 (.A1(u5_mul_69_18_n_639),
    .A2(u5_mul_69_18_n_519),
    .B1(u5_mul_69_18_n_431),
    .B2(u5_mul_69_18_n_372),
    .Y(u5_mul_69_18_n_768));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28108 (.A1(u5_mul_69_18_n_306),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_492),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_767));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28109 (.A1(u5_mul_69_18_n_626),
    .A2(u5_mul_69_18_n_377),
    .B1(u5_mul_69_18_n_1),
    .B2(u5_mul_69_18_n_274),
    .Y(u5_mul_69_18_n_766));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28110 (.A1(u5_mul_69_18_n_235),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_404),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_765));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28111 (.A1(u5_mul_69_18_n_412),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_555),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_764));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28112 (.A1(u5_mul_69_18_n_365),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_340),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_763));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28113 (.A1(u5_mul_69_18_n_417),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_411),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_762));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28114 (.A1(u5_mul_69_18_n_360),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_319),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_761));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28115 (.A1(u5_mul_69_18_n_408),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_323),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_760));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28116 (.A1(u5_mul_69_18_n_558),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_333),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_759));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28117 (.A1(u5_mul_69_18_n_629),
    .A2(u5_mul_69_18_n_492),
    .B1(u5_mul_69_18_n_430),
    .B2(u5_mul_69_18_n_275),
    .Y(u5_mul_69_18_n_758));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28118 (.A1(u5_mul_69_18_n_370),
    .A2(u5_mul_69_18_n_644),
    .B1(u5_mul_69_18_n_407),
    .B2(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_757));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28119 (.A1(u5_mul_69_18_n_311),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_376),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_756));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28120 (.A1(u5_mul_69_18_n_471),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_353),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_755));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28121 (.A1(u5_mul_69_18_n_485),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_579),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_754));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28122 (.A1(u5_mul_69_18_n_332),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_278),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_753));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28123 (.A1(u5_mul_69_18_n_573),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_298),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_752));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28124 (.A1(u5_mul_69_18_n_444),
    .A2(u5_mul_69_18_n_639),
    .B1(u5_mul_69_18_n_461),
    .B2(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_751));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28125 (.A1(u5_mul_69_18_n_373),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_239),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_750));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28126 (.A1(u5_mul_69_18_n_290),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_365),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_749));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28127 (.A1(u5_mul_69_18_n_516),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_420),
    .B2(u5_mul_69_18_n_308),
    .Y(u5_mul_69_18_n_748));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28128 (.A1(u5_mul_69_18_n_566),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_337),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_747));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28129 (.A1(u5_mul_69_18_n_455),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_556),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_746));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28130 (.A1(u5_mul_69_18_n_533),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_482),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_745));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28131 (.A1(u5_mul_69_18_n_542),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_272),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_744));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28132 (.A1(u5_mul_69_18_n_392),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_230),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_743));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28133 (.A1(u5_mul_69_18_n_333),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_445),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_742));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28134 (.A1(u5_mul_69_18_n_493),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_453),
    .B2(u5_mul_69_18_n_28),
    .Y(u5_mul_69_18_n_741));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28135 (.A1(u5_mul_69_18_n_456),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_360),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_740));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28136 (.A1(u5_mul_69_18_n_230),
    .A2(u5_mul_69_18_n_71),
    .B1(u5_mul_69_18_n_573),
    .B2(u5_mul_69_18_n_70),
    .Y(u5_mul_69_18_n_739));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28137 (.A1(u5_mul_69_18_n_560),
    .A2(u5_mul_69_18_n_636),
    .B1(u5_mul_69_18_n_558),
    .B2(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_738));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28138 (.A1(u5_mul_69_18_n_635),
    .A2(u5_mul_69_18_n_277),
    .B1(u5_mul_69_18_n_9),
    .B2(u5_mul_69_18_n_462),
    .Y(u5_mul_69_18_n_737));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28139 (.A1(u5_mul_69_18_n_576),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_566),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_736));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28140 (.A1(u5_mul_69_18_n_353),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_348),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_735));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28141 (.A1(u5_mul_69_18_n_418),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_609),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_734));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28142 (.A1(u5_mul_69_18_n_555),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_495),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_733));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28143 (.A1(u5_mul_69_18_n_563),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_400),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_732));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28144 (.A1(u5_mul_69_18_n_554),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_524),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_731));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28145 (.A1(u5_mul_69_18_n_543),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_232),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_730));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28146 (.A1(u5_mul_69_18_n_474),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_11),
    .B2(u5_mul_69_18_n_487),
    .Y(u5_mul_69_18_n_729));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28147 (.A1(u5_mul_69_18_n_639),
    .A2(u5_mul_69_18_n_238),
    .B1(u5_mul_69_18_n_431),
    .B2(u5_mul_69_18_n_403),
    .Y(u5_mul_69_18_n_728));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28148 (.A1(u5_mul_69_18_n_310),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_325),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_727));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28149 (.A1(u5_mul_69_18_n_362),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_300),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_726));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28150 (.A1(u5_mul_69_18_n_339),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_488),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_725));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28151 (.A1(u5_mul_69_18_n_520),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_572),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_691));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28152 (.A1(u5_mul_69_18_n_371),
    .A2(u5_mul_69_18_n_623),
    .B1(u5_mul_69_18_n_505),
    .B2(u5_mul_69_18_n_425),
    .Y(u5_mul_69_18_n_723));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28153 (.A1(u5_mul_69_18_n_285),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_309),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_722));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28154 (.A1(u5_mul_69_18_n_491),
    .A2(u5_mul_69_18_n_625),
    .B1(u5_mul_69_18_n_295),
    .B2(u5_mul_69_18_n_424),
    .Y(u5_mul_69_18_n_721));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28155 (.A1(u5_mul_69_18_n_413),
    .A2(u5_mul_69_18_n_622),
    .B1(u5_mul_69_18_n_318),
    .B2(u5_mul_69_18_n_28),
    .Y(u5_mul_69_18_n_720));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28156 (.A1(u5_mul_69_18_n_644),
    .A2(u5_mul_69_18_n_398),
    .B1(u5_mul_69_18_n_2),
    .B2(u5_mul_69_18_n_387),
    .Y(u5_mul_69_18_n_719));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28157 (.A1(u5_mul_69_18_n_309),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_486),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_718));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28158 (.A1(u5_mul_69_18_n_582),
    .A2(u5_mul_69_18_n_624),
    .B1(u5_mul_69_18_n_451),
    .B2(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_717));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28159 (.A1(u5_mul_69_18_n_470),
    .A2(u5_mul_69_18_n_621),
    .B1(u5_mul_69_18_n_521),
    .B2(u5_mul_69_18_n_426),
    .Y(u5_mul_69_18_n_716));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28160 (.A1(u5_mul_69_18_n_644),
    .A2(u5_mul_69_18_n_328),
    .B1(u5_mul_69_18_n_2),
    .B2(u5_mul_69_18_n_366),
    .Y(u5_mul_69_18_n_715));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28161 (.A1(u5_mul_69_18_n_465),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_475),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_714));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28162 (.A1(u5_mul_69_18_n_608),
    .A2(u5_mul_69_18_n_629),
    .B1(u5_mul_69_18_n_469),
    .B2(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_713));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28163 (.A1(u5_mul_69_18_n_280),
    .A2(u5_mul_69_18_n_638),
    .B1(u5_mul_69_18_n_456),
    .B2(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_712));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28164 (.A1(u5_mul_69_18_n_291),
    .A2(u5_mul_69_18_n_628),
    .B1(u5_mul_69_18_n_313),
    .B2(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_711));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28165 (.A1(u5_mul_69_18_n_231),
    .A2(u5_mul_69_18_n_641),
    .B1(u5_mul_69_18_n_442),
    .B2(u5_mul_69_18_n_427),
    .Y(u5_mul_69_18_n_710));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28166 (.A1(u5_mul_69_18_n_459),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_362),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_709));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28167 (.A1(u5_mul_69_18_n_330),
    .A2(u5_mul_69_18_n_640),
    .B1(u5_mul_69_18_n_518),
    .B2(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_708));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28168 (.A1(u5_mul_69_18_n_540),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_454),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_707));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28169 (.A1(u5_mul_69_18_n_323),
    .A2(u5_mul_69_18_n_643),
    .B1(u5_mul_69_18_n_327),
    .B2(u5_mul_69_18_n_420),
    .Y(u5_mul_69_18_n_706));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28170 (.A1(u5_mul_69_18_n_559),
    .A2(u5_mul_69_18_n_626),
    .B1(u5_mul_69_18_n_312),
    .B2(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_705));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28171 (.A1(u5_mul_69_18_n_350),
    .A2(u5_mul_69_18_n_637),
    .B1(u5_mul_69_18_n_234),
    .B2(u5_mul_69_18_n_421),
    .Y(u5_mul_69_18_n_703));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28172 (.A1(u5_mul_69_18_n_638),
    .A2(u5_mul_69_18_n_319),
    .B1(u5_mul_69_18_n_10),
    .B2(u5_mul_69_18_n_317),
    .Y(u5_mul_69_18_n_700));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28173 (.A1(u5_mul_69_18_n_410),
    .A2(u5_mul_69_18_n_642),
    .B1(u5_mul_69_18_n_394),
    .B2(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_699));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28174 (.A1(u5_mul_69_18_n_502),
    .A2(u5_mul_69_18_n_627),
    .B1(u5_mul_69_18_n_294),
    .B2(u5_mul_69_18_n_429),
    .Y(u5_mul_69_18_n_698));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28175 (.A1(u5_mul_69_18_n_341),
    .A2(u5_mul_69_18_n_630),
    .B1(u5_mul_69_18_n_334),
    .B2(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_696));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28176 (.A1(u5_mul_69_18_n_624),
    .A2(u5_mul_69_18_n_511),
    .B1(u5_mul_69_18_n_6),
    .B2(u5_mul_69_18_n_569),
    .Y(u5_mul_69_18_n_694));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28177 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_115),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_256),
    .Y(u5_mul_69_18_n_690));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28178 (.A(u5_mul_69_18_n_79),
    .B(u5_mul_69_18_n_620),
    .Y(u5_mul_69_18_n_689));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28179 (.A(u5_mul_69_18_n_82),
    .B(u5_mul_69_18_n_616),
    .Y(u5_mul_69_18_n_688));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28180 (.A(u5_mul_69_18_n_123),
    .B(u5_mul_69_18_n_614),
    .Y(u5_mul_69_18_n_687));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28181 (.A(u5_mul_69_18_n_92),
    .B(u5_mul_69_18_n_611),
    .Y(u5_mul_69_18_n_686));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28182 (.A(u5_mul_69_18_n_141),
    .B(u5_mul_69_18_n_615),
    .Y(u5_mul_69_18_n_685));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28183 (.A(u5_mul_69_18_n_139),
    .B(u5_mul_69_18_n_610),
    .Y(u5_mul_69_18_n_684));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28184 (.A(u5_mul_69_18_n_74),
    .B(u5_mul_69_18_n_618),
    .Y(u5_mul_69_18_n_683));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28185 (.A(u5_mul_69_18_n_134),
    .B(u5_mul_69_18_n_612),
    .Y(u5_mul_69_18_n_682));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28186 (.A(u5_mul_69_18_n_87),
    .B(u5_mul_69_18_n_619),
    .Y(u5_mul_69_18_n_681));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28187 (.A(u5_mul_69_18_n_129),
    .B(u5_mul_69_18_n_613),
    .Y(u5_mul_69_18_n_680));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28188 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_253),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_265),
    .Y(u5_mul_69_18_n_679));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28189 (.A(u5_mul_69_18_n_34),
    .B(u5_mul_69_18_n_617),
    .Y(u5_mul_69_18_n_678));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28190 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_262),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_253),
    .Y(u5_mul_69_18_n_677));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28191 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_259),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_266),
    .Y(u5_mul_69_18_n_676));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28192 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_265),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_259),
    .Y(u5_mul_69_18_n_675));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28193 (.A1(u5_mul_69_18_n_69),
    .A2(u5_mul_69_18_n_247),
    .B1(u5_mul_69_18_n_53),
    .B2(u5_mul_69_18_n_68),
    .Y(u5_mul_69_18_n_674));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28194 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_256),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_261),
    .Y(u5_mul_69_18_n_673));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28195 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_255),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_262),
    .Y(u5_mul_69_18_n_672));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28196 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_261),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_270),
    .Y(u5_mul_69_18_n_671));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28197 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_268),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_260),
    .Y(u5_mul_69_18_n_670));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28198 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_254),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_267),
    .Y(u5_mul_69_18_n_669));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28199 (.A1(u5_mul_69_18_n_69),
    .A2(u5_mul_69_18_n_264),
    .B1(u5_mul_69_18_n_68),
    .B2(u5_mul_69_18_n_251),
    .Y(u5_mul_69_18_n_668));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28200 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_269),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_245),
    .Y(u5_mul_69_18_n_667));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28201 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_250),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_258),
    .Y(u5_mul_69_18_n_666));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28202 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_263),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_248),
    .Y(u5_mul_69_18_n_665));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28203 (.A1(u5_mul_69_18_n_69),
    .A2(u5_mul_69_18_n_257),
    .B1(u5_mul_69_18_n_68),
    .B2(u5_mul_69_18_n_264),
    .Y(u5_mul_69_18_n_664));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28204 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_248),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_254),
    .Y(u5_mul_69_18_n_663));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28205 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_260),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_269),
    .Y(u5_mul_69_18_n_662));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g28206 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_266),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_263),
    .Y(u5_mul_69_18_n_661));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28207 (.A1(u5_mul_69_18_n_164),
    .A2(u5_mul_69_18_n_270),
    .B1(n_3303),
    .B2(u5_mul_69_18_n_255),
    .Y(u5_mul_69_18_n_660));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28208 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_267),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_268),
    .Y(u5_mul_69_18_n_659));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28209 (.A1(u5_mul_69_18_n_165),
    .A2(u5_mul_69_18_n_252),
    .B1(u5_mul_69_18_n_153),
    .B2(u5_mul_69_18_n_243),
    .Y(u5_mul_69_18_n_658));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28210 (.A1(u5_mul_69_18_n_69),
    .A2(u5_mul_69_18_n_246),
    .B1(u5_mul_69_18_n_68),
    .B2(u5_mul_69_18_n_249),
    .Y(u5_mul_69_18_n_657));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28211 (.A1(u5_mul_69_18_n_69),
    .A2(u5_mul_69_18_n_244),
    .B1(u5_mul_69_18_n_68),
    .B2(u5_mul_69_18_n_247),
    .Y(u5_mul_69_18_n_656));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28212 (.A(u5_mul_69_18_n_644),
    .Y(u5_mul_69_18_n_643));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28213 (.A(u5_mul_69_18_n_642),
    .Y(u5_mul_69_18_n_641));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28214 (.A(u5_mul_69_18_n_640),
    .Y(u5_mul_69_18_n_639));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28215 (.A(u5_mul_69_18_n_638),
    .Y(u5_mul_69_18_n_637));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28219 (.A(u5_mul_69_18_n_636),
    .Y(u5_mul_69_18_n_71));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28223 (.A(u5_mul_69_18_n_635),
    .Y(u5_mul_69_18_n_636));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28225 (.A(u5_mul_69_18_n_32),
    .Y(u5_mul_69_18_n_634));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28226 (.A(u5_mul_69_18_n_632),
    .Y(u5_mul_69_18_n_633));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28227 (.A(n_3302),
    .B(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_655));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28228 (.A(u5_mul_69_18_n_117),
    .B(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_654));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28229 (.A(n_3302),
    .B(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_653));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28230 (.A(u5_mul_69_18_n_118),
    .B(u5_mul_69_18_n_430),
    .Y(u5_mul_69_18_n_652));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28231 (.A(u5_mul_69_18_n_9),
    .B(n_3302),
    .Y(u5_mul_69_18_n_651));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28232 (.A(u5_mul_69_18_n_117),
    .B(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_650));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28233 (.A(u5_mul_69_18_n_118),
    .B(u5_mul_69_18_n_431),
    .Y(u5_mul_69_18_n_649));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28234 (.A(u5_mul_69_18_n_118),
    .B(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_648));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28235 (.A(u5_mul_69_18_n_118),
    .B(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_647));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28236 (.A(u5_mul_69_18_n_116),
    .B(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_646));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28237 (.A(u5_mul_69_18_n_116),
    .B(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_645));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28238 (.A1(n_14156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u5_mul_69_18_n_196),
    .C(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_644));
 A2O1A1Ixp33_ASAP7_75t_R u5_mul_69_18_g28239 (.A1(n_14160),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u5_mul_69_18_n_200),
    .C(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_642));
 A2O1A1Ixp33_ASAP7_75t_R u5_mul_69_18_g28240 (.A1(n_14148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B(u5_mul_69_18_n_193),
    .C(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_640));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28241 (.A1(n_14140),
    .A2(u5_mul_69_18_n_125),
    .B(u5_mul_69_18_n_199),
    .C(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_638));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28242 (.A1(n_14132),
    .A2(u5_mul_69_18_n_40),
    .B(u5_mul_69_18_n_202),
    .C(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_635));
 A2O1A1Ixp33_ASAP7_75t_R u5_mul_69_18_g28243 (.A1(u5_mul_69_18_n_146),
    .A2(n_14164),
    .B(u5_mul_69_18_n_203),
    .C(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_632));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28244 (.A(u5_mul_69_18_n_630),
    .Y(u5_mul_69_18_n_629));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28245 (.A(u5_mul_69_18_n_628),
    .Y(u5_mul_69_18_n_627));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28246 (.A(u5_mul_69_18_n_626),
    .Y(u5_mul_69_18_n_625));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28247 (.A(u5_mul_69_18_n_624),
    .Y(u5_mul_69_18_n_623));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28248 (.A(u5_mul_69_18_n_622),
    .Y(u5_mul_69_18_n_621));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28249 (.A(u5_mul_69_18_n_118),
    .B(n_14148),
    .C(u5_mul_69_18_n_123),
    .Y(u5_mul_69_18_n_620));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28250 (.A(u5_mul_69_18_n_118),
    .B(n_14136),
    .C(u5_mul_69_18_n_74),
    .Y(u5_mul_69_18_n_619));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28251 (.A(n_3302),
    .B(n_14132),
    .C(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_618));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28252 (.A(u5_mul_69_18_n_117),
    .B(n_14164),
    .C(u5_mul_69_18_n_143),
    .Y(u5_mul_69_18_n_617));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28253 (.A(n_3302),
    .B(n_14128),
    .C(u5_mul_69_18_n_94),
    .Y(u5_mul_69_18_n_616));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28254 (.A(u5_mul_69_18_n_117),
    .B(n_14160),
    .C(u5_mul_69_18_n_139),
    .Y(u5_mul_69_18_n_615));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28255 (.A(u5_mul_69_18_n_118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .C(u5_mul_69_18_n_129),
    .Y(u5_mul_69_18_n_614));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28256 (.A(u5_mul_69_18_n_118),
    .B(n_14140),
    .C(u5_mul_69_18_n_88),
    .Y(u5_mul_69_18_n_613));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28257 (.A(u5_mul_69_18_n_117),
    .B(n_14152),
    .C(u5_mul_69_18_n_79),
    .Y(u5_mul_69_18_n_612));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28258 (.A(u5_mul_69_18_n_99),
    .B(n_3302),
    .C(n_14178),
    .Y(u5_mul_69_18_n_611));
 MAJIxp5_ASAP7_75t_R u5_mul_69_18_g28259 (.A(u5_mul_69_18_n_117),
    .B(n_14156),
    .C(u5_mul_69_18_n_134),
    .Y(u5_mul_69_18_n_610));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28260 (.A1(u5_mul_69_18_n_153),
    .A2(u5_mul_69_18_n_165),
    .B(u5_mul_69_18_n_96),
    .Y(u5_mul_69_18_n_631));
 A2O1A1Ixp33_ASAP7_75t_R u5_mul_69_18_g28261 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u5_mul_69_18_n_197),
    .C(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_630));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28262 (.A1(n_14136),
    .A2(u5_mul_69_18_n_85),
    .B(u5_mul_69_18_n_198),
    .C(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_628));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28263 (.A1(n_14128),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B(u5_mul_69_18_n_201),
    .C(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_626));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28264 (.A1(n_14152),
    .A2(u5_mul_69_18_n_130),
    .B(u5_mul_69_18_n_195),
    .C(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_624));
 O2A1O1Ixp33_ASAP7_75t_R u5_mul_69_18_g28265 (.A1(n_14178),
    .A2(u5_mul_69_18_n_89),
    .B(u5_mul_69_18_n_194),
    .C(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_622));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28266 (.A(u5_mul_69_18_n_608),
    .Y(u5_mul_69_18_n_609));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28267 (.A(u5_mul_69_18_n_582),
    .Y(u5_mul_69_18_n_583));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28268 (.A(u5_mul_69_18_n_579),
    .Y(u5_mul_69_18_n_580));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28269 (.A(u5_mul_69_18_n_576),
    .Y(u5_mul_69_18_n_577));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28270 (.A(u5_mul_69_18_n_574),
    .Y(u5_mul_69_18_n_575));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28271 (.A(u5_mul_69_18_n_570),
    .Y(u5_mul_69_18_n_571));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28272 (.A(u5_mul_69_18_n_567),
    .Y(u5_mul_69_18_n_568));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28273 (.A(u5_mul_69_18_n_551),
    .Y(u5_mul_69_18_n_552));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28274 (.A(u5_mul_69_18_n_548),
    .Y(u5_mul_69_18_n_549));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28275 (.A(u5_mul_69_18_n_546),
    .Y(u5_mul_69_18_n_547));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28276 (.A(u5_mul_69_18_n_544),
    .Y(u5_mul_69_18_n_545));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28277 (.A(u5_mul_69_18_n_541),
    .Y(u5_mul_69_18_n_542));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28278 (.A(u5_mul_69_18_n_539),
    .Y(u5_mul_69_18_n_540));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28279 (.A(u5_mul_69_18_n_537),
    .Y(u5_mul_69_18_n_538));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28280 (.A(u5_mul_69_18_n_535),
    .Y(u5_mul_69_18_n_536));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28281 (.A(u5_mul_69_18_n_532),
    .Y(u5_mul_69_18_n_533));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28282 (.A(u5_mul_69_18_n_529),
    .Y(u5_mul_69_18_n_530));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28283 (.A(u5_mul_69_18_n_527),
    .Y(u5_mul_69_18_n_528));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28284 (.A(u5_mul_69_18_n_525),
    .Y(u5_mul_69_18_n_526));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28285 (.A(u5_mul_69_18_n_522),
    .Y(u5_mul_69_18_n_523));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28286 (.A(u5_mul_69_18_n_518),
    .Y(u5_mul_69_18_n_519));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28287 (.A(u5_mul_69_18_n_513),
    .Y(u5_mul_69_18_n_514));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28288 (.A(u5_mul_69_18_n_508),
    .Y(u5_mul_69_18_n_509));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28289 (.A(u5_mul_69_18_n_506),
    .Y(u5_mul_69_18_n_507));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28290 (.A(u5_mul_69_18_n_503),
    .Y(u5_mul_69_18_n_504));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28291 (.A(u5_mul_69_18_n_501),
    .Y(u5_mul_69_18_n_502));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28292 (.A(u5_mul_69_18_n_496),
    .Y(u5_mul_69_18_n_497));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28293 (.A(u5_mul_69_18_n_483),
    .Y(u5_mul_69_18_n_484));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28294 (.A(u5_mul_69_18_n_480),
    .Y(u5_mul_69_18_n_481));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28295 (.A(u5_mul_69_18_n_477),
    .Y(u5_mul_69_18_n_478));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28296 (.A(u5_mul_69_18_n_475),
    .Y(u5_mul_69_18_n_476));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28297 (.A(u5_mul_69_18_n_471),
    .Y(u5_mul_69_18_n_472));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28298 (.A(u5_mul_69_18_n_466),
    .Y(u5_mul_69_18_n_467));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28299 (.A(u5_mul_69_18_n_454),
    .Y(u5_mul_69_18_n_455));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28300 (.A(u5_mul_69_18_n_449),
    .Y(u5_mul_69_18_n_450));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28301 (.A(u5_mul_69_18_n_443),
    .Y(u5_mul_69_18_n_444));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28302 (.A(u5_mul_69_18_n_440),
    .Y(u5_mul_69_18_n_441));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28303 (.A(u5_mul_69_18_n_437),
    .Y(u5_mul_69_18_n_438));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28304 (.A(u5_mul_69_18_n_435),
    .Y(u5_mul_69_18_n_436));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28305 (.A(u5_mul_69_18_n_432),
    .Y(u5_mul_69_18_n_433));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28306 (.A(u5_mul_69_18_n_11),
    .Y(u5_mul_69_18_n_431));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28307 (.A(u5_mul_69_18_n_8),
    .Y(u5_mul_69_18_n_430));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28308 (.A(u5_mul_69_18_n_0),
    .Y(u5_mul_69_18_n_429));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28313 (.A(u5_mul_69_18_n_428),
    .Y(u5_mul_69_18_n_70));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28316 (.A(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_428));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28318 (.A(u5_mul_69_18_n_3),
    .Y(u5_mul_69_18_n_427));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28319 (.A(u5_mul_69_18_n_7),
    .Y(u5_mul_69_18_n_426));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28320 (.A(u5_mul_69_18_n_6),
    .Y(u5_mul_69_18_n_425));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28321 (.A(u5_mul_69_18_n_1),
    .Y(u5_mul_69_18_n_424));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28322 (.A(u5_mul_69_18_n_30),
    .Y(u5_mul_69_18_n_423));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28323 (.A(u5_mul_69_18_n_5),
    .Y(u5_mul_69_18_n_422));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28324 (.A(u5_mul_69_18_n_10),
    .Y(u5_mul_69_18_n_421));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28325 (.A(u5_mul_69_18_n_2),
    .Y(u5_mul_69_18_n_420));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28326 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_123),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_56),
    .Y(u5_mul_69_18_n_608));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28327 (.A1(n_13884),
    .A2(u5_mul_69_18_n_33),
    .B(u5_mul_69_18_n_192),
    .Y(u5_mul_69_18_n_607));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28328 (.A1(u5_mul_69_18_n_151),
    .A2(n_3336),
    .B(u5_mul_69_18_n_175),
    .Y(u5_mul_69_18_n_606));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28329 (.A1(u5_mul_69_18_n_152),
    .A2(n_3344),
    .B(u5_mul_69_18_n_185),
    .Y(u5_mul_69_18_n_605));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28330 (.A1(u5_mul_69_18_n_151),
    .A2(n_3353),
    .B(u5_mul_69_18_n_168),
    .Y(u5_mul_69_18_n_604));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28331 (.A1(u5_mul_69_18_n_152),
    .A2(n_3345),
    .B(u5_mul_69_18_n_213),
    .Y(u5_mul_69_18_n_603));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28332 (.A1(u5_mul_69_18_n_151),
    .A2(n_3341),
    .B(u5_mul_69_18_n_173),
    .Y(u5_mul_69_18_n_602));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28333 (.A1(u5_mul_69_18_n_152),
    .A2(n_3294),
    .B(u5_mul_69_18_n_218),
    .Y(u5_mul_69_18_n_601));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28334 (.A1(u5_mul_69_18_n_152),
    .A2(n_3305),
    .B(u5_mul_69_18_n_206),
    .Y(u5_mul_69_18_n_600));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28335 (.A1(u5_mul_69_18_n_152),
    .A2(n_3306),
    .B(u5_mul_69_18_n_190),
    .Y(u5_mul_69_18_n_599));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28336 (.A1(u5_mul_69_18_n_149),
    .A2(n_3297),
    .B(u5_mul_69_18_n_179),
    .Y(u5_mul_69_18_n_598));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28337 (.A1(u5_mul_69_18_n_149),
    .A2(n_3310),
    .B(u5_mul_69_18_n_170),
    .Y(u5_mul_69_18_n_597));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28338 (.A1(u5_mul_69_18_n_152),
    .A2(n_3355),
    .B(u5_mul_69_18_n_180),
    .Y(u5_mul_69_18_n_596));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28339 (.A1(u5_mul_69_18_n_149),
    .A2(n_3354),
    .B(u5_mul_69_18_n_210),
    .Y(u5_mul_69_18_n_595));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28340 (.A1(u5_mul_69_18_n_151),
    .A2(n_3337),
    .B(u5_mul_69_18_n_174),
    .Y(u5_mul_69_18_n_594));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28341 (.A1(u5_mul_69_18_n_149),
    .A2(n_3347),
    .B(u5_mul_69_18_n_186),
    .Y(u5_mul_69_18_n_593));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28342 (.A1(u5_mul_69_18_n_151),
    .A2(n_3350),
    .B(u5_mul_69_18_n_209),
    .Y(u5_mul_69_18_n_592));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28343 (.A1(u5_mul_69_18_n_151),
    .A2(n_3311),
    .B(u5_mul_69_18_n_211),
    .Y(u5_mul_69_18_n_591));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28344 (.A1(u5_mul_69_18_n_149),
    .A2(n_3351),
    .B(u5_mul_69_18_n_182),
    .Y(u5_mul_69_18_n_590));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28345 (.A1(u5_mul_69_18_n_149),
    .A2(n_3349),
    .B(u5_mul_69_18_n_204),
    .Y(u5_mul_69_18_n_589));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28346 (.A1(u5_mul_69_18_n_152),
    .A2(n_3299),
    .B(u5_mul_69_18_n_171),
    .Y(u5_mul_69_18_n_588));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28347 (.A1(u5_mul_69_18_n_151),
    .A2(n_3348),
    .B(u5_mul_69_18_n_216),
    .Y(u5_mul_69_18_n_587));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28348 (.A1(u5_mul_69_18_n_151),
    .A2(n_3358),
    .B(u5_mul_69_18_n_189),
    .Y(u5_mul_69_18_n_586));
 OAI21xp33_ASAP7_75t_R u5_mul_69_18_g28349 (.A1(u5_mul_69_18_n_149),
    .A2(n_3292),
    .B(u5_mul_69_18_n_167),
    .Y(u5_mul_69_18_n_585));
 OR2x2_ASAP7_75t_R u5_mul_69_18_g28350 (.A(u5_mul_69_18_n_52),
    .B(u5_n_2),
    .Y(u5_mul_69_18_n_584));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28351 (.A1(u5_mul_69_18_n_134),
    .A2(u5_mul_69_18_n_102),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_62),
    .Y(u5_mul_69_18_n_582));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28352 (.A1(n_3353),
    .A2(u5_mul_69_18_n_59),
    .B1(u5_mul_69_18_n_154),
    .B2(u5_mul_69_18_n_128),
    .Y(u5_mul_69_18_n_581));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28353 (.A1(n_3358),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_110),
    .B2(u5_mul_69_18_n_37),
    .Y(u5_mul_69_18_n_579));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28354 (.A1(u5_mul_69_18_n_159),
    .A2(u5_mul_69_18_n_142),
    .B1(n_3351),
    .B2(u5_mul_69_18_n_66),
    .Y(u5_mul_69_18_n_578));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28355 (.A1(n_3337),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_106),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_576));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28356 (.A1(n_3351),
    .A2(u5_mul_69_18_n_61),
    .B1(u5_mul_69_18_n_159),
    .B2(u5_mul_69_18_n_133),
    .Y(u5_mul_69_18_n_574));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28357 (.A1(n_3311),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_155),
    .B2(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_573));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28358 (.A1(u5_mul_69_18_n_48),
    .A2(n_3305),
    .B1(u5_mul_69_18_n_88),
    .B2(u5_mul_69_18_n_111),
    .Y(u5_mul_69_18_n_572));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28359 (.A1(u5_mul_69_18_n_91),
    .A2(u5_mul_69_18_n_162),
    .B1(u5_mul_69_18_n_50),
    .B2(n_3354),
    .Y(u5_mul_69_18_n_570));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28360 (.A1(u5_mul_69_18_n_156),
    .A2(u5_mul_69_18_n_133),
    .B1(n_3292),
    .B2(u5_mul_69_18_n_61),
    .Y(u5_mul_69_18_n_569));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28361 (.A1(u5_mul_69_18_n_55),
    .A2(n_3341),
    .B1(u5_mul_69_18_n_122),
    .B2(u5_mul_69_18_n_161),
    .Y(u5_mul_69_18_n_567));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28362 (.A1(n_3358),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_110),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_566));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28363 (.A1(n_3350),
    .A2(u5_mul_69_18_n_43),
    .B1(u5_mul_69_18_n_112),
    .B2(u5_mul_69_18_n_36),
    .Y(u5_mul_69_18_n_565));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28364 (.A1(u5_mul_69_18_n_112),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_564));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28365 (.A1(u5_mul_69_18_n_143),
    .A2(u5_mul_69_18_n_102),
    .B1(u5_mul_69_18_n_144),
    .B2(n_3345),
    .Y(u5_mul_69_18_n_563));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28366 (.A1(n_3354),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_73),
    .Y(u5_mul_69_18_n_562));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28367 (.A1(u5_mul_69_18_n_102),
    .A2(u5_mul_69_18_n_94),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_561));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28368 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_73),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_560));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28369 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_83),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_45),
    .Y(u5_mul_69_18_n_559));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28370 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_73),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_558));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28371 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_142),
    .B1(n_13884),
    .B2(u5_mul_69_18_n_66),
    .Y(u5_mul_69_18_n_557));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28372 (.A1(u5_mul_69_18_n_162),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3354),
    .B2(u5_mul_69_18_n_55),
    .Y(u5_mul_69_18_n_556));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28373 (.A1(u5_mul_69_18_n_64),
    .A2(n_3311),
    .B1(u5_mul_69_18_n_138),
    .B2(u5_mul_69_18_n_155),
    .Y(u5_mul_69_18_n_555));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28374 (.A1(u5_mul_69_18_n_57),
    .A2(n_3294),
    .B1(u5_mul_69_18_n_123),
    .B2(u5_mul_69_18_n_107),
    .Y(u5_mul_69_18_n_554));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28375 (.A1(u5_mul_69_18_n_100),
    .A2(u5_mul_69_18_n_94),
    .B1(n_3306),
    .B2(u5_mul_69_18_n_51),
    .Y(u5_mul_69_18_n_553));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28376 (.A1(n_3347),
    .A2(u5_mul_69_18_n_72),
    .B1(u5_mul_69_18_n_103),
    .B2(u5_mul_69_18_n_73),
    .Y(u5_mul_69_18_n_551));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28377 (.A1(u5_mul_69_18_n_107),
    .A2(u5_mul_69_18_n_74),
    .B1(n_3294),
    .B2(u5_mul_69_18_n_40),
    .Y(u5_mul_69_18_n_550));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28378 (.A1(u5_mul_69_18_n_67),
    .A2(n_3306),
    .B1(u5_mul_69_18_n_143),
    .B2(u5_mul_69_18_n_100),
    .Y(u5_mul_69_18_n_548));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28379 (.A1(u5_mul_69_18_n_110),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3358),
    .B2(u5_mul_69_18_n_56),
    .Y(u5_mul_69_18_n_546));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28380 (.A1(u5_mul_69_18_n_38),
    .A2(u5_mul_69_18_n_156),
    .B1(u5_mul_69_18_n_47),
    .B2(n_3292),
    .Y(u5_mul_69_18_n_544));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28381 (.A1(n_3299),
    .A2(u5_mul_69_18_n_60),
    .B1(u5_mul_69_18_n_105),
    .B2(u5_mul_69_18_n_129),
    .Y(u5_mul_69_18_n_543));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28382 (.A1(n_3305),
    .A2(u5_mul_69_18_n_46),
    .B1(u5_mul_69_18_n_111),
    .B2(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_541));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28383 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_56),
    .Y(u5_mul_69_18_n_539));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28384 (.A1(u5_mul_69_18_n_62),
    .A2(n_3294),
    .B1(u5_mul_69_18_n_134),
    .B2(u5_mul_69_18_n_107),
    .Y(u5_mul_69_18_n_537));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28385 (.A1(u5_mul_69_18_n_82),
    .A2(u5_mul_69_18_n_100),
    .B1(u5_mul_69_18_n_46),
    .B2(n_3306),
    .Y(u5_mul_69_18_n_535));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28386 (.A1(n_3344),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_37),
    .B2(u5_mul_69_18_n_113),
    .Y(u5_mul_69_18_n_534));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28387 (.A1(n_3345),
    .A2(u5_mul_69_18_n_57),
    .B1(u5_mul_69_18_n_123),
    .B2(u5_mul_69_18_n_102),
    .Y(u5_mul_69_18_n_532));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28388 (.A1(u5_mul_69_18_n_162),
    .A2(u5_mul_69_18_n_36),
    .B1(n_3354),
    .B2(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_531));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28389 (.A1(u5_mul_69_18_n_111),
    .A2(u5_mul_69_18_n_134),
    .B1(n_3305),
    .B2(u5_mul_69_18_n_132),
    .Y(u5_mul_69_18_n_529));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28390 (.A1(n_13883),
    .A2(u5_mul_69_18_n_55),
    .B1(u5_mul_69_18_n_108),
    .B2(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_527));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28391 (.A1(n_3348),
    .A2(u5_mul_69_18_n_47),
    .B1(u5_mul_69_18_n_157),
    .B2(u5_mul_69_18_n_38),
    .Y(u5_mul_69_18_n_525));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28392 (.A1(n_3306),
    .A2(u5_mul_69_18_n_57),
    .B1(u5_mul_69_18_n_123),
    .B2(u5_mul_69_18_n_100),
    .Y(u5_mul_69_18_n_524));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28393 (.A1(u5_mul_69_18_n_143),
    .A2(u5_mul_69_18_n_107),
    .B1(u5_mul_69_18_n_144),
    .B2(n_3294),
    .Y(u5_mul_69_18_n_522));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28394 (.A1(n_13883),
    .A2(u5_mul_69_18_n_50),
    .B1(u5_mul_69_18_n_108),
    .B2(u5_mul_69_18_n_91),
    .Y(u5_mul_69_18_n_521));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28395 (.A1(u5_mul_69_18_n_48),
    .A2(n_3299),
    .B1(u5_mul_69_18_n_88),
    .B2(u5_mul_69_18_n_105),
    .Y(u5_mul_69_18_n_520));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28396 (.A1(n_3351),
    .A2(u5_mul_69_18_n_42),
    .B1(u5_mul_69_18_n_159),
    .B2(u5_mul_69_18_n_78),
    .Y(u5_mul_69_18_n_518));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28397 (.A1(u5_mul_69_18_n_129),
    .A2(u5_mul_69_18_n_160),
    .B1(u5_mul_69_18_n_60),
    .B2(n_3355),
    .Y(u5_mul_69_18_n_517));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28398 (.A1(u5_mul_69_18_n_65),
    .A2(n_3355),
    .B1(u5_mul_69_18_n_139),
    .B2(u5_mul_69_18_n_160),
    .Y(u5_mul_69_18_n_516));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28399 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_133),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_61),
    .Y(u5_mul_69_18_n_515));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28400 (.A1(n_3294),
    .A2(u5_mul_69_18_n_46),
    .B1(u5_mul_69_18_n_107),
    .B2(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_513));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28401 (.A1(u5_mul_69_18_n_78),
    .A2(u5_mul_69_18_n_156),
    .B1(u5_mul_69_18_n_42),
    .B2(n_3292),
    .Y(u5_mul_69_18_n_512));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28402 (.A1(u5_mul_69_18_n_133),
    .A2(u5_mul_69_18_n_101),
    .B1(u5_mul_69_18_n_61),
    .B2(n_3297),
    .Y(u5_mul_69_18_n_511));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28403 (.A1(n_3341),
    .A2(u5_mul_69_18_n_58),
    .B1(u5_mul_69_18_n_161),
    .B2(u5_mul_69_18_n_128),
    .Y(u5_mul_69_18_n_510));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28404 (.A1(u5_mul_69_18_n_160),
    .A2(u5_mul_69_18_n_94),
    .B1(n_3355),
    .B2(u5_mul_69_18_n_51),
    .Y(u5_mul_69_18_n_508));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28405 (.A1(u5_mul_69_18_n_111),
    .A2(u5_mul_69_18_n_123),
    .B1(n_3305),
    .B2(u5_mul_69_18_n_57),
    .Y(u5_mul_69_18_n_506));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28406 (.A1(n_3347),
    .A2(u5_mul_69_18_n_61),
    .B1(u5_mul_69_18_n_103),
    .B2(u5_mul_69_18_n_133),
    .Y(u5_mul_69_18_n_505));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28407 (.A1(u5_mul_69_18_n_160),
    .A2(u5_mul_69_18_n_88),
    .B1(u5_mul_69_18_n_48),
    .B2(n_3355),
    .Y(u5_mul_69_18_n_503));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28408 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_38),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_501));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28409 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_127),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_500));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28410 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_127),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_499));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28411 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_111),
    .B1(n_3305),
    .B2(u5_mul_69_18_n_65),
    .Y(u5_mul_69_18_n_498));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28412 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_133),
    .B1(n_13883),
    .B2(u5_mul_69_18_n_61),
    .Y(u5_mul_69_18_n_496));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28413 (.A1(n_3348),
    .A2(u5_mul_69_18_n_64),
    .B1(u5_mul_69_18_n_157),
    .B2(u5_mul_69_18_n_138),
    .Y(u5_mul_69_18_n_495));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28414 (.A1(n_3297),
    .A2(u5_mul_69_18_n_50),
    .B1(u5_mul_69_18_n_101),
    .B2(u5_mul_69_18_n_91),
    .Y(u5_mul_69_18_n_494));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28415 (.A1(u5_mul_69_18_n_161),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3341),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_493));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28416 (.A1(u5_mul_69_18_n_121),
    .A2(u5_mul_69_18_n_159),
    .B1(u5_mul_69_18_n_55),
    .B2(n_3351),
    .Y(u5_mul_69_18_n_492));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28417 (.A1(n_3336),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_104),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_491));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28418 (.A1(u5_mul_69_18_n_133),
    .A2(u5_mul_69_18_n_109),
    .B1(u5_mul_69_18_n_61),
    .B2(n_3349),
    .Y(u5_mul_69_18_n_490));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28419 (.A1(u5_mul_69_18_n_134),
    .A2(u5_mul_69_18_n_160),
    .B1(u5_mul_69_18_n_62),
    .B2(n_3355),
    .Y(u5_mul_69_18_n_489));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28420 (.A1(u5_mul_69_18_n_62),
    .A2(n_3348),
    .B1(u5_mul_69_18_n_37),
    .B2(u5_mul_69_18_n_157),
    .Y(u5_mul_69_18_n_488));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28421 (.A1(n_3336),
    .A2(u5_mul_69_18_n_43),
    .B1(u5_mul_69_18_n_104),
    .B2(u5_mul_69_18_n_36),
    .Y(u5_mul_69_18_n_487));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28422 (.A1(u5_mul_69_18_n_60),
    .A2(n_3345),
    .B1(u5_mul_69_18_n_129),
    .B2(u5_mul_69_18_n_102),
    .Y(u5_mul_69_18_n_486));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28423 (.A1(n_3337),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_106),
    .B2(u5_mul_69_18_n_37),
    .Y(u5_mul_69_18_n_485));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28424 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_94),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_51),
    .Y(u5_mul_69_18_n_483));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28425 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_123),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_57),
    .Y(u5_mul_69_18_n_482));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28426 (.A1(n_3310),
    .A2(u5_mul_69_18_n_66),
    .B1(u5_mul_69_18_n_158),
    .B2(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_480));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28427 (.A1(n_3354),
    .A2(u5_mul_69_18_n_64),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_137),
    .Y(u5_mul_69_18_n_479));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28428 (.A1(u5_mul_69_18_n_110),
    .A2(u5_mul_69_18_n_128),
    .B1(n_3358),
    .B2(u5_mul_69_18_n_59),
    .Y(u5_mul_69_18_n_477));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28429 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_87),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_49),
    .Y(u5_mul_69_18_n_475));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28430 (.A1(n_3344),
    .A2(u5_mul_69_18_n_43),
    .B1(u5_mul_69_18_n_113),
    .B2(u5_mul_69_18_n_36),
    .Y(u5_mul_69_18_n_474));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28431 (.A1(u5_mul_69_18_n_138),
    .A2(u5_mul_69_18_n_112),
    .B1(u5_mul_69_18_n_64),
    .B2(n_3350),
    .Y(u5_mul_69_18_n_473));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28432 (.A1(n_3358),
    .A2(u5_mul_69_18_n_67),
    .B1(u5_mul_69_18_n_141),
    .B2(u5_mul_69_18_n_110),
    .Y(u5_mul_69_18_n_471));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28433 (.A1(u5_mul_69_18_n_50),
    .A2(n_3292),
    .B1(u5_mul_69_18_n_91),
    .B2(u5_mul_69_18_n_156),
    .Y(u5_mul_69_18_n_470));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28434 (.A1(u5_mul_69_18_n_112),
    .A2(u5_mul_69_18_n_123),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_57),
    .Y(u5_mul_69_18_n_469));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28435 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_55),
    .Y(u5_mul_69_18_n_468));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28436 (.A1(u5_mul_69_18_n_79),
    .A2(u5_mul_69_18_n_102),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_466));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28437 (.A1(u5_mul_69_18_n_112),
    .A2(u5_mul_69_18_n_87),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_49),
    .Y(u5_mul_69_18_n_465));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28438 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_36),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_464));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28439 (.A1(n_3305),
    .A2(u5_mul_69_18_n_51),
    .B1(u5_mul_69_18_n_111),
    .B2(u5_mul_69_18_n_94),
    .Y(u5_mul_69_18_n_463));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28440 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_74),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_40),
    .Y(u5_mul_69_18_n_462));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28441 (.A1(u5_mul_69_18_n_79),
    .A2(u5_mul_69_18_n_107),
    .B1(u5_mul_69_18_n_43),
    .B2(n_3294),
    .Y(u5_mul_69_18_n_461));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28442 (.A1(n_3348),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_157),
    .B2(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_460));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28443 (.A1(n_3337),
    .A2(u5_mul_69_18_n_43),
    .B1(u5_mul_69_18_n_106),
    .B2(u5_mul_69_18_n_36),
    .Y(u5_mul_69_18_n_459));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28444 (.A1(u5_mul_69_18_n_160),
    .A2(u5_mul_69_18_n_74),
    .B1(u5_mul_69_18_n_40),
    .B2(n_3355),
    .Y(u5_mul_69_18_n_458));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28445 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_37),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_62),
    .Y(u5_mul_69_18_n_457));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28446 (.A1(u5_mul_69_18_n_157),
    .A2(u5_mul_69_18_n_128),
    .B1(n_3348),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_456));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28447 (.A1(u5_mul_69_18_n_55),
    .A2(n_3348),
    .B1(u5_mul_69_18_n_122),
    .B2(u5_mul_69_18_n_157),
    .Y(u5_mul_69_18_n_454));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28448 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_50),
    .Y(u5_mul_69_18_n_453));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28449 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_100),
    .B1(u5_mul_69_18_n_65),
    .B2(n_3306),
    .Y(u5_mul_69_18_n_452));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28450 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_134),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_62),
    .Y(u5_mul_69_18_n_451));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28451 (.A1(u5_mul_69_18_n_144),
    .A2(n_3355),
    .B1(u5_mul_69_18_n_143),
    .B2(u5_mul_69_18_n_160),
    .Y(u5_mul_69_18_n_449));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28452 (.A1(n_3341),
    .A2(u5_mul_69_18_n_64),
    .B1(u5_mul_69_18_n_138),
    .B2(u5_mul_69_18_n_161),
    .Y(u5_mul_69_18_n_448));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28453 (.A1(u5_mul_69_18_n_100),
    .A2(u5_mul_69_18_n_74),
    .B1(n_3306),
    .B2(u5_mul_69_18_n_40),
    .Y(u5_mul_69_18_n_447));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28454 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_56),
    .Y(u5_mul_69_18_n_446));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28455 (.A1(u5_mul_69_18_n_73),
    .A2(u5_mul_69_18_n_156),
    .B1(u5_mul_69_18_n_72),
    .B2(n_3292),
    .Y(u5_mul_69_18_n_445));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28456 (.A1(u5_mul_69_18_n_43),
    .A2(n_3355),
    .B1(u5_mul_69_18_n_79),
    .B2(u5_mul_69_18_n_160),
    .Y(u5_mul_69_18_n_443));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28457 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_141),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_67),
    .Y(u5_mul_69_18_n_442));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28458 (.A1(u5_mul_69_18_n_138),
    .A2(u5_mul_69_18_n_110),
    .B1(u5_mul_69_18_n_63),
    .B2(n_3358),
    .Y(u5_mul_69_18_n_440));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28459 (.A1(u5_mul_69_18_n_113),
    .A2(u5_mul_69_18_n_129),
    .B1(n_3344),
    .B2(u5_mul_69_18_n_60),
    .Y(u5_mul_69_18_n_439));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28460 (.A1(u5_mul_69_18_n_101),
    .A2(u5_mul_69_18_n_38),
    .B1(n_3297),
    .B2(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_437));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28461 (.A1(u5_mul_69_18_n_160),
    .A2(u5_mul_69_18_n_84),
    .B1(u5_mul_69_18_n_46),
    .B2(n_3355),
    .Y(u5_mul_69_18_n_435));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28462 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_38),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_434));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28463 (.A1(u5_mul_69_18_n_87),
    .A2(u5_mul_69_18_n_161),
    .B1(u5_mul_69_18_n_49),
    .B2(n_3341),
    .Y(u5_mul_69_18_n_432));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28475 (.A(u5_mul_69_18_n_416),
    .Y(u5_mul_69_18_n_417));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28476 (.A(u5_mul_69_18_n_414),
    .Y(u5_mul_69_18_n_415));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28477 (.A(u5_mul_69_18_n_409),
    .Y(u5_mul_69_18_n_410));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28478 (.A(u5_mul_69_18_n_407),
    .Y(u5_mul_69_18_n_408));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28479 (.A(u5_mul_69_18_n_404),
    .Y(u5_mul_69_18_n_405));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28480 (.A(u5_mul_69_18_n_400),
    .Y(u5_mul_69_18_n_401));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28481 (.A(u5_mul_69_18_n_397),
    .Y(u5_mul_69_18_n_398));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28482 (.A(u5_mul_69_18_n_394),
    .Y(u5_mul_69_18_n_395));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28483 (.A(u5_mul_69_18_n_392),
    .Y(u5_mul_69_18_n_393));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28484 (.A(u5_mul_69_18_n_390),
    .Y(u5_mul_69_18_n_391));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28485 (.A(u5_mul_69_18_n_388),
    .Y(u5_mul_69_18_n_389));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28486 (.A(u5_mul_69_18_n_382),
    .Y(u5_mul_69_18_n_383));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28487 (.A(u5_mul_69_18_n_380),
    .Y(u5_mul_69_18_n_381));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28488 (.A(u5_mul_69_18_n_378),
    .Y(u5_mul_69_18_n_379));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28489 (.A(u5_mul_69_18_n_376),
    .Y(u5_mul_69_18_n_377));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28490 (.A(u5_mul_69_18_n_372),
    .Y(u5_mul_69_18_n_373));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28491 (.A(u5_mul_69_18_n_368),
    .Y(u5_mul_69_18_n_369));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28492 (.A(u5_mul_69_18_n_366),
    .Y(u5_mul_69_18_n_367));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28493 (.A(u5_mul_69_18_n_363),
    .Y(u5_mul_69_18_n_364));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28494 (.A(u5_mul_69_18_n_356),
    .Y(u5_mul_69_18_n_357));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28495 (.A(u5_mul_69_18_n_354),
    .Y(u5_mul_69_18_n_355));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28496 (.A(u5_mul_69_18_n_349),
    .Y(u5_mul_69_18_n_350));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28497 (.A(u5_mul_69_18_n_344),
    .Y(u5_mul_69_18_n_345));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28498 (.A(u5_mul_69_18_n_341),
    .Y(u5_mul_69_18_n_342));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28499 (.A(u5_mul_69_18_n_338),
    .Y(u5_mul_69_18_n_339));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28500 (.A(u5_mul_69_18_n_335),
    .Y(u5_mul_69_18_n_336));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28501 (.A(u5_mul_69_18_n_331),
    .Y(u5_mul_69_18_n_332));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28502 (.A(u5_mul_69_18_n_329),
    .Y(u5_mul_69_18_n_330));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28503 (.A(u5_mul_69_18_n_327),
    .Y(u5_mul_69_18_n_328));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28504 (.A(u5_mul_69_18_n_325),
    .Y(u5_mul_69_18_n_326));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28505 (.A(u5_mul_69_18_n_321),
    .Y(u5_mul_69_18_n_322));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28506 (.A(u5_mul_69_18_n_313),
    .Y(u5_mul_69_18_n_314));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28507 (.A(u5_mul_69_18_n_311),
    .Y(u5_mul_69_18_n_312));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28509 (.A(u5_mul_69_18_n_307),
    .Y(u5_mul_69_18_n_308));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28510 (.A(u5_mul_69_18_n_304),
    .Y(u5_mul_69_18_n_305));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28511 (.A(u5_mul_69_18_n_300),
    .Y(u5_mul_69_18_n_301));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28512 (.A(u5_mul_69_18_n_295),
    .Y(u5_mul_69_18_n_296));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28513 (.A(u5_mul_69_18_n_293),
    .Y(u5_mul_69_18_n_294));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28514 (.A(u5_mul_69_18_n_289),
    .Y(u5_mul_69_18_n_290));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28516 (.A(u5_mul_69_18_n_285),
    .Y(u5_mul_69_18_n_286));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28517 (.A(u5_mul_69_18_n_282),
    .Y(u5_mul_69_18_n_283));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28518 (.A(u5_mul_69_18_n_279),
    .Y(u5_mul_69_18_n_280));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28519 (.A(u5_mul_69_18_n_275),
    .Y(u5_mul_69_18_n_276));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28520 (.A(u5_mul_69_18_n_272),
    .Y(u5_mul_69_18_n_273));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28521 (.A(u5_mul_69_18_n_257),
    .Y(u5_mul_69_18_n_258));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28522 (.A(u5_mul_69_18_n_251),
    .Y(u5_mul_69_18_n_252));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28523 (.A(u5_mul_69_18_n_249),
    .Y(u5_mul_69_18_n_250));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28524 (.A(u5_mul_69_18_n_245),
    .Y(u5_mul_69_18_n_246));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28525 (.A(u5_mul_69_18_n_243),
    .Y(u5_mul_69_18_n_244));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28526 (.A(u5_mul_69_18_n_238),
    .Y(u5_mul_69_18_n_239));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28527 (.A(u5_mul_69_18_n_232),
    .Y(u5_mul_69_18_n_233));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28528 (.A1(u5_mul_69_18_n_65),
    .A2(u5_mul_69_18_n_117),
    .B1(u5_mul_69_18_n_139),
    .B2(u5_mul_69_18_n_116),
    .Y(u5_mul_69_18_n_229));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28529 (.A1(u5_mul_69_18_n_144),
    .A2(u5_mul_69_18_n_117),
    .B1(u5_mul_69_18_n_143),
    .B2(u5_mul_69_18_n_116),
    .Y(u5_mul_69_18_n_228));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28530 (.A1(u5_mul_69_18_n_84),
    .A2(u5_mul_69_18_n_115),
    .B1(u5_mul_69_18_n_46),
    .B2(n_3302),
    .Y(u5_mul_69_18_n_227));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28531 (.A1(u5_mul_69_18_n_43),
    .A2(u5_mul_69_18_n_117),
    .B1(u5_mul_69_18_n_79),
    .B2(u5_mul_69_18_n_54),
    .Y(u5_mul_69_18_n_226));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28532 (.A1(u5_mul_69_18_n_74),
    .A2(u5_mul_69_18_n_54),
    .B1(u5_mul_69_18_n_40),
    .B2(n_3302),
    .Y(u5_mul_69_18_n_225));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28534 (.A1(u5_mul_69_18_n_88),
    .A2(u5_mul_69_18_n_54),
    .B1(u5_mul_69_18_n_48),
    .B2(u5_mul_69_18_n_118),
    .Y(u5_mul_69_18_n_223));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28535 (.A1(u5_mul_69_18_n_54),
    .A2(u5_mul_69_18_n_129),
    .B1(u5_mul_69_18_n_117),
    .B2(u5_mul_69_18_n_60),
    .Y(u5_mul_69_18_n_222));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28536 (.A1(n_3302),
    .A2(u5_mul_69_18_n_93),
    .B1(u5_mul_69_18_n_92),
    .B2(u5_mul_69_18_n_115),
    .Y(u5_mul_69_18_n_221));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28537 (.A1(u5_mul_69_18_n_134),
    .A2(u5_mul_69_18_n_116),
    .B1(u5_mul_69_18_n_62),
    .B2(u5_mul_69_18_n_117),
    .Y(u5_mul_69_18_n_220));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28538 (.A1(u5_mul_69_18_n_57),
    .A2(u5_mul_69_18_n_117),
    .B1(u5_mul_69_18_n_123),
    .B2(u5_mul_69_18_n_54),
    .Y(u5_mul_69_18_n_219));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28539 (.A1(n_3350),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_37),
    .B2(u5_mul_69_18_n_112),
    .Y(u5_mul_69_18_n_419));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28540 (.A1(u5_mul_69_18_n_56),
    .A2(n_3344),
    .B1(u5_mul_69_18_n_122),
    .B2(u5_mul_69_18_n_113),
    .Y(u5_mul_69_18_n_418));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28541 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_79),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_416));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28542 (.A1(u5_mul_69_18_n_49),
    .A2(n_3294),
    .B1(u5_mul_69_18_n_88),
    .B2(u5_mul_69_18_n_107),
    .Y(u5_mul_69_18_n_414));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28543 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_413));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28544 (.A1(u5_mul_69_18_n_64),
    .A2(n_3353),
    .B1(u5_mul_69_18_n_138),
    .B2(u5_mul_69_18_n_154),
    .Y(u5_mul_69_18_n_412));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28545 (.A1(n_3305),
    .A2(u5_mul_69_18_n_77),
    .B1(u5_mul_69_18_n_79),
    .B2(u5_mul_69_18_n_111),
    .Y(u5_mul_69_18_n_411));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28546 (.A1(u5_mul_69_18_n_142),
    .A2(u5_mul_69_18_n_101),
    .B1(u5_mul_69_18_n_66),
    .B2(n_3297),
    .Y(u5_mul_69_18_n_409));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28547 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_137),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_63),
    .Y(u5_mul_69_18_n_407));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28548 (.A1(n_3354),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_406));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28549 (.A1(u5_mul_69_18_n_45),
    .A2(n_3351),
    .B1(u5_mul_69_18_n_83),
    .B2(u5_mul_69_18_n_159),
    .Y(u5_mul_69_18_n_404));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28550 (.A1(u5_mul_69_18_n_101),
    .A2(u5_mul_69_18_n_78),
    .B1(n_3297),
    .B2(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_403));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28551 (.A1(u5_mul_69_18_n_37),
    .A2(u5_mul_69_18_n_161),
    .B1(u5_mul_69_18_n_62),
    .B2(n_3341),
    .Y(u5_mul_69_18_n_402));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28552 (.A1(u5_mul_69_18_n_143),
    .A2(u5_mul_69_18_n_105),
    .B1(u5_mul_69_18_n_67),
    .B2(n_3299),
    .Y(u5_mul_69_18_n_400));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28553 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_87),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_49),
    .Y(u5_mul_69_18_n_399));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28554 (.A1(u5_mul_69_18_n_63),
    .A2(n_3347),
    .B1(u5_mul_69_18_n_137),
    .B2(u5_mul_69_18_n_103),
    .Y(u5_mul_69_18_n_397));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28555 (.A1(n_3345),
    .A2(u5_mul_69_18_n_46),
    .B1(u5_mul_69_18_n_102),
    .B2(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_396));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28556 (.A1(n_3292),
    .A2(u5_mul_69_18_n_66),
    .B1(u5_mul_69_18_n_156),
    .B2(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_394));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28557 (.A1(n_3341),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_161),
    .B2(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_392));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28558 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_82),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_45),
    .Y(u5_mul_69_18_n_390));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28559 (.A1(u5_mul_69_18_n_79),
    .A2(u5_mul_69_18_n_100),
    .B1(u5_mul_69_18_n_43),
    .B2(n_3306),
    .Y(u5_mul_69_18_n_388));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28560 (.A1(u5_mul_69_18_n_159),
    .A2(u5_mul_69_18_n_137),
    .B1(n_3351),
    .B2(u5_mul_69_18_n_63),
    .Y(u5_mul_69_18_n_387));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28561 (.A1(u5_mul_69_18_n_159),
    .A2(u5_mul_69_18_n_73),
    .B1(n_3351),
    .B2(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_386));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28562 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_36),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_385));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28563 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_129),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_59),
    .Y(u5_mul_69_18_n_384));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28564 (.A1(n_3353),
    .A2(u5_mul_69_18_n_45),
    .B1(u5_mul_69_18_n_154),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_382));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28565 (.A1(n_3344),
    .A2(u5_mul_69_18_n_49),
    .B1(u5_mul_69_18_n_113),
    .B2(u5_mul_69_18_n_87),
    .Y(u5_mul_69_18_n_380));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28566 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_38),
    .B1(n_13883),
    .B2(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_378));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28567 (.A1(n_3292),
    .A2(u5_mul_69_18_n_45),
    .B1(u5_mul_69_18_n_156),
    .B2(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_376));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28568 (.A1(n_3348),
    .A2(u5_mul_69_18_n_50),
    .B1(u5_mul_69_18_n_157),
    .B2(u5_mul_69_18_n_92),
    .Y(u5_mul_69_18_n_375));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28569 (.A1(u5_mul_69_18_n_138),
    .A2(u5_mul_69_18_n_106),
    .B1(u5_mul_69_18_n_63),
    .B2(n_3337),
    .Y(u5_mul_69_18_n_374));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28570 (.A1(u5_mul_69_18_n_78),
    .A2(u5_mul_69_18_n_158),
    .B1(u5_mul_69_18_n_42),
    .B2(n_3310),
    .Y(u5_mul_69_18_n_372));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28571 (.A1(n_3354),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_133),
    .Y(u5_mul_69_18_n_371));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28572 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_137),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_63),
    .Y(u5_mul_69_18_n_370));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28573 (.A1(n_3344),
    .A2(u5_mul_69_18_n_51),
    .B1(u5_mul_69_18_n_113),
    .B2(u5_mul_69_18_n_94),
    .Y(u5_mul_69_18_n_368));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28574 (.A1(u5_mul_69_18_n_137),
    .A2(u5_mul_69_18_n_108),
    .B1(u5_mul_69_18_n_63),
    .B2(n_13883),
    .Y(u5_mul_69_18_n_366));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28575 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_39),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_41),
    .Y(u5_mul_69_18_n_365));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28576 (.A1(u5_mul_69_18_n_55),
    .A2(n_3349),
    .B1(u5_mul_69_18_n_121),
    .B2(u5_mul_69_18_n_109),
    .Y(u5_mul_69_18_n_363));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28577 (.A1(u5_mul_69_18_n_43),
    .A2(n_3358),
    .B1(u5_mul_69_18_n_36),
    .B2(u5_mul_69_18_n_110),
    .Y(u5_mul_69_18_n_362));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28578 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_87),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_49),
    .Y(u5_mul_69_18_n_361));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28579 (.A1(u5_mul_69_18_n_162),
    .A2(u5_mul_69_18_n_128),
    .B1(n_3354),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_360));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28580 (.A1(u5_mul_69_18_n_141),
    .A2(u5_mul_69_18_n_112),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_67),
    .Y(u5_mul_69_18_n_359));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28581 (.A1(n_3311),
    .A2(u5_mul_69_18_n_67),
    .B1(u5_mul_69_18_n_155),
    .B2(u5_mul_69_18_n_141),
    .Y(u5_mul_69_18_n_358));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28582 (.A1(n_3305),
    .A2(u5_mul_69_18_n_67),
    .B1(u5_mul_69_18_n_143),
    .B2(u5_mul_69_18_n_111),
    .Y(u5_mul_69_18_n_356));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28583 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_354));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28584 (.A1(n_3341),
    .A2(u5_mul_69_18_n_66),
    .B1(u5_mul_69_18_n_141),
    .B2(u5_mul_69_18_n_161),
    .Y(u5_mul_69_18_n_353));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28585 (.A1(u5_mul_69_18_n_132),
    .A2(n_3306),
    .B1(u5_mul_69_18_n_134),
    .B2(u5_mul_69_18_n_100),
    .Y(u5_mul_69_18_n_352));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28586 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_83),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_45),
    .Y(u5_mul_69_18_n_351));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28587 (.A1(u5_mul_69_18_n_101),
    .A2(u5_mul_69_18_n_127),
    .B1(n_3297),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_349));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28588 (.A1(n_3353),
    .A2(u5_mul_69_18_n_67),
    .B1(u5_mul_69_18_n_141),
    .B2(u5_mul_69_18_n_154),
    .Y(u5_mul_69_18_n_348));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28589 (.A1(u5_mul_69_18_n_107),
    .A2(u5_mul_69_18_n_94),
    .B1(n_3294),
    .B2(u5_mul_69_18_n_51),
    .Y(u5_mul_69_18_n_347));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28590 (.A1(u5_mul_69_18_n_49),
    .A2(n_3358),
    .B1(u5_mul_69_18_n_87),
    .B2(u5_mul_69_18_n_110),
    .Y(u5_mul_69_18_n_346));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28591 (.A1(n_3349),
    .A2(u5_mul_69_18_n_66),
    .B1(u5_mul_69_18_n_109),
    .B2(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_344));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28592 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_78),
    .B1(n_13884),
    .B2(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_343));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28593 (.A1(n_3297),
    .A2(u5_mul_69_18_n_55),
    .B1(u5_mul_69_18_n_101),
    .B2(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_341));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28594 (.A1(u5_mul_69_18_n_110),
    .A2(u5_mul_69_18_n_39),
    .B1(n_3358),
    .B2(u5_mul_69_18_n_41),
    .Y(u5_mul_69_18_n_340));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28595 (.A1(u5_mul_69_18_n_37),
    .A2(u5_mul_69_18_n_155),
    .B1(u5_mul_69_18_n_62),
    .B2(n_3311),
    .Y(u5_mul_69_18_n_338));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28596 (.A1(n_3341),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_161),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_337));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28597 (.A1(n_3354),
    .A2(u5_mul_69_18_n_66),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_335));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28598 (.A1(n_3292),
    .A2(u5_mul_69_18_n_55),
    .B1(u5_mul_69_18_n_156),
    .B2(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_334));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28599 (.A1(u5_mul_69_18_n_101),
    .A2(u5_mul_69_18_n_73),
    .B1(n_3297),
    .B2(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_333));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28600 (.A1(u5_mul_69_18_n_91),
    .A2(u5_mul_69_18_n_103),
    .B1(u5_mul_69_18_n_50),
    .B2(n_3347),
    .Y(u5_mul_69_18_n_331));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28601 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_78),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_329));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28602 (.A1(n_3292),
    .A2(u5_mul_69_18_n_63),
    .B1(u5_mul_69_18_n_156),
    .B2(u5_mul_69_18_n_137),
    .Y(u5_mul_69_18_n_327));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28603 (.A1(u5_mul_69_18_n_39),
    .A2(u5_mul_69_18_n_104),
    .B1(u5_mul_69_18_n_41),
    .B2(n_3336),
    .Y(u5_mul_69_18_n_325));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28604 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_73),
    .B1(n_13884),
    .B2(u5_mul_69_18_n_72),
    .Y(u5_mul_69_18_n_324));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28605 (.A1(n_3297),
    .A2(u5_mul_69_18_n_63),
    .B1(u5_mul_69_18_n_101),
    .B2(u5_mul_69_18_n_137),
    .Y(u5_mul_69_18_n_323));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28606 (.A1(u5_mul_69_18_n_50),
    .A2(n_3310),
    .B1(u5_mul_69_18_n_91),
    .B2(u5_mul_69_18_n_158),
    .Y(u5_mul_69_18_n_321));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28607 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_105),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_65),
    .Y(u5_mul_69_18_n_320));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28608 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_127),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_319));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28609 (.A1(u5_mul_69_18_n_110),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3358),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_318));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28610 (.A1(u5_mul_69_18_n_159),
    .A2(u5_mul_69_18_n_127),
    .B1(n_3351),
    .B2(u5_mul_69_18_n_58),
    .Y(u5_mul_69_18_n_317));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28611 (.A1(u5_mul_69_18_n_157),
    .A2(u5_mul_69_18_n_36),
    .B1(n_3348),
    .B2(u5_mul_69_18_n_43),
    .Y(u5_mul_69_18_n_316));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28612 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_87),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_49),
    .Y(u5_mul_69_18_n_315));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28613 (.A1(u5_mul_69_18_n_102),
    .A2(u5_mul_69_18_n_88),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_48),
    .Y(u5_mul_69_18_n_313));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28614 (.A1(n_3297),
    .A2(u5_mul_69_18_n_45),
    .B1(u5_mul_69_18_n_101),
    .B2(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_311));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28615 (.A1(u5_mul_69_18_n_113),
    .A2(u5_mul_69_18_n_39),
    .B1(n_3344),
    .B2(u5_mul_69_18_n_41),
    .Y(u5_mul_69_18_n_310));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28616 (.A1(u5_mul_69_18_n_60),
    .A2(n_3306),
    .B1(u5_mul_69_18_n_129),
    .B2(u5_mul_69_18_n_100),
    .Y(u5_mul_69_18_n_309));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28617 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_107),
    .B1(u5_mul_69_18_n_65),
    .B2(n_3294),
    .Y(u5_mul_69_18_n_307));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28618 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_122),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_55),
    .Y(u5_mul_69_18_n_306));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28619 (.A1(n_3354),
    .A2(u5_mul_69_18_n_47),
    .B1(u5_mul_69_18_n_162),
    .B2(u5_mul_69_18_n_38),
    .Y(u5_mul_69_18_n_304));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28620 (.A1(u5_mul_69_18_n_66),
    .A2(n_3348),
    .B1(u5_mul_69_18_n_141),
    .B2(u5_mul_69_18_n_157),
    .Y(u5_mul_69_18_n_303));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28621 (.A1(n_3336),
    .A2(u5_mul_69_18_n_62),
    .B1(u5_mul_69_18_n_104),
    .B2(u5_mul_69_18_n_37),
    .Y(u5_mul_69_18_n_302));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28622 (.A1(n_3341),
    .A2(u5_mul_69_18_n_43),
    .B1(u5_mul_69_18_n_36),
    .B2(u5_mul_69_18_n_161),
    .Y(u5_mul_69_18_n_300));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28623 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_142),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_66),
    .Y(u5_mul_69_18_n_299));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28624 (.A1(n_3348),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_157),
    .B2(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_298));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28625 (.A1(u5_mul_69_18_n_57),
    .A2(n_3355),
    .B1(u5_mul_69_18_n_123),
    .B2(u5_mul_69_18_n_160),
    .Y(u5_mul_69_18_n_297));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28626 (.A1(n_3350),
    .A2(u5_mul_69_18_n_45),
    .B1(u5_mul_69_18_n_112),
    .B2(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_295));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28627 (.A1(u5_mul_69_18_n_38),
    .A2(u5_mul_69_18_n_159),
    .B1(u5_mul_69_18_n_47),
    .B2(n_3351),
    .Y(u5_mul_69_18_n_293));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28628 (.A1(n_13883),
    .A2(u5_mul_69_18_n_58),
    .B1(u5_mul_69_18_n_108),
    .B2(u5_mul_69_18_n_127),
    .Y(u5_mul_69_18_n_292));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28629 (.A1(u5_mul_69_18_n_100),
    .A2(u5_mul_69_18_n_88),
    .B1(n_3306),
    .B2(u5_mul_69_18_n_48),
    .Y(u5_mul_69_18_n_291));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28630 (.A1(n_3350),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_112),
    .B2(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_289));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28631 (.A1(u5_mul_69_18_n_111),
    .A2(u5_mul_69_18_n_39),
    .B1(n_3305),
    .B2(u5_mul_69_18_n_41),
    .Y(u5_mul_69_18_n_288));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28632 (.A1(u5_mul_69_18_n_158),
    .A2(u5_mul_69_18_n_38),
    .B1(n_3310),
    .B2(u5_mul_69_18_n_47),
    .Y(u5_mul_69_18_n_287));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28633 (.A1(u5_mul_69_18_n_60),
    .A2(n_3294),
    .B1(u5_mul_69_18_n_129),
    .B2(u5_mul_69_18_n_107),
    .Y(u5_mul_69_18_n_285));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28634 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_128),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_59),
    .Y(u5_mul_69_18_n_284));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28635 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_91),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_50),
    .Y(u5_mul_69_18_n_282));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28636 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_102),
    .B1(u5_mul_69_18_n_65),
    .B2(n_3345),
    .Y(u5_mul_69_18_n_281));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28637 (.A1(n_3311),
    .A2(u5_mul_69_18_n_59),
    .B1(u5_mul_69_18_n_155),
    .B2(u5_mul_69_18_n_128),
    .Y(u5_mul_69_18_n_279));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28638 (.A1(n_3351),
    .A2(u5_mul_69_18_n_50),
    .B1(u5_mul_69_18_n_159),
    .B2(u5_mul_69_18_n_91),
    .Y(u5_mul_69_18_n_278));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28639 (.A1(u5_mul_69_18_n_102),
    .A2(u5_mul_69_18_n_74),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_40),
    .Y(u5_mul_69_18_n_277));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28640 (.A1(u5_mul_69_18_n_121),
    .A2(u5_mul_69_18_n_158),
    .B1(u5_mul_69_18_n_55),
    .B2(n_3310),
    .Y(u5_mul_69_18_n_275));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28641 (.A1(u5_mul_69_18_n_108),
    .A2(u5_mul_69_18_n_83),
    .B1(fracta_mul[23]),
    .B2(u5_mul_69_18_n_45),
    .Y(u5_mul_69_18_n_274));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28642 (.A1(u5_mul_69_18_n_82),
    .A2(u5_mul_69_18_n_113),
    .B1(u5_mul_69_18_n_44),
    .B2(n_3344),
    .Y(u5_mul_69_18_n_272));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28643 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_92),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_93),
    .Y(u5_mul_69_18_n_271));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28644 (.A1(u5_mul_69_18_n_100),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3306),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_270));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28645 (.A1(u5_mul_69_18_n_162),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3354),
    .B2(u5_mul_69_18_n_53),
    .Y(u5_mul_69_18_n_269));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28646 (.A1(u5_mul_69_18_n_155),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3311),
    .B2(u5_mul_69_18_n_97),
    .Y(u5_mul_69_18_n_268));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28647 (.A1(u5_mul_69_18_n_154),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3353),
    .B2(u5_mul_69_18_n_97),
    .Y(u5_mul_69_18_n_267));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28648 (.A1(u5_mul_69_18_n_112),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_97),
    .Y(u5_mul_69_18_n_266));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28649 (.A1(u5_mul_69_18_n_113),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3344),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_265));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28650 (.A1(u5_mul_69_18_n_53),
    .A2(n_3349),
    .B1(u5_mul_69_18_n_96),
    .B2(u5_mul_69_18_n_109),
    .Y(u5_mul_69_18_n_264));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28651 (.A1(u5_mul_69_18_n_106),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_97),
    .Y(u5_mul_69_18_n_263));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28652 (.A1(u5_mul_69_18_n_105),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3299),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_262));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28653 (.A1(u5_mul_69_18_n_107),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3294),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_261));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28654 (.A1(u5_mul_69_18_n_157),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3348),
    .B2(u5_mul_69_18_n_97),
    .Y(u5_mul_69_18_n_260));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28655 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_259));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28656 (.A1(u5_mul_69_18_n_53),
    .A2(n_3310),
    .B1(u5_mul_69_18_n_96),
    .B2(u5_mul_69_18_n_158),
    .Y(u5_mul_69_18_n_257));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28657 (.A1(u5_mul_69_18_n_160),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3355),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_256));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28658 (.A1(u5_mul_69_18_n_102),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3345),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_255));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28659 (.A1(u5_mul_69_18_n_161),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3341),
    .B2(u5_mul_69_18_n_53),
    .Y(u5_mul_69_18_n_254));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28660 (.A1(u5_mul_69_18_n_111),
    .A2(u5_mul_69_18_n_99),
    .B1(n_3305),
    .B2(u5_mul_69_18_n_52),
    .Y(u5_mul_69_18_n_253));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28661 (.A1(u5_mul_69_18_n_53),
    .A2(n_3297),
    .B1(u5_mul_69_18_n_96),
    .B2(u5_mul_69_18_n_101),
    .Y(u5_mul_69_18_n_251));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28662 (.A1(u5_mul_69_18_n_53),
    .A2(n_3351),
    .B1(u5_mul_69_18_n_96),
    .B2(u5_mul_69_18_n_159),
    .Y(u5_mul_69_18_n_249));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28663 (.A1(u5_mul_69_18_n_110),
    .A2(u5_mul_69_18_n_98),
    .B1(n_3358),
    .B2(u5_mul_69_18_n_53),
    .Y(u5_mul_69_18_n_248));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28664 (.A1(n_13883),
    .A2(u5_mul_69_18_n_53),
    .B1(u5_mul_69_18_n_108),
    .B2(u5_mul_69_18_n_96),
    .Y(u5_mul_69_18_n_247));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28665 (.A1(u5_mul_69_18_n_103),
    .A2(u5_mul_69_18_n_96),
    .B1(n_3347),
    .B2(u5_mul_69_18_n_53),
    .Y(u5_mul_69_18_n_245));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28666 (.A1(u5_mul_69_18_n_156),
    .A2(u5_mul_69_18_n_96),
    .B1(n_3292),
    .B2(u5_mul_69_18_n_53),
    .Y(u5_mul_69_18_n_243));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28667 (.A1(u5_mul_69_18_n_139),
    .A2(u5_mul_69_18_n_113),
    .B1(n_3344),
    .B2(u5_mul_69_18_n_65),
    .Y(u5_mul_69_18_n_242));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28668 (.A1(u5_mul_69_18_n_104),
    .A2(u5_mul_69_18_n_139),
    .B1(n_3336),
    .B2(u5_mul_69_18_n_64),
    .Y(u5_mul_69_18_n_241));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28669 (.A1(u5_mul_69_18_n_141),
    .A2(u5_mul_69_18_n_106),
    .B1(n_3337),
    .B2(u5_mul_69_18_n_67),
    .Y(u5_mul_69_18_n_240));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28670 (.A1(u5_mul_69_18_n_109),
    .A2(u5_mul_69_18_n_78),
    .B1(n_3349),
    .B2(u5_mul_69_18_n_42),
    .Y(u5_mul_69_18_n_238));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28671 (.A1(n_3299),
    .A2(u5_mul_69_18_n_46),
    .B1(u5_mul_69_18_n_105),
    .B2(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_237));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28672 (.A1(u5_mul_69_18_n_112),
    .A2(u5_mul_69_18_n_128),
    .B1(n_3350),
    .B2(u5_mul_69_18_n_59),
    .Y(u5_mul_69_18_n_236));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28673 (.A1(n_3347),
    .A2(u5_mul_69_18_n_44),
    .B1(u5_mul_69_18_n_103),
    .B2(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_235));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28674 (.A1(u5_mul_69_18_n_58),
    .A2(n_3292),
    .B1(u5_mul_69_18_n_127),
    .B2(u5_mul_69_18_n_156),
    .Y(u5_mul_69_18_n_234));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28675 (.A1(n_3305),
    .A2(u5_mul_69_18_n_60),
    .B1(u5_mul_69_18_n_111),
    .B2(u5_mul_69_18_n_129),
    .Y(u5_mul_69_18_n_232));
 OAI22xp33_ASAP7_75t_R u5_mul_69_18_g28676 (.A1(u5_mul_69_18_n_143),
    .A2(u5_mul_69_18_n_113),
    .B1(u5_mul_69_18_n_144),
    .B2(n_3344),
    .Y(u5_mul_69_18_n_231));
 AOI22xp33_ASAP7_75t_R u5_mul_69_18_g28677 (.A1(n_3353),
    .A2(u5_mul_69_18_n_41),
    .B1(u5_mul_69_18_n_154),
    .B2(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_230));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28678 (.A(u5_mul_69_18_n_218),
    .Y(u5_mul_69_18_n_217));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28679 (.A(u5_mul_69_18_n_216),
    .Y(u5_mul_69_18_n_215));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28680 (.A(u5_mul_69_18_n_213),
    .Y(u5_mul_69_18_n_214));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28681 (.A(u5_mul_69_18_n_211),
    .Y(u5_mul_69_18_n_212));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28682 (.A(u5_mul_69_18_n_209),
    .Y(u5_mul_69_18_n_208));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28683 (.A(u5_mul_69_18_n_206),
    .Y(u5_mul_69_18_n_207));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28684 (.A(u5_mul_69_18_n_204),
    .Y(u5_mul_69_18_n_205));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28685 (.A(u5_mul_69_18_n_146),
    .B(n_14164),
    .Y(u5_mul_69_18_n_203));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28686 (.A(n_14132),
    .B(u5_mul_69_18_n_40),
    .Y(u5_mul_69_18_n_202));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28687 (.A(n_14128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .Y(u5_mul_69_18_n_201));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28688 (.A(n_14160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .Y(u5_mul_69_18_n_200));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28689 (.A(n_14140),
    .B(u5_mul_69_18_n_125),
    .Y(u5_mul_69_18_n_199));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28690 (.A(n_14136),
    .B(u5_mul_69_18_n_85),
    .Y(u5_mul_69_18_n_198));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .Y(u5_mul_69_18_n_197));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28692 (.A(n_14156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .Y(u5_mul_69_18_n_196));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28693 (.A(n_14152),
    .B(u5_mul_69_18_n_130),
    .Y(u5_mul_69_18_n_195));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28694 (.A(n_14178),
    .B(u5_mul_69_18_n_89),
    .Y(u5_mul_69_18_n_194));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28695 (.A(n_14148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(u5_mul_69_18_n_193));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28696 (.A(u5_mul_69_18_n_152),
    .B(n_3294),
    .Y(u5_mul_69_18_n_218));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28697 (.A(u5_mul_69_18_n_151),
    .B(n_3348),
    .Y(u5_mul_69_18_n_216));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28698 (.A(n_3345),
    .B(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_213));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28699 (.A(n_3311),
    .B(u5_mul_69_18_n_35),
    .Y(u5_mul_69_18_n_211));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28700 (.A(u5_mul_69_18_n_151),
    .B(n_3354),
    .Y(u5_mul_69_18_n_210));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28701 (.A(u5_mul_69_18_n_151),
    .B(n_3350),
    .Y(u5_mul_69_18_n_209));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28702 (.A(u5_mul_69_18_n_152),
    .B(n_3305),
    .Y(u5_mul_69_18_n_206));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28703 (.A(n_3349),
    .B(u5_mul_69_18_n_149),
    .Y(u5_mul_69_18_n_204));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28704 (.A(u5_mul_69_18_n_190),
    .Y(u5_mul_69_18_n_191));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28705 (.A(u5_mul_69_18_n_189),
    .Y(u5_mul_69_18_n_188));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28706 (.A(u5_mul_69_18_n_186),
    .Y(u5_mul_69_18_n_187));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28707 (.A(u5_mul_69_18_n_185),
    .Y(u5_mul_69_18_n_184));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28708 (.A(u5_mul_69_18_n_182),
    .Y(u5_mul_69_18_n_183));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28709 (.A(u5_mul_69_18_n_180),
    .Y(u5_mul_69_18_n_181));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28710 (.A(u5_mul_69_18_n_179),
    .Y(u5_mul_69_18_n_178));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28711 (.A(u5_mul_69_18_n_175),
    .Y(u5_mul_69_18_n_176));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28712 (.A(u5_mul_69_18_n_171),
    .Y(u5_mul_69_18_n_172));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28713 (.A(u5_mul_69_18_n_168),
    .Y(u5_mul_69_18_n_169));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28714 (.A(u5_mul_69_18_n_167),
    .Y(u5_mul_69_18_n_166));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28717 (.A(u5_mul_69_18_n_165),
    .Y(u5_mul_69_18_n_69));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28720 (.A(u5_mul_69_18_n_164),
    .Y(u5_mul_69_18_n_165));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28721 (.A(u5_mul_69_18_n_34),
    .B(u5_mul_69_18_n_117),
    .Y(u5_mul_69_18_n_163));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28723 (.A(u5_mul_69_18_n_149),
    .B(fracta_mul[23]),
    .Y(u5_mul_69_18_n_192));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28724 (.A(n_3306),
    .B(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_190));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28725 (.A(u5_mul_69_18_n_35),
    .B(n_3358),
    .Y(u5_mul_69_18_n_189));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28726 (.A(n_3347),
    .B(u5_mul_69_18_n_149),
    .Y(u5_mul_69_18_n_186));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28727 (.A(u5_mul_69_18_n_34),
    .B(n_3344),
    .Y(u5_mul_69_18_n_185));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28728 (.A(u5_mul_69_18_n_149),
    .B(n_3351),
    .Y(u5_mul_69_18_n_182));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28729 (.A(n_3355),
    .B(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_180));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28730 (.A(u5_mul_69_18_n_33),
    .B(n_3297),
    .Y(u5_mul_69_18_n_179));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28731 (.A(u5_mul_69_18_n_148),
    .B(u5_mul_69_18_n_116),
    .Y(u5_mul_69_18_n_177));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28732 (.A(n_3336),
    .B(u5_mul_69_18_n_35),
    .Y(u5_mul_69_18_n_175));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28733 (.A(u5_mul_69_18_n_151),
    .B(n_3337),
    .Y(u5_mul_69_18_n_174));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28734 (.A(u5_mul_69_18_n_151),
    .B(n_3341),
    .Y(u5_mul_69_18_n_173));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28735 (.A(u5_mul_69_18_n_152),
    .B(n_3299),
    .Y(u5_mul_69_18_n_171));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28736 (.A(u5_mul_69_18_n_149),
    .B(n_3310),
    .Y(u5_mul_69_18_n_170));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28737 (.A(u5_mul_69_18_n_151),
    .B(n_3353),
    .Y(u5_mul_69_18_n_168));
 NAND2xp33_ASAP7_75t_R u5_mul_69_18_g28738 (.A(u5_mul_69_18_n_149),
    .B(n_3292),
    .Y(u5_mul_69_18_n_167));
 NOR2xp33_ASAP7_75t_R u5_mul_69_18_g28739 (.A(n_3303),
    .B(u5_mul_69_18_n_95),
    .Y(u5_mul_69_18_n_164));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28747 (.A(n_3354),
    .Y(u5_mul_69_18_n_162));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28748 (.A(n_3341),
    .Y(u5_mul_69_18_n_161));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28749 (.A(n_3355),
    .Y(u5_mul_69_18_n_160));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28750 (.A(n_3351),
    .Y(u5_mul_69_18_n_159));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28751 (.A(n_3310),
    .Y(u5_mul_69_18_n_158));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28752 (.A(n_3348),
    .Y(u5_mul_69_18_n_157));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28753 (.A(n_3292),
    .Y(u5_mul_69_18_n_156));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28754 (.A(n_3311),
    .Y(u5_mul_69_18_n_155));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28755 (.A(n_3353),
    .Y(u5_mul_69_18_n_154));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28760 (.A(u5_mul_69_18_n_153),
    .Y(u5_mul_69_18_n_68));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28761 (.A(n_3303),
    .Y(u5_mul_69_18_n_153));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28763 (.A(u5_mul_69_18_n_149),
    .Y(u5_mul_69_18_n_150));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28764 (.A(u5_mul_69_18_n_151),
    .Y(u5_mul_69_18_n_149));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28765 (.A(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_151));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28766 (.A(u5_mul_69_18_n_152),
    .Y(u5_mul_69_18_n_148));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28767 (.A(fractb_mul[23]),
    .Y(u5_mul_69_18_n_152));
 INVxp67_ASAP7_75t_L u5_mul_69_18_g28768 (.A(fractb_mul[23]),
    .Y(u5_mul_69_18_n_146));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28771 (.A(u5_mul_69_18_n_143),
    .Y(u5_mul_69_18_n_144));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28783 (.A(u5_mul_69_18_n_141),
    .Y(u5_mul_69_18_n_142));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28784 (.A(u5_mul_69_18_n_142),
    .Y(u5_mul_69_18_n_66));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28786 (.A(u5_mul_69_18_n_141),
    .Y(u5_mul_69_18_n_67));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28792 (.A(u5_mul_69_18_n_143),
    .Y(u5_mul_69_18_n_141));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28813 (.A(u5_mul_69_18_n_137),
    .Y(u5_mul_69_18_n_63));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28815 (.A(u5_mul_69_18_n_138),
    .Y(u5_mul_69_18_n_137));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28822 (.A(u5_mul_69_18_n_138),
    .Y(u5_mul_69_18_n_64));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28823 (.A(u5_mul_69_18_n_139),
    .Y(u5_mul_69_18_n_138));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u5_mul_69_18_n_139));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28841 (.A(u5_mul_69_18_n_133),
    .Y(u5_mul_69_18_n_61));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28847 (.A(u5_mul_69_18_n_37),
    .Y(u5_mul_69_18_n_133));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28854 (.A(u5_mul_69_18_n_134),
    .Y(u5_mul_69_18_n_132));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28860 (.A(n_14154),
    .Y(u5_mul_69_18_n_134));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28862 (.A(n_14154),
    .Y(u5_mul_69_18_n_130));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28872 (.A(u5_mul_69_18_n_127),
    .Y(u5_mul_69_18_n_58));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28882 (.A(u5_mul_69_18_n_128),
    .Y(u5_mul_69_18_n_127));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28884 (.A(u5_mul_69_18_n_128),
    .Y(u5_mul_69_18_n_59));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28888 (.A(u5_mul_69_18_n_129),
    .Y(u5_mul_69_18_n_128));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28892 (.A(n_14142),
    .Y(u5_mul_69_18_n_129));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28894 (.A(n_14142),
    .Y(u5_mul_69_18_n_125));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28904 (.A(u5_mul_69_18_n_122),
    .Y(u5_mul_69_18_n_56));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28909 (.A(u5_mul_69_18_n_121),
    .Y(u5_mul_69_18_n_55));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28916 (.A(u5_mul_69_18_n_122),
    .Y(u5_mul_69_18_n_121));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28920 (.A(u5_mul_69_18_n_123),
    .Y(u5_mul_69_18_n_122));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28923 (.A(n_14146),
    .Y(u5_mul_69_18_n_123));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28928 (.A(u5_mul_69_18_n_117),
    .Y(u5_mul_69_18_n_116));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28934 (.A(u5_mul_69_18_n_118),
    .Y(u5_mul_69_18_n_117));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28936 (.A(u5_mul_69_18_n_118),
    .Y(u5_mul_69_18_n_54));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28939 (.A(n_3302),
    .Y(u5_mul_69_18_n_118));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28947 (.A(n_3344),
    .Y(u5_mul_69_18_n_113));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28948 (.A(n_3350),
    .Y(u5_mul_69_18_n_112));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28949 (.A(n_3305),
    .Y(u5_mul_69_18_n_111));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28950 (.A(n_3358),
    .Y(u5_mul_69_18_n_110));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28951 (.A(n_3349),
    .Y(u5_mul_69_18_n_109));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28952 (.A(n_13883),
    .Y(u5_mul_69_18_n_108));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28953 (.A(n_3294),
    .Y(u5_mul_69_18_n_107));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28954 (.A(n_3337),
    .Y(u5_mul_69_18_n_106));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28955 (.A(n_3299),
    .Y(u5_mul_69_18_n_105));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28956 (.A(n_3336),
    .Y(u5_mul_69_18_n_104));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28957 (.A(n_3347),
    .Y(u5_mul_69_18_n_103));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28958 (.A(n_3345),
    .Y(u5_mul_69_18_n_102));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28959 (.A(n_3297),
    .Y(u5_mul_69_18_n_101));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28960 (.A(n_3306),
    .Y(u5_mul_69_18_n_100));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28962 (.A(u5_mul_69_18_n_98),
    .Y(u5_mul_69_18_n_97));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28965 (.A(u5_mul_69_18_n_96),
    .Y(u5_mul_69_18_n_53));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28973 (.A(u5_mul_69_18_n_98),
    .Y(u5_mul_69_18_n_96));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28978 (.A(u5_mul_69_18_n_99),
    .Y(u5_mul_69_18_n_98));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g28989 (.A(n_14124),
    .Y(u5_mul_69_18_n_99));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28990 (.A(n_14124),
    .Y(u5_mul_69_18_n_95));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28993 (.A(u5_mul_69_18_n_94),
    .Y(u5_mul_69_18_n_51));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g28995 (.A(u5_mul_69_18_n_92),
    .Y(u5_mul_69_18_n_93));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29005 (.A(u5_mul_69_18_n_91),
    .Y(u5_mul_69_18_n_50));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29009 (.A(u5_mul_69_18_n_92),
    .Y(u5_mul_69_18_n_91));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29013 (.A(u5_mul_69_18_n_94),
    .Y(u5_mul_69_18_n_92));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29019 (.A(n_14126),
    .Y(u5_mul_69_18_n_94));
 INVx1_ASAP7_75t_R u5_mul_69_18_g29021 (.A(n_14126),
    .Y(u5_mul_69_18_n_89));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29044 (.A(u5_mul_69_18_n_87),
    .Y(u5_mul_69_18_n_49));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29045 (.A(u5_mul_69_18_n_88),
    .Y(u5_mul_69_18_n_87));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29050 (.A(u5_mul_69_18_n_88),
    .Y(u5_mul_69_18_n_48));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u5_mul_69_18_n_88));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u5_mul_69_18_n_85));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29063 (.A(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_83));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29068 (.A(u5_mul_69_18_n_83),
    .Y(u5_mul_69_18_n_45));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29070 (.A(u5_mul_69_18_n_82),
    .Y(u5_mul_69_18_n_44));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29074 (.A(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_82));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29078 (.A(u5_mul_69_18_n_84),
    .Y(u5_mul_69_18_n_46));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29082 (.A(n_14130),
    .Y(u5_mul_69_18_n_84));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29092 (.A(u5_mul_69_18_n_78),
    .Y(u5_mul_69_18_n_42));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29100 (.A(u5_mul_69_18_n_36),
    .Y(u5_mul_69_18_n_78));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29107 (.A(u5_mul_69_18_n_79),
    .Y(u5_mul_69_18_n_77));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29113 (.A(n_14150),
    .Y(u5_mul_69_18_n_79));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29123 (.A(u5_mul_69_18_n_73),
    .Y(u5_mul_69_18_n_72));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29131 (.A(u5_mul_69_18_n_39),
    .Y(u5_mul_69_18_n_73));
 INVxp33_ASAP7_75t_R u5_mul_69_18_g29140 (.A(u5_mul_69_18_n_74),
    .Y(u5_mul_69_18_n_40));
 HB1xp67_ASAP7_75t_R u5_mul_69_18_g29146 (.A(n_14134),
    .Y(u5_mul_69_18_n_74));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29438 (.A(n_14303),
    .B(u5_mul_69_18_n_1875),
    .Y(u5_mul_69_18_n_26));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29439 (.A(u5_mul_69_18_n_1849),
    .B(n_14306),
    .Y(u5_mul_69_18_n_25));
 OR2x2_ASAP7_75t_R u5_mul_69_18_g29440 (.A(u5_mul_69_18_n_1826),
    .B(n_14312),
    .Y(u5_mul_69_18_n_24));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29441 (.A(n_14316),
    .B(u5_mul_69_18_n_1794),
    .Y(u5_mul_69_18_n_23));
 OR2x2_ASAP7_75t_R u5_mul_69_18_g29442 (.A(u5_mul_69_18_n_1753),
    .B(n_14315),
    .Y(u5_mul_69_18_n_22));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29444 (.A(u5_mul_69_18_n_1737),
    .B(u5_mul_69_18_n_1708),
    .Y(u5_mul_69_18_n_20));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29445 (.A(u5_mul_69_18_n_1664),
    .B(n_14332),
    .Y(u5_mul_69_18_n_19));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29450 (.A(u5_mul_69_18_n_984),
    .B(n_14397),
    .Y(u5_mul_69_18_n_14));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g29451 (.A(u5_mul_69_18_n_833),
    .B(u5_mul_69_18_n_680),
    .Y(u5_mul_69_18_n_13));
 AO22x1_ASAP7_75t_R u5_mul_69_18_g29452 (.A1(u5_mul_69_18_n_288),
    .A2(u5_mul_69_18_n_635),
    .B1(u5_mul_69_18_n_310),
    .B2(u5_mul_69_18_n_9),
    .Y(u5_mul_69_18_n_12));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g29453 (.A(n_14148),
    .B(n_14146),
    .Y(u5_mul_69_18_n_11));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29454 (.A(n_14140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u5_mul_69_18_n_10));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29455 (.A(n_14132),
    .B(n_14130),
    .Y(u5_mul_69_18_n_9));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g29456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .B(n_14142),
    .Y(u5_mul_69_18_n_8));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29457 (.A(n_14124),
    .B(n_14178),
    .Y(u5_mul_69_18_n_7));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29458 (.A(n_14152),
    .B(n_14150),
    .Y(u5_mul_69_18_n_6));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g29459 (.A(n_14164),
    .B(u5_mul_69_18_n_143),
    .Y(u5_mul_69_18_n_5));
 AND2x2_ASAP7_75t_R u5_mul_69_18_g29460 (.A(n_3303),
    .B(n_3302),
    .Y(u5_n_2));
 XNOR2xp5_ASAP7_75t_R u5_mul_69_18_g29461 (.A(n_14160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u5_mul_69_18_n_3));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29462 (.A(n_14156),
    .B(n_14154),
    .Y(u5_mul_69_18_n_2));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29463 (.A(n_14128),
    .B(n_14126),
    .Y(u5_mul_69_18_n_1));
 XOR2xp5_ASAP7_75t_R u5_mul_69_18_g29464 (.A(n_14136),
    .B(n_14134),
    .Y(u5_mul_69_18_n_0));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[0]  (.CLK(clk),
    .D(n_742),
    .QN(u5_prod1[0]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[10]  (.CLK(clk),
    .D(n_14221),
    .QN(u5_prod1[10]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[11]  (.CLK(clk),
    .D(n_14196),
    .QN(u5_prod1[11]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[12]  (.CLK(clk),
    .D(n_14234),
    .QN(u5_prod1[12]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[13]  (.CLK(clk),
    .D(n_14257),
    .QN(u5_prod1[13]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[14]  (.CLK(clk),
    .D(n_14231),
    .QN(u5_prod1[14]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[15]  (.CLK(clk),
    .D(n_14243),
    .QN(u5_prod1[15]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[16]  (.CLK(clk),
    .D(n_14201),
    .QN(u5_prod1[16]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[17]  (.CLK(clk),
    .D(n_14226),
    .QN(u5_prod1[17]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[18]  (.CLK(clk),
    .D(n_14186),
    .QN(u5_prod1[18]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[19]  (.CLK(clk),
    .D(n_14267),
    .QN(u5_prod1[19]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[1]  (.CLK(clk),
    .D(n_14266),
    .QN(u5_prod1[1]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[20]  (.CLK(clk),
    .D(n_14222),
    .QN(u5_prod1[20]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[21]  (.CLK(clk),
    .D(n_14263),
    .QN(u5_prod1[21]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[22]  (.CLK(clk),
    .D(n_14241),
    .QN(u5_prod1[22]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[23]  (.CLK(clk),
    .D(n_14191),
    .QN(u5_prod1[23]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[24]  (.CLK(clk),
    .D(n_14230),
    .QN(u5_prod1[24]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[25]  (.CLK(clk),
    .D(n_14255),
    .QN(u5_prod1[25]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[26]  (.CLK(clk),
    .D(n_14233),
    .QN(u5_prod1[26]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[27]  (.CLK(clk),
    .D(n_14229),
    .QN(u5_prod1[27]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[28]  (.CLK(clk),
    .D(n_14252),
    .QN(u5_prod1[28]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[29]  (.CLK(clk),
    .D(n_14225),
    .QN(u5_prod1[29]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[2]  (.CLK(clk),
    .D(n_14262),
    .QN(u5_prod1[2]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[30]  (.CLK(clk),
    .D(n_14203),
    .QN(u5_prod1[30]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[31]  (.CLK(clk),
    .D(n_14193),
    .QN(u5_prod1[31]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[32]  (.CLK(clk),
    .D(n_14261),
    .QN(u5_prod1[32]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[33]  (.CLK(clk),
    .D(n_14236),
    .QN(u5_prod1[33]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[34]  (.CLK(clk),
    .D(n_14256),
    .QN(u5_prod1[34]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[35]  (.CLK(clk),
    .D(n_14250),
    .QN(u5_prod1[35]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[36]  (.CLK(clk),
    .D(n_14200),
    .QN(u5_prod1[36]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[37]  (.CLK(clk),
    .D(n_14244),
    .QN(u5_prod1[37]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[38]  (.CLK(clk),
    .D(n_14237),
    .QN(u5_prod1[38]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[39]  (.CLK(clk),
    .D(n_14245),
    .QN(u5_prod1[39]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[3]  (.CLK(clk),
    .D(n_14254),
    .QN(u5_prod1[3]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[40]  (.CLK(clk),
    .D(n_14249),
    .QN(u5_prod1[40]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[41]  (.CLK(clk),
    .D(n_14194),
    .QN(u5_prod1[41]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[42]  (.CLK(clk),
    .D(n_14183),
    .QN(u5_prod1[42]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[43]  (.CLK(clk),
    .D(n_14215),
    .QN(u5_prod1[43]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[44]  (.CLK(clk),
    .D(n_14220),
    .QN(u5_prod1[44]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[45]  (.CLK(clk),
    .D(n_14209),
    .QN(u5_prod1[45]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[46]  (.CLK(clk),
    .D(n_14212),
    .QN(u5_prod1[46]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[47]  (.CLK(clk),
    .D(n_14205),
    .QN(u5_prod1[47]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[4]  (.CLK(clk),
    .D(n_14235),
    .QN(u5_prod1[4]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[5]  (.CLK(clk),
    .D(n_14251),
    .QN(u5_prod1[5]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[6]  (.CLK(clk),
    .D(n_14210),
    .QN(u5_prod1[6]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[7]  (.CLK(clk),
    .D(n_14228),
    .QN(u5_prod1[7]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[8]  (.CLK(clk),
    .D(n_14218),
    .QN(u5_prod1[8]));
 DFFHQNx1_ASAP7_75t_R \u5_prod1_reg[9]  (.CLK(clk),
    .D(n_14247),
    .QN(u5_prod1[9]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[0]  (.CLK(clk),
    .D(n_945),
    .QN(prod[0]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[10]  (.CLK(clk),
    .D(n_902),
    .QN(prod[10]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[11]  (.CLK(clk),
    .D(n_935),
    .QN(prod[11]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[12]  (.CLK(clk),
    .D(n_933),
    .QN(prod[12]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[13]  (.CLK(clk),
    .D(n_882),
    .QN(prod[13]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[14]  (.CLK(clk),
    .D(n_883),
    .QN(prod[14]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[15]  (.CLK(clk),
    .D(n_952),
    .QN(prod[15]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[16]  (.CLK(clk),
    .D(n_903),
    .QN(prod[16]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[17]  (.CLK(clk),
    .D(n_973),
    .QN(prod[17]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[18]  (.CLK(clk),
    .D(n_887),
    .QN(prod[18]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[19]  (.CLK(clk),
    .D(n_890),
    .QN(prod[19]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[1]  (.CLK(clk),
    .D(n_922),
    .QN(prod[1]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[20]  (.CLK(clk),
    .D(n_970),
    .QN(prod[20]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[21]  (.CLK(clk),
    .D(n_915),
    .QN(prod[21]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[22]  (.CLK(clk),
    .D(n_954),
    .QN(prod[22]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[23]  (.CLK(clk),
    .D(n_980),
    .QN(prod[23]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[24]  (.CLK(clk),
    .D(n_932),
    .QN(prod[24]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[25]  (.CLK(clk),
    .D(n_889),
    .QN(prod[25]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[26]  (.CLK(clk),
    .D(n_911),
    .QN(prod[26]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[27]  (.CLK(clk),
    .D(n_934),
    .QN(prod[27]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[28]  (.CLK(clk),
    .D(n_927),
    .QN(prod[28]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[29]  (.CLK(clk),
    .D(n_919),
    .QN(prod[29]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[2]  (.CLK(clk),
    .D(n_966),
    .QN(prod[2]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[30]  (.CLK(clk),
    .D(n_914),
    .QN(prod[30]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[31]  (.CLK(clk),
    .D(n_930),
    .QN(prod[31]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[32]  (.CLK(clk),
    .D(n_892),
    .QN(prod[32]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[33]  (.CLK(clk),
    .D(n_941),
    .QN(prod[33]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[34]  (.CLK(clk),
    .D(n_885),
    .QN(prod[34]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[35]  (.CLK(clk),
    .D(n_965),
    .QN(prod[35]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[36]  (.CLK(clk),
    .D(n_913),
    .QN(prod[36]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[37]  (.CLK(clk),
    .D(n_979),
    .QN(prod[37]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[38]  (.CLK(clk),
    .D(n_918),
    .QN(prod[38]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[39]  (.CLK(clk),
    .D(n_983),
    .QN(prod[39]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[3]  (.CLK(clk),
    .D(n_896),
    .QN(prod[3]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[40]  (.CLK(clk),
    .D(n_943),
    .QN(prod[40]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[41]  (.CLK(clk),
    .D(n_906),
    .QN(prod[41]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[42]  (.CLK(clk),
    .D(n_912),
    .QN(prod[42]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[43]  (.CLK(clk),
    .D(n_931),
    .QN(prod[43]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[44]  (.CLK(clk),
    .D(n_968),
    .QN(prod[44]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[45]  (.CLK(clk),
    .D(n_937),
    .QN(prod[45]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[46]  (.CLK(clk),
    .D(n_938),
    .QN(prod[46]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[47]  (.CLK(clk),
    .D(n_957),
    .QN(prod[47]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[4]  (.CLK(clk),
    .D(n_949),
    .QN(prod[4]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[5]  (.CLK(clk),
    .D(n_978),
    .QN(prod[5]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[6]  (.CLK(clk),
    .D(n_888),
    .QN(prod[6]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[7]  (.CLK(clk),
    .D(n_928),
    .QN(prod[7]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[8]  (.CLK(clk),
    .D(n_916),
    .QN(prod[8]));
 DFFHQNx1_ASAP7_75t_R \u5_prod_reg[9]  (.CLK(clk),
    .D(n_894),
    .QN(prod[9]));
 DFFHQNx1_ASAP7_75t_L \u6_quo1_reg[0]  (.CLK(clk),
    .D(n_14080),
    .QN(n_14081));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[10]  (.CLK(clk),
    .D(n_14184),
    .QN(u6_quo1[10]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[11]  (.CLK(clk),
    .D(n_737),
    .QN(u6_quo1[11]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[12]  (.CLK(clk),
    .D(n_14204),
    .QN(u6_quo1[12]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[13]  (.CLK(clk),
    .D(n_740),
    .QN(u6_quo1[13]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[14]  (.CLK(clk),
    .D(n_14199),
    .QN(u6_quo1[14]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[15]  (.CLK(clk),
    .D(n_856),
    .QN(u6_quo1[15]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[16]  (.CLK(clk),
    .D(n_14190),
    .QN(u6_quo1[16]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[17]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9087),
    .QN(u6_quo1[17]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[18]  (.CLK(clk),
    .D(n_14248),
    .QN(u6_quo1[18]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[19]  (.CLK(clk),
    .D(n_851),
    .QN(u6_quo1[19]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[1]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13674),
    .QN(n_14085));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[20]  (.CLK(clk),
    .D(n_830),
    .QN(u6_quo1[20]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[21]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7921),
    .QN(u6_quo1[21]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[22]  (.CLK(clk),
    .D(n_14224),
    .QN(u6_quo1[22]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[23]  (.CLK(clk),
    .D(n_853),
    .QN(u6_quo1[23]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[24]  (.CLK(clk),
    .D(n_14219),
    .QN(u6_quo1[24]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[25]  (.CLK(clk),
    .D(n_769),
    .QN(u6_quo1[25]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[26]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1468),
    .QN(u6_quo1[26]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[27]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6181),
    .QN(u6_quo1[27]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[28]  (.CLK(clk),
    .D(n_849),
    .QN(u6_quo1[28]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[29]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5680),
    .QN(u6_quo1[29]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[2]  (.CLK(clk),
    .D(n_14192),
    .QN(u6_quo1[2]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[30]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5226),
    .QN(u6_quo1[30]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[31]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5177),
    .QN(u6_quo1[31]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[32]  (.CLK(clk),
    .D(n_848),
    .QN(u6_quo1[32]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[33]  (.CLK(clk),
    .D(n_817),
    .QN(u6_quo1[33]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[34]  (.CLK(clk),
    .D(n_14197),
    .QN(u6_quo1[34]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[35]  (.CLK(clk),
    .D(n_833),
    .QN(u6_quo1[35]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[36]  (.CLK(clk),
    .D(n_838),
    .QN(u6_quo1[36]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[37]  (.CLK(clk),
    .D(n_852),
    .QN(u6_quo1[37]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[38]  (.CLK(clk),
    .D(n_866),
    .QN(u6_quo1[38]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[39]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3572),
    .QN(u6_quo1[39]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[3]  (.CLK(clk),
    .D(n_839),
    .QN(u6_quo1[3]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[40]  (.CLK(clk),
    .D(n_810),
    .QN(u6_quo1[40]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[41]  (.CLK(clk),
    .D(n_809),
    .QN(u6_quo1[41]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[42]  (.CLK(clk),
    .D(n_771),
    .QN(u6_quo1[42]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[43]  (.CLK(clk),
    .D(n_847),
    .QN(u6_quo1[43]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[44]  (.CLK(clk),
    .D(n_761),
    .QN(u6_quo1[44]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[45]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3012),
    .QN(u6_quo1[45]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[46]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2927),
    .QN(u6_quo1[46]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[47]  (.CLK(clk),
    .D(n_870),
    .QN(u6_quo1[47]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[48]  (.CLK(clk),
    .D(n_763),
    .QN(u6_quo1[48]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[49]  (.CLK(clk),
    .D(n_14214),
    .QN(u6_quo1[49]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[4]  (.CLK(clk),
    .D(n_14264),
    .QN(u6_quo1[4]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[5]  (.CLK(clk),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12549),
    .QN(u6_quo1[5]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[6]  (.CLK(clk),
    .D(n_733),
    .QN(u6_quo1[6]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[7]  (.CLK(clk),
    .D(n_844),
    .QN(u6_quo1[7]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[8]  (.CLK(clk),
    .D(n_805),
    .QN(u6_quo1[8]));
 DFFHQNx1_ASAP7_75t_R \u6_quo1_reg[9]  (.CLK(clk),
    .D(n_854),
    .QN(u6_quo1[9]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[0]  (.CLK(clk),
    .D(n_14082),
    .QN(quo[0]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[10]  (.CLK(clk),
    .D(n_891),
    .QN(quo[10]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[11]  (.CLK(clk),
    .D(n_971),
    .QN(quo[11]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[12]  (.CLK(clk),
    .D(n_976),
    .QN(quo[12]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[13]  (.CLK(clk),
    .D(n_886),
    .QN(quo[13]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[14]  (.CLK(clk),
    .D(n_929),
    .QN(quo[14]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[15]  (.CLK(clk),
    .D(n_967),
    .QN(quo[15]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[16]  (.CLK(clk),
    .D(n_982),
    .QN(quo[16]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[17]  (.CLK(clk),
    .D(n_944),
    .QN(quo[17]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[18]  (.CLK(clk),
    .D(n_895),
    .QN(quo[18]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[19]  (.CLK(clk),
    .D(n_956),
    .QN(quo[19]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[1]  (.CLK(clk),
    .D(n_14086),
    .QN(quo[1]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[20]  (.CLK(clk),
    .D(n_909),
    .QN(quo[20]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[21]  (.CLK(clk),
    .D(n_897),
    .QN(quo[21]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[22]  (.CLK(clk),
    .D(n_953),
    .QN(quo[22]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[23]  (.CLK(clk),
    .D(n_908),
    .QN(quo[23]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[24]  (.CLK(clk),
    .D(n_984),
    .QN(quo[24]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[25]  (.CLK(clk),
    .D(n_964),
    .QN(quo[25]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[26]  (.CLK(clk),
    .D(n_901),
    .QN(quo[26]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[27]  (.CLK(clk),
    .D(n_962),
    .QN(quo[27]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[28]  (.CLK(clk),
    .D(n_904),
    .QN(quo[28]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[29]  (.CLK(clk),
    .D(n_961),
    .QN(quo[29]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[2]  (.CLK(clk),
    .D(n_898),
    .QN(quo[2]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[30]  (.CLK(clk),
    .D(n_963),
    .QN(quo[30]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[31]  (.CLK(clk),
    .D(n_921),
    .QN(quo[31]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[32]  (.CLK(clk),
    .D(n_905),
    .QN(quo[32]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[33]  (.CLK(clk),
    .D(n_975),
    .QN(quo[33]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[34]  (.CLK(clk),
    .D(n_958),
    .QN(quo[34]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[35]  (.CLK(clk),
    .D(n_955),
    .QN(quo[35]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[36]  (.CLK(clk),
    .D(n_985),
    .QN(quo[36]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[37]  (.CLK(clk),
    .D(n_910),
    .QN(quo[37]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[38]  (.CLK(clk),
    .D(n_917),
    .QN(quo[38]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[39]  (.CLK(clk),
    .D(n_920),
    .QN(quo[39]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[3]  (.CLK(clk),
    .D(n_977),
    .QN(quo[3]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[40]  (.CLK(clk),
    .D(n_974),
    .QN(quo[40]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[41]  (.CLK(clk),
    .D(n_936),
    .QN(quo[41]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[42]  (.CLK(clk),
    .D(n_981),
    .QN(quo[42]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[43]  (.CLK(clk),
    .D(n_923),
    .QN(quo[43]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[44]  (.CLK(clk),
    .D(n_950),
    .QN(quo[44]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[45]  (.CLK(clk),
    .D(n_907),
    .QN(quo[45]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[46]  (.CLK(clk),
    .D(n_946),
    .QN(quo[46]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[47]  (.CLK(clk),
    .D(n_969),
    .QN(quo[47]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[48]  (.CLK(clk),
    .D(n_959),
    .QN(quo[48]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[49]  (.CLK(clk),
    .D(n_947),
    .QN(quo[49]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[4]  (.CLK(clk),
    .D(n_951),
    .QN(quo[4]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[5]  (.CLK(clk),
    .D(n_960),
    .QN(quo[5]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[6]  (.CLK(clk),
    .D(n_972),
    .QN(quo[6]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[7]  (.CLK(clk),
    .D(n_893),
    .QN(quo[7]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[8]  (.CLK(clk),
    .D(n_900),
    .QN(quo[8]));
 DFFHQNx1_ASAP7_75t_R \u6_quo_reg[9]  (.CLK(clk),
    .D(n_948),
    .QN(quo[9]));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_481));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2414));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_480));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1580));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233843 (.A(n_14271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_478));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233845 (.A(n_14271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_479));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_476));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2120));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_drc_bufs233871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_475));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_474));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2188));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_464));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1860));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_455));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_382));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs233972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2338));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs234010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_451));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs234012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1581));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs234141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_436));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_drc_bufs234214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_428));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_drc_bufs234275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_424));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_drc_bufs234760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2120),
    .Y(n_14012));
 BUFx6f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_473));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt233884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_472));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt233886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_471));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_fopt233897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_466));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_467));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt233927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1727));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_461));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_460));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_459));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_458));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt233982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_454));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt233984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_453));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt233999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_452));
 BUFx4f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_450));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt234023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_449));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_447));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_446));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_441));
 BUFx4f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_440));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234133 (.A(u6_rem_96_22_Y_u6_div_90_17_n_437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_438));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_437));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_435));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_434));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_fopt234189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_432));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_431));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_427));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_421));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_fopt234365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_420));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234375 (.A(u6_rem_96_22_Y_u6_div_90_17_n_417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_419));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234376 (.A(u6_rem_96_22_Y_u6_div_90_17_n_417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_418));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt234378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_462));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_416));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_415));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_417));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt234397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1336));
 BUFx6f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt234401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_414));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt3 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_397));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt4 (.A(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_396));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt5 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_477));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_fopt6 (.A(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_470));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_fopt8 (.A(u6_rem_96_22_Y_u6_div_90_17_n_468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_469));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_fopt9 (.A(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_468));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13733),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13710),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13658),
    .Y(u6_n_149));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13702),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13738),
    .Y(u6_n_148));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13700),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13743),
    .Y(u6_n_145));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214370 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13736),
    .Y(u6_n_147));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214371 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13665),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13728),
    .Y(u6_n_143));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214372 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13608),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13717),
    .Y(u6_n_136));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214373 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13719),
    .Y(u6_n_135));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13718),
    .Y(u6_n_134));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13667),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13730),
    .Y(u6_n_146));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13666),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13726),
    .Y(u6_n_144));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214377 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13644),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13720),
    .Y(u6_n_137));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13729),
    .Y(u6_n_142));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214379 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13662),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13724),
    .Y(u6_n_141));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13634),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13723),
    .Y(u6_n_140));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214381 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13631),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13722),
    .Y(u6_n_139));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13607),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13721),
    .Y(u6_n_138));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13743));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214384 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13599),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13714),
    .Y(u6_n_133));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13713),
    .Y(u6_n_132));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13517),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13712),
    .Y(u6_n_130));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13711),
    .Y(u6_n_129));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214388 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13738));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214389 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13558),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13715),
    .Y(u6_n_131));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214390 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13736));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214391 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13432),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13709),
    .Y(u6_n_128));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13734));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13733));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214394 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13706),
    .Y(u6_n_127));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214395 (.A1(n_14271),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_n_126));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214396 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13730));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214397 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13729));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214398 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13728));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13727));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214400 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13726));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214401 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13725));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13724));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214403 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13723));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214404 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13722));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214405 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13721));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214406 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13720));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214407 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13719));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214408 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13718));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214409 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13717));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214410 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13677),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13366),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13716));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214411 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13552),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13715));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214412 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13714));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214413 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13713));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214414 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13712));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214415 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13711));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13710));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13434),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13709));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13708));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13707));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13706));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B(n_14271),
    .Y(u6_n_76));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214422 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13704));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13703));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13702));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13701));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13700));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214427_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_456));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214429 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13204),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13632),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13697));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214430 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13653),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13696));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214431 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13695));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214432 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13694));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13650),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13693));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214434 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(n_14280),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13692));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214435 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13605),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13691));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214436 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13201),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13606),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13690));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214437 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13645),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13689));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214438 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13688));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214439 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13573),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13687));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B(u6_n_77),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13699));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13686));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13685));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214444 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13684));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214445 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13589),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13683));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214446 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13555),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13682));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214447 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13516),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13681));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214448 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13680));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214449 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2341),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13433),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13679));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13678));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13677));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214454 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13373),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13676));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214455 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13675));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214456 (.A(u6_n_77),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13674));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_494),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13672));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214458 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13301),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13671));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13502),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13670));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214460 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13528),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13669));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214461 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13668));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214462 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13565),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2409),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13623),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13480),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13529),
    .Y(u6_n_77));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13667));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13666));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13665));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13664));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13663));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13642),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13662));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13658));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13629),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13657));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13287),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13656));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214475 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2411),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13655));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13661));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13660));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13659));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214479 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13654));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13653));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13409),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2411),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13410),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13652));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13651));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214483 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13650));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13649));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214485 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13628),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13282),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13648));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13646));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13645));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13644));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214490 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2344),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13643));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2358),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13618),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13642));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214492 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13641));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214493 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13277),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2408),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13640));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214494 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2408),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13647));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214495 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2409),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_372),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2413));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13638));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13639));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214499 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13580),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13541),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13637));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13636));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13618),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13634));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13633));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13632));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13631));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2408),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13630));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214507 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13550),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2412));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2411));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214511 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13591),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2410));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2407),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13629));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214513 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13590),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2397),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13628));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2406),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2360),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13627));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214515 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2378),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13626));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13625));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214517 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13534),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13624));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214518 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13549),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13623));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214519 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13525),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13622));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214520 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13591),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13407),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13590),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13621));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13620));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13615));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13290),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13614));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214525 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13582),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13613));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214526 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13584),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13612));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214527 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13246),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13611));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214528 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13587),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13610));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214529 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13609));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214530 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13401),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13619));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214531 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13400),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13618));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2404),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13616));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2408));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13587),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13608));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13607));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13606));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13605));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13604));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13603));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13602));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13601));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13600));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13599));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214546 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13543),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13444),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_13442),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13442),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13566),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2409));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13598));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214548 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2372),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13307),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13597));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13596));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13554),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13595));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2391),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13594));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214552 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13593));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214553 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2384),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2385),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13468),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13592));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2407));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214558 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2406));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13590));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214560 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13545),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13591));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13589));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13588));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13584));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13582));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13581));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13580));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214569 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13579));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13548),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13578));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214571 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13587));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214572 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2386),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13586));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214573 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2387),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13585));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214574 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13583));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2400),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2405));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214576 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13477),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2404));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13577));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13576));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13534),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13575));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13453),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13574));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13573));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13572));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214584 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2400),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13571));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13544),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13570));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13569));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13567));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13565));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214589 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2358),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13438),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2373),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13322),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13564));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214590 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13319),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13323),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13563));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13247),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13562));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214592 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13404),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13535),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13568));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214593 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2354),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13561));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214594 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13560));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214595 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2359),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2362),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13302),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13566));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13558));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13372),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13557));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13556));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13555));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214600 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13536),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13554));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13553));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13552));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214603 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13420),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13559));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13480),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13551));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2397),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13510),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_13425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13550));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2395),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13405),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13549));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13548));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2403));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214610 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13547));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2396),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13546));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2402));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214616 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13416),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2389),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_13414),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13446),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13416),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13545));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214617 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13544));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2401));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2400));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214622 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13464),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13543));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214623 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13542));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13541));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214625 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13496),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_872),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13540));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13539));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13537));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13533));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214629 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_424),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13529));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13405),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13528));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13527));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214632 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2366),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13472),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13538));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13425),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13526));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13525));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13454),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13536));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2395),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13535));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13421),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13534));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214639 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2379),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13532));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214640 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13381),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13531));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214641 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13414),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13530));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13522));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13520));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214645 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13518));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13517));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13516));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13452),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13515));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13440),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13514));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13471),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2399));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2374),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13524));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13523));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214654 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13424),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13521));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13417),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13519));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214656 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13436),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13513));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214657 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2388),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13512));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13511));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13508));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13506));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13504));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13510));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13503));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214667 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2398));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214668 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_848),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13509));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2397));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2367),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13502));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13507));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214672 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13501));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214673 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13500));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13499));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2360),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13505));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214676 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13498));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2396));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214679 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13238),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13376),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13237),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13495));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214680 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13378),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13237),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13377),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13494));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13493));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13344),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13492));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13437),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13491));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13468),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13490));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13489));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13488));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13475),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13487));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214688 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13366),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_848),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13486));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13497));
 AO211x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13364),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13496));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13484));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13479));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13477));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13475));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13472));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13470));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13467));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13465));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13464));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13380),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13463));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13462));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13461));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13460));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13485));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13459));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13483));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13458));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13482));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13481));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13480));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2387),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13478));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13476));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13474));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13457));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13456));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13473));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13471));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2395));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13469));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13455));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13468));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13454));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13466));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13451));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13449));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13445));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13441));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13439));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13437));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13436));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214743 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13435));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214744 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13231),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13434));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214745 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2342),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13433));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13432));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13263),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13431));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13251),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13430));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13429));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2363),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13428));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13257),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2353),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13427));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2357),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13323),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13315),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13453));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214753 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13236),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13452));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214754 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2371),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13450));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13296),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13448));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214756 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2364),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2394));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13247),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13447));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214758 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13446));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214759 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2346),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2393));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13302),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13444));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2348),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13443));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13322),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13313),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13442));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214763 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13440));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2392));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2368),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13438));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2391));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214767 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2390));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214768 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13195),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13223),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2389));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214769 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2342),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13220),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2388));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13423));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13421));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13419));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13412));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13410));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13408));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13406));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13404));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13402));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13426));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13425));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13401));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13400));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_243),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13424));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2387));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13295),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13422));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13420));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2347),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13418));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2386));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13417));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2354),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13416));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13415));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13414));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2350),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13413));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214799 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13399));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13398));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13397));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2382),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13411));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13409));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13395));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13394));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13393));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13316),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13392));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13391));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13407));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214811 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13390));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13389));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214813 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13388));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13387));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13386));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13385));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13384));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13383));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13382));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2385));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13405));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2384));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214823 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13106),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13403));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13381));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13378));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13376));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13374));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13372));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13370));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13368));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13366));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13365));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12948),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13196),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13364));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214836 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13363));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13362));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13380));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_797),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13361));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13379));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2374),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13360));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13359));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13358));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13357));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_822),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_823),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13356));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13355));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13274),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13354));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2346),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13353));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214849 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13199),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13352));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13276),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13351));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13273),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13350));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13349));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13271),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13348));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13347));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13346));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214856 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_514),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13345));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214857 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13344));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13343));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13342));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13341));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13340));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13339));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13338));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13337));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13377));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214866 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2813),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13336));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214867 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13375));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2363),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13335));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2383));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13373));
 AO211x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13229),
    .C(n_14465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13371));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13369));
 OR3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13160),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13367));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13334));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13331));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13327));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13325));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13324));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13321));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13320));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13317));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13316));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13315));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13313));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13311));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13309));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13308));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214905 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13306));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13304));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13301));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13300));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13298));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13297));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13294));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13293));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13291));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13289));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13288));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13286));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13285));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13284));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13281));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13280));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13333));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13332));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13279));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2382));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13330));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13329));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2381));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13328));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13278));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13326));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2380));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2379));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2378));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2377));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13277));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13323));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2376));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13322));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2375));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13319));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13318));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2374));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2373));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2372));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13314));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13312));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13310));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2371));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2370));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2369));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2368));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13307));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g214969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13305));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13303));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13302));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2367));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13299));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2366));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2365));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13296));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13295));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2364));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13292));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2363));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13290));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2362));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2361));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2360));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13287));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2359));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2358));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2357));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13283));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13282));
 AOI211x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g214991 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13094),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13134),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2356));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13276));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13273));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13271));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13268));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13266));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g214998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13262));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13261));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13260));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13259));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13250));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13246));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13245));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13241));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2344));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13237));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13235));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13234));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2341),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13233));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215022 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2341),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13232));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215023 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2340),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13231));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215024 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12856),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13230));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215025 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13157),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13229));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215026 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13112),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2336),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12660),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_13155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13228));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215027 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13227));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_35),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13226));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13225));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13275));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13274));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13224));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13272));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13223));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13222));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13221));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13270));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13220));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13219));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13218));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13269));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13217));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13267));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13265));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13264));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13263));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2355));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2354));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2353));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2352));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2351));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2350));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13258));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13257));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13256));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13255));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13254));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13253));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13252));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13251));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2349));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2348));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13249));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13248));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13247));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2347));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2346));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13244));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13243));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13242));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2345));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13240));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13239));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13238));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13236));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13215));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13213));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13211));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13209));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13207));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13206));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13203));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13201));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13199));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13197));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13196));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215087 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13072),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13216));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215088 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13097),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13214));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215089 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13095),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13212));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215090 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13062),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13210));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215091 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13073),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13208));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13205));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13204));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215094 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13202));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13200));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215096 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13034),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13198));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13195));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13193));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13191));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13188));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13186));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13183));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215107 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13182));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13181));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215109 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13180));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_494),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2343));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2342));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215112 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13022),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13194));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13192));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13190));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13189));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215116 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13008),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13187));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215117 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_363),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13185));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215118 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13184));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2340));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215123 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13178));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13177));
 AOI221xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215125 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13105),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2336),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12656),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13176));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215126 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_369),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12654),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13175));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215127 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13174));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215128 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13076),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13173));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215129 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13172));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215130 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13074),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13171));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215131 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13170));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215132 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13169));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13168));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215134 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13124),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13167));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215135 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13123),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2284),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13179));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215136 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2341));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215137 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12976),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13166));
 OAI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215138 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13049),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12663),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13165));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215139 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_362),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13164));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215140 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13163));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13161));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215143 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13116),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13160));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215144 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13159));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13158));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13157));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13156));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13155));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13154));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13153));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215151 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13115),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13152));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215152 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2305),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13151));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13150));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215154 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13033),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13149));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215155 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_367),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12657),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13148));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215156 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12726),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13147));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215157 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12639),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13146));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215158 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12661),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13145));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215159 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13046),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13144));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13070),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13143));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215161 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13050),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12644),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13142));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215162 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13045),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13141));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215163 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2339),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13140));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13093),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13138));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215166 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13137));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215167 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2335),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13136));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12818),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13135));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13089),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13099),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_13119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13134));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13133));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13011),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13132));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215172 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13041),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13131));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215173 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13066),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13130));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215174 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12898),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12897),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13129));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215175 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12977),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13128));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215176 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12620),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13127));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13126));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215178 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13125));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13121));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13119));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13118));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13117));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12727),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12753),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13116));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .B(u6_n_79),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13115));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12768),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13114));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12751),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13113));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12972),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13124));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215189 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13123));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215190 (.A(u6_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13122));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13078),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13120));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13084),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13112));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13111));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215194 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12823),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13086),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13110));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215195 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_365),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13109));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13082),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13108));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13107));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13085),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13106));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13105));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215202 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12746),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13104));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215203 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13103));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13101),
    .Y(u6_n_79));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13099));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2293),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13098));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215210 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12970),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2339));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215211 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13017),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13035),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13101));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215212 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13023),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13100));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13097));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13063),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13096));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13064),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13095));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13094));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215217 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13068),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12747),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13093));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215218 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12727),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13092));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13089));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215222 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13044),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12940),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13087));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13086));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215224 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2333),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2282),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13085));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215225 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2281),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13084));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215226 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2332),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13083));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12763),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13082));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215228 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12756),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13059),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13081));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215229 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13091));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13052),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13090));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12956),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13088));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215237 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13079));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2335));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2336));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13077));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13076));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13075));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13059),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13074));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13073));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13072));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13071));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13054),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13070));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13051),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13069));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13058),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12883),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13080));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13078));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215252 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2318),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13068));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215253 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_366),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12869),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13067));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215254 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12735),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2285),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13066));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215255 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12954),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13065));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215257 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2319),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2334));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215258 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12762),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13064));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215259 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12684),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13063));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13062));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13061));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13059));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2331));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13057));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215270 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12990),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13056));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215271 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12755),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13055));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215272 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12698),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13054));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215273 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13030),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13053));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13052));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215275 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12851),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2333));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215276 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12878),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2332));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215277 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12880),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13060));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215278 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13058));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215279 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12965),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13029),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2330));
 OAI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215280 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13000),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12995),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13013),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2316),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13051));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13028),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13050));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215282 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2324),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12830),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_13030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13049));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12813),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13048));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13047));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13046));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13045));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12993),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13044));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13043));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215289 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12694),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13042));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13041));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13040));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215292 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2283),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12988),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2289),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12927),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13039));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215293 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13010),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12904),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13038));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2329));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13037));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215299 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13004),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13036));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2328));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215303 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12966),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13035));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13034));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13033));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13031));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13030));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2324));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215313 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2275),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13028));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215314 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12727),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12753),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12702),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2327));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215315 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2305),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12703),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2326));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215316 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2322),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2271),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13027));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2325));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215318 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2322),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12939),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13032));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215319 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2314),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_12882),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12882),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2320),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13029));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13026));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215322 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12908),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13025));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215323 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12907),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13024));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12962),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13023));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13022));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12691),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_13002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13021));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2323));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2281),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2287),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12742),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13020));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215331 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12764),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12770),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13019));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13018));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12953),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13017));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215335 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2274),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12987),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13016));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215336 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12978),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13015));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13014));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12997),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13013));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13012));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12987),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13011));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215341 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12732),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12992),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13010));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12975),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13009));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12974),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13008));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215344 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12934),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13007));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13006));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2322));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215350 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2309),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2315),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_12881),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12881),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12906),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13005));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2321));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2308),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12900),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_12873),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12873),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12905),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13004));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12947),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12922),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13003));
 OA21x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2314),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13001));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12951),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13000));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12858),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_866),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12999));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12998));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12996));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12994));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12991));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12989));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12884),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12872),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12986));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215367 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12985));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12947),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12984));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2291),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12997));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12971),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12995));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12927),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12993));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215372 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12924),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12992));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12967),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12904),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12990));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12988));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2315),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12987));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12982));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12980));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12977));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12976));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12887),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12983));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2320));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215384 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12902),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12975));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12974));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12901),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12973));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12886),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12981));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215388 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12874),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12979));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215389 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12978));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12972));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12970));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12968));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12966));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12934),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12965));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12964));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12907),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12875),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12963));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12962));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215398 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12856),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12971));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12961));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12960));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12969));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12932),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12959));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12967));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12958));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12956));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12954));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12952));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12950));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12892),
    .B(n_13848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12946));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12792),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12945));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215412 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2300),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12957));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12955));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12953));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12944));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2261),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12951));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12949));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2450),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12948));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12943));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12629),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12817),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_432),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12947));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12939));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12936));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12931));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12930));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12928));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12926));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12923));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12922));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12921));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12942));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12941));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2319));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2318));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12940));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12938));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12920));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12937));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12935));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12883),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12934));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2317));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12933));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215446 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12726),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12919));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215447 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12726),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12918));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12917));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12932));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2316));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12929));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12927));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12925));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12924));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12916));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12912));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12910));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12903));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12902));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12901));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2313));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215468 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12667),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12899));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12796),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12898));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12709),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12897));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215471 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12896));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215472 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12895));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12683),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12894));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12893));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215475 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12583),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12892));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2273),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12666),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12891));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12688),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12890));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215478 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2286),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12889));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215479 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12888));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215480 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2295),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12915));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2276),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12914));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2272),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12913));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2260),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12911));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215484 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2270),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12909));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12758),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2282),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12908));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12879),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12907));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215487 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12695),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12906));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215488 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12687),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12905));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12904));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215490 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2278),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2315));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12710),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2314));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215492 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12670),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12671),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12900));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12885));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12880));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12878));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12875));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12871));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12870));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12866));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12864));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12862));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12860));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12858));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12856));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12855));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12854));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12853));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12852));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12851));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_243),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12887));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12886));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12850));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12884));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12883));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12772),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12882));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12881));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215521 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12661),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12879));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12877));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2271),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12876));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12874));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12688),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12873));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12872));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2312));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12869));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12849));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12848));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12868));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12744),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12867));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12847));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12846));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12752),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12845));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215536 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12844));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12843));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12842));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12764),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12841));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12840));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2295),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12865));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12839));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12838));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12837));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12836));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12835));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12834));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12863));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12861));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12655),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2311));
 AO211x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_432),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_360),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12609),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12859));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215552 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12556),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12857));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12833));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12831));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12829));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12827));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12821));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12819));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12818));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12622),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12817));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12816));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12815));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12814));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12813));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12783),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12812));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12784),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12811));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12810));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12809));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12832));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12808));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12807));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12806));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12805));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215582 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12804));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12803));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12802));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2273),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12801));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12830));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2272),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12800));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12799));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12798));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12797));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12828));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12716),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12826));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2275),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12825));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12796));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12824));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215596 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12634),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12795));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2310));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215598 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12635),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12794));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2309));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215600 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12793));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215601 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12630),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12792));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2308));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12791));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215604 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_754),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2818),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12790));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12789));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12690),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12788));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12787));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12823));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12822));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_830),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2307));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12820));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12786));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12782));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12779));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12776));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12774));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12773));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12771));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12769));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12768));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12765));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12763));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12762));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12760));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12759));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12758));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12756));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12755));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12752));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12751));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12750));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12749));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12748));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12745));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12744));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12742));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12739));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12738));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12737));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12734));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2285),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12733));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12732));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12730),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12731));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12729));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2281));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12726));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2279));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12785));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12724));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12784));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12783));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12781));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12780));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12778));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12777));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2306));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12723));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12722));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12775));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2305));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12772));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12770));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2304));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12767));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12766));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12764));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2303));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2302));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2301));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2300));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12761));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2299));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2298));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12757));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2297));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2296));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2295));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2294));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12754));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2293));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12753));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2292));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2291));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2290));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2289));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2910),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2288));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12747));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12746));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12743));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12741));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12740));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2287));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2286));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12736));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12735));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2285));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2284));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2283));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12730));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2282));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12728));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12727));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2280));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215740 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12725));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12720));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12718));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12716));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12714));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12711));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12709));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12707));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12705));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12701));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12700));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12699));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12697));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12696));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12693));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12691));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12690));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12689));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12686));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12685));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12684));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12681));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12680));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12679));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12601),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12555),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12678));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12677));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12580),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12676));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12675));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12721));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12719));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12717));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12715));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2278));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12713));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215799 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12712));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12710));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12674));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12673));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12672));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12671));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12670));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12708));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12706));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12669));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12668));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12704));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12703));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12702));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2277));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2276));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2275));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2274));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12698));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2273));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2272));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12667));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2271));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2270));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2269));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12695));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12694));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12666));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12692));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2268));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2267));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2266));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2265));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2264));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2263));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12688));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2262));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12687));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2261));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2260));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12665));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2259));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2258));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12683));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12682));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12663));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12661));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12659));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12657));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12655));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12653));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12650));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12648));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12646));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12644));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12642));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2257));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12639));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12664));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12662));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12660));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215863 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_358),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12658));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12656));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12654));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12618),
    .B(n_14466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12652));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12651));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215868 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12486),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12487),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12649));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215869 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12461),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12463),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12647));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12645));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12441),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12643));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12411),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12641));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215873 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12640));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12637));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12635));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12633));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12630));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12629));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215880 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12628));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215881 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_436),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12627));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215882 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12626));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12625));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12624));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215887 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12622));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2256));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12638));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12636));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215891 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12558),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12634));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215892 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12632));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215893 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12631));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12620));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215895 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12619));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215896 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12618));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215897 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12617));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215898 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12526),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12616));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215899 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12615));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215900 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12614));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215901 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12613));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215902 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12562),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12612));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12611));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12610));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12621));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12609));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215907 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12608));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215908 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12409),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12607));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215909 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12606));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215910 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12605));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215911 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12473),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12604));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215912 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12603));
 OAI33xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215913 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_12549),
    .B1(u6_n_81),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .B3(u6_rem_96_22_Y_u6_div_90_17_n_12369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12602));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12601));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12600));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215916 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12599));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215918 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_436),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12543),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12597));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215919 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12056),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12596));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215920 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12539),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12595));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215921 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12594));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215922 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12521),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12593));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215923 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12075),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12484),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12592));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215924 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12517),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12591));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215925 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12462),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12590));
 AOI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215926 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12525),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12077),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12589));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215927 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12488),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12588));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12490),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12587));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215930 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12544),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12585));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215931 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12584));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215932 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12542),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2240),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12598));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12583));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12579));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215935 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_436),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12578));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215936 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12443),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12577));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215937 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12439),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12576));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12481),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12575));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12574));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12573));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215941 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12552),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12572));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12571));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12512),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12570));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215945 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12547),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12568));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12567));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_357),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12582));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215948 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12060),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12581));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215949 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12355),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12047),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12580));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12565));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12563));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12562));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215953 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2228),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12561));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12560));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .B(u6_n_81),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12566));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12564));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12559));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12558));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12541),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12557));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12556));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12555));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12554));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12553));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12552));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12505),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12196),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12296),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12551));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215967 (.A(u6_n_81),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12549));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215968 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12535),
    .Y(u6_n_81));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12547));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12548));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12363),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12546));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215972 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2214),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12545));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215973 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12510),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12544));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215974 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12263),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12510),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12262),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12543));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12541));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12483),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12539));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12538));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12537));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12536));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12489),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12535));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12534));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215983 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12533));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215984 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12532));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215985 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2210),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12531));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215986 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12161),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12530));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12529));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215988 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12504),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12528));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215989 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12542));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215990 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12540));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g215991 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2243),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12417),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12480),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12449),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12527));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12526));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12525));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12524));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12523));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12522));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12521));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g215998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12520));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g215999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12519));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12518));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12517));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12516));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12515));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12514));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12513));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216006 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12184),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12512));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216007 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12187),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12294),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12511));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12509));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216009 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12510));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12507));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216011 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12508));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216014 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12502));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12501));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216016 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12135),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12500));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12177),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12499));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216018 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12498));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216019 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12471),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12497));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216020 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2195),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12467),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12496));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12274),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12506));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216022 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12300),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12470),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12505));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216023 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12318),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2255));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216024 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12312),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12504));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216025 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12347),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2254));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216026 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12503));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12494));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12493));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12492));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12471),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12491));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12490));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216033 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12415),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12489));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12488));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12487));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12486));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12485));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12467),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12484));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216039 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12102),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12483));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216040 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12398),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12495));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12482));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12481));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216043 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12367),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12480));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216044 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2234),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12428),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12288),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12365),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12479));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12478));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12477));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216047 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12454),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12476));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12457),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12343),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12436),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12475));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12452),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12474));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12473));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12472));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12471));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12469));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12467));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2249));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2250));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12356),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12402),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12466));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216065 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2253));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216066 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2252));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216067 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12431),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12470));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216068 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12432),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2251));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216069 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12468));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216070 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2248));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12464));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12432),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12463));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12435),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12462));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12461));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216076 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12460));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216077 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12459));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216078 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12458));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216079 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2247));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216080 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12431),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12316),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12465));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216082 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12397),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12423),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12455));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216083 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12286),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12454));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12416),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12344),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12453));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216085 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2200),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12452));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216086 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12118),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12451));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216087 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12109),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12450));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216088 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12179),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12421),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12457));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216089 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2210),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2216),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12191),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12456));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216090 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12158),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2215),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12178),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2246));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12449));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216092 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12425),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12447));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216093 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12381),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12446));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216094 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12384),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12445));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12444));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12443));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12442));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12441));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12440));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12420),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12439));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216101 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12448));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12347),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12438));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216103 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12437));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216104 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12160),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2223),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12436));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12435));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216106 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12359),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12434));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12432));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216108 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12358),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2236),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12433));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12431));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216110 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12430));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12423),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12429));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12426));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12422));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216116 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12335),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12421));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216117 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2237),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12420));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216118 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2236),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12419));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216119 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2238),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2203),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12418));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216120 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2226),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12362),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12428));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216121 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12364),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12427));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12417));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216123 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2219),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12425));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2236),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12424));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216125 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2237),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2245));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216126 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12308),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2244));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216127 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12423));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12416));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12411));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12410));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2236),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12409));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12348),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12408));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216134 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12333),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12407));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216135 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12341),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12406));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216136 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12405));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216137 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12346),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12404));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2240),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2234),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12415));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216139 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12290),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2243));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216140 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12339),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12414));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12364),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12287),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12413));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216142 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12412));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12381),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12401));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12400));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12399));
 NAND2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12398));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12397));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12403));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12363),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12395));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12394));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12402));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12393));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12392));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12391));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12390));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216158 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11940),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11542),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12250),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12389));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12388));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12387));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12386));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12385));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12383));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12379));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12374));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216168 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12372));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216169 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12369));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12367));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12363));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12362));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12360));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12359));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12306),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12358));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12357));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12356));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216179 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12355));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12315),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2242));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12384));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2241));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216183 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12382));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12354));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12381));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12380));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12353));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12378));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12377));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12376));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12375));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12352));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12373));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12371));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12370));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216196 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12097),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12368));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12366));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12365));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12364));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2240));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12053),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12361));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12351));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12345));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12342));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12340));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12336));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12334));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12332));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12330));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12328));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2237));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216220 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12163),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12326));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216221 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12183),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12175),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12325));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216222 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12199),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12324));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216223 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12123),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12323));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216224 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12114),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12322));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216225 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12129),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12321));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216226 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12165),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12320));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12136),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12319));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216228 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12172),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12103),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12350));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12179),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12349));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12348));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2210),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2232),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_12191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12347));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2202),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12346));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12284),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12344));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12343));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2204),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12139),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12341));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12126),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2208),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12339));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12189),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12338));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216238 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12190),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12337));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216239 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12112),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12335));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216240 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12333));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216241 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2231),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12331));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216242 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2230),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2239));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12121),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12329));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2238));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12089),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12327));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2236));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12316));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12310));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12307));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12303));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12299));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12297));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12295));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12293));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12290));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12289));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12286));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12285));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12284));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12283));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12282));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12187),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12318));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12317));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12315));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2235));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12196),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12314));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12313));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12312));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216272 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12311));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12309));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2203),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12308));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12306));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12305));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12304));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12281));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12280));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12279));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12302));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12278));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216283 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12066),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12277));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12301));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12300));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12276));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216287 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12157),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12275));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12274));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12273));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12298));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216291 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12084),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12296));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12272));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12271));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12270));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12269));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12268));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12294));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12188),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12267));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12266));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216300 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12265));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12264));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12292));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12291));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12288));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12287));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2234));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12263));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12261));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12258));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12256));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12253));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12251));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12050),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12250));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12049),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12249));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216316 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_356),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12248));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12247));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216318 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12246));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216319 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12245));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216320 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12244));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216321 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12243));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216322 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12242));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12262));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12241));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12240));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216326 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_12066),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12239));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_209),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12238));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216328 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12237));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12236));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12235));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12234));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12233));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12232));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_514),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12231));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12230));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12229));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2208),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12228));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12227));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12226));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12225));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12224));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216342 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12058),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_830),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12223));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_514),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12222));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12221));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12220));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12260));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2196),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12259));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12060),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12219));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216349 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12218));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12217));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12216));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12215));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2233));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12060),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12214));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12257));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216356 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12255));
 NOR3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12054),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12051),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12254));
 OA211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216358 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12024),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12055),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12252));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12213));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12211));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12209));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12207));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12204));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12201));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12200));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12198));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216374 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12197));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12195));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12194));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12193));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12188));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216386 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12186));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12184));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12182));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12180));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12177));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12176));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12174));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12173));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12171));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12169));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12168));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12166));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12164));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12161));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12160));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12159));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12157));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12155));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12154));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12212));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12153));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12210));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12208));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12206));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12152));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12205));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12203));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12202));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12151));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12150));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2232));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2231));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2230));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2229));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12199));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2228));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2227));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2226));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12196));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2225));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2224));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2223));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12192));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12191));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12190));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12189));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2222));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2221));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12187));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12185));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12183));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12181));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12179));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12178));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2220));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12175));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2219));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2218));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2217));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12172));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12170));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2216));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12167));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2215));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2214));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12165));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12163));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12162));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2213));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2212));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2211));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2210));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12158));
 OA211x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216471 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12011),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_12044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12156));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12149));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12147));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12145));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12143));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12137));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12135));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12133));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12131));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12130));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12128));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12125));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12122));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12120));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12118));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12117));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12115));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12113));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12111));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12109));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12108));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12106));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12104));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12102));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12046),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12045),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12100));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216515 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12099));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216516 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12098));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216517 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12097));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12096));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12148));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12146));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12095));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_25),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2209));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12144));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12094));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12142));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12093));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12141));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12140));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12092));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12091));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12090));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12089));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12088));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12139));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_79),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12138));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2208));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2207));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12136));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12134));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2206));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12132));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2205));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2204));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2203));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2202));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12129));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12127));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12126));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12124));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12123));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12121));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2201));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2200));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12119));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_25),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2199));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12116));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2198));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2197));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12114));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12112));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12110));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2196));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12107));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_25),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12105));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2195));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12103));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2194));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2193));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12101));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12087));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12084));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12082));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12080));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12077));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12075));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12073));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12071));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12068));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12066));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_49),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2192));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2191));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216586 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11890),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12086));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216587 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11949),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12085));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216588 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11920),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12083));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12081));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12079));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11922),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12078));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216592 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_354),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12076));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216593 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11908),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12074));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216594 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11878),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12072));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216595 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11952),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12070));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12069));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11982),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12067));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12062));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12060));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12058));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12056));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12055));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216603 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12013),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11512),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12054));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12053));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216606 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12052));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12051));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216608 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11610),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12050));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216609 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2125),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12049));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216610 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11779),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12065));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216611 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11825),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12064));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216612 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12063));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216613 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12061));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12059));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216615 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11875),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12057));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12047));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216617 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11640),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12046));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11815),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12045));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216619 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12044));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216620 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11980),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12043));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216621 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11954),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12042));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216622 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12041));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216623 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12040));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12039));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216625 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12038));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216626 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11918),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12037));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216627 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12036));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216628 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12035));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216629 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12048));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216630 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_49),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12034));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216631 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12033));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216632 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12032));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216633 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12031));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216634 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12030));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216635 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12029));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12028));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12027));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216638 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12026));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216639 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12025));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12024));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12023));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12022));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216643 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11940),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11602),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11983),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12021));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12018));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11600),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12017));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216647 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11971),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12016));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12004),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .Y(u6_n_82));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12014));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11702),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12020));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2190),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2165),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_11621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12019));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12013));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12012));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12011));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11977),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11976),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12010));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11992),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12009));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12008));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12007));
 INVx5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12005));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12004));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216661 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11526),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12003));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216662 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11507),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12002));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216663 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12001));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216664 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11516),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12000));
 AOI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216665 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_355),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2188),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11521),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11999));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216666 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11998));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216667 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11919),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11997));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216668 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11996));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216669 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11622),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11995));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216670 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11606),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11994));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216671 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11993));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216672 (.A(u6_n_83),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12006));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216673_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_444));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11992));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216675 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11872),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11991));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216676 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11494),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11990));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216677 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11826),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11989));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216678 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11847),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11496),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11988));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216679 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_474),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11987));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11986));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11985));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11984));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11983));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11982));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11981));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11980));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216687 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2185),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_475),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11979));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11978));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216689 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11605),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11646),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11977));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11935),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11760),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11976));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11974),
    .Y(u6_n_83));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216692 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11860),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11974));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216693 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11973));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216694 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11561),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2187),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11972));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2187),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11971));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11944),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11970));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2190));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11966));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11965));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11964));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11963));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11962));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216706 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11608),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11961));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216707 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11544),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11939),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11960));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216708 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11959));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216709 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2153),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11958));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216710 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11628),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11957));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216711 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11969));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216712 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11819),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2189));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216713 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11932),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11968));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216714 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11884),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11967));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11956));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11955));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11954));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11928),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11953));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11952));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11951));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11950));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11931),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11949));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11930),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11948));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11947));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216728 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11832),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11907),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11897),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11823),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11946));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11945));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216731 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11912),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2187));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216732 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2127),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11944));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216733 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11881),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11898),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11863),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11943));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11942));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11940));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216736 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11855),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11901),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11941));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11937));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2186));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216743 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11829),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11934));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216744 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11933));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11932));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2183),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11931));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11896),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11930));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11894),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11929));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11901),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11928));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11927));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11905),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11939));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2183),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11744),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11938));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216753 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2177),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11936));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216754 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11802),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11935));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11925));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11894),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11923));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11922));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11921));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11730),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11920));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11906),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11919));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11903),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11918));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11887),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11917));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11916));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11915));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216766 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11904),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11914));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216767 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11776),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11926));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216768 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2182),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11924));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11913));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11912));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11911));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11798),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11910));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11880),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11909));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11667),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11908));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11906));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11905));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11903));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11900));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216783 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11899));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216784 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11706),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11898));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216785 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11707),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11897));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11647),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11650),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2184));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11907));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11870),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2183));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2181),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11904));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2175),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11902));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11839),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11901));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11893));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11892));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11891));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11890));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11869),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11889));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216798 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11888));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2181),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11887));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11792),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11896));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11895));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11770),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11894));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11886));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11831),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11884));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11545),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2137),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11551),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11883));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11609),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11634),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11638),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11882));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11830),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11881));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2141),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2143),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11620),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11885));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11880));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216810 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11566),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11879));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11878));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11877));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11876));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11875));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11849),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11836),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11874));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11873));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11872));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2179),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11871));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11870));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11869));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11868));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2181));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216828 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11604),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11865));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216829 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11842),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11864));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216830 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11786),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11812),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2182));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216831 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11811),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11867));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11866));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2178),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11862));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11861));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11823),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11860));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11834),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11859));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11841),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11863));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11833),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11752),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2180));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11749),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11857));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_424),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11856));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11855));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216844 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11854));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11570),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11853));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216846 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2133),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11852));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216847 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11716),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11858));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11851));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216851 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11765),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11848));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11847));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216854 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11766),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2170),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11767),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11846));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11787),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11845));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216856 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11844));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216857 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11850));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216858 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11793),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11849));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11711),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2179));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11840));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11839));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11838));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11837));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216866 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11747),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11836));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216867 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2178));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2159),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2142),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2177));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11843));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2145),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11750),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11842));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11541),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11699),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11841));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11835));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11831));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11828));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11826));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11825));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2169),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11824));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216880 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2126),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11834));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216881 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2176));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216882 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11587),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11833));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11807),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11832));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11701),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2125),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11830));
 NAND4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2166),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2140),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11829));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216886 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2160),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11827));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11821));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11819));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11817));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11815));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216892 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11813));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11812));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11811));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216895 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11810));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11809));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11808));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11807));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11823));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11822));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2175));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11764),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11806));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11820));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11805));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216905 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11804));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11758),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11803));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216907 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11802));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11818));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11801));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11800));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11799));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11816));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11814));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11794));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11792));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11790));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11788));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2171));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2168));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216933 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11617),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11785));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216934 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2134),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11784));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216935 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2130),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11783));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216936 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_348),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11782));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216937 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11528),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11781));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11780));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216939 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11502),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11779));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216940 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2174));
 NAND4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11629),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11609),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11798));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11555),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11797));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11585),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2173));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11778));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11616),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2141),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2172));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11549),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11545),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11796));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216947 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11579),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11795));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216948 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2163),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11793));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216949 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11791));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216950 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11499),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11789));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216951 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2132),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11787));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2170));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216953 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2169));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11501),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11532),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11786));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11774));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11767));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11764));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11761));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11758));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11756));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11754));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11753));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11751));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2165));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11748));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11747));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11746));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11777));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11776));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11745));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11744));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11775));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11773));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11743));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11772));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11742));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11771));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g216982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11770));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216983 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11741));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g216984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11769));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216985 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11768));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11766));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11765));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11740));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11763));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11739));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11738));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11737));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11762));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11736));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11735));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11760));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11734));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11733));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g216999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11732));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2440),
    .B(n_14028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11759));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11731));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11730));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217003 (.A(n_14028),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11757));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11729));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11728));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11727));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217007 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11523),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11726));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11725));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11724));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11723));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11722));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11721));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2440),
    .B(n_14028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11755));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2167));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11512),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11752));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2166));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11750));
 OA211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217018 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11484),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11749));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11719));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11716));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11711));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11708));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11706));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11704));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11701));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217029 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11252),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11503),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11700));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217030 (.A1(n_14019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11485),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11133),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11699));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11698));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217032 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11697));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217033 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11696));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217034 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11695));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11720));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11694));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11718));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_130),
    .B(n_14028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11717));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11693));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11692));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11691));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11690));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217043 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11512),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11689));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11688));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2137),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11687));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11686));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11685));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11684));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11683));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11682));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11715));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11681));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217053 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11488),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11680));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11679));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11678));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11677));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11676));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11675));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11714));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11674));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11713));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217062 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11673));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11712));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11710));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217065 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11494),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11672));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11671));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217067 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11493),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11670));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217068 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11669));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217069 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_502),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11709));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11668));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217071 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_514),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11667));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217072 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11666));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11707));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2164));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11705));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_130),
    .B(n_14028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11703));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11702));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11665));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11663));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11661));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11658));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11656));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11654));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11652));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11649));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11646));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11645));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11644));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11642));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11641));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11640));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11639));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11637));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11636));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11635));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11633));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11631));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11629));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11628));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11626));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11625));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11624));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217126 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11621));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11619));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11618));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11616));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11614));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11610));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11608));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11606));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11605));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11604));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11602));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217144 (.A(n_14028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11600));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11664));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11662));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11660));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11599));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11598));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11597));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11659));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11657));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11655));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11653));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11651));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11650));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11648));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2163));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11647));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2162));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2161));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11643));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2160));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2159));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2158));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2157));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2156));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217168 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2155));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217169 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11638));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2154));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2153));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2152));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2151));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11634));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11632));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2150));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11630));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2149));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2148));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11627));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2147));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2146));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11623));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11622));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11620));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2145));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2144));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11617));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11615));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2143));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11613));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11612));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11611));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11609));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11607));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2142));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2141));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2140));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217199 (.A(n_14026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11603));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217201 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11594));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11592));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11589));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11588));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11586));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11584));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11582));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11581));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11578));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11576));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11574));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11573));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11571));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11570));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11568));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11567));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11564));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11563));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11562));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11561));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11559));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217237 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11557));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11556));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11554));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11552));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11549));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11547));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11544));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11542));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11541));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11540));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11539));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_389),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11538));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11596));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11595));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11593));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11537));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11591));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11536));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11535));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11534));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11533));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11532));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11590));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11531));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11530));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2139));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11587));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11585));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2138));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11583));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2137));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2136));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217272 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11579));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11577));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11529));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11575));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2135));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11572));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2134));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2133));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2132));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11569));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2131));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2130));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11566));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11565));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2129));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2128));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2127));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11560));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11558));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11528));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2126));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11475),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11555));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11448),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11553));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11551));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11550));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11548));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11527));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11546));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11545));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2125));
 OA221x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217303 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_396),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11161),
    .C(n_14025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11543));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11525));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11523));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11521));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11518));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11516));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11515));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11512));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11510));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11508));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11506));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11504));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11503));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11351),
    .A2(n_14019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11526));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11471),
    .B(n_14017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11524));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11470),
    .B(n_14032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11522));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11459),
    .B(n_14020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11520));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217321 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11469),
    .B(n_14018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11519));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217322 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11468),
    .B(n_14023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11517));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11466),
    .B(n_14022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11514));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11478),
    .B(n_14030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11513));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217325 (.A(n_14015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11511));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217326 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11367),
    .A2(n_14019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11509));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11309),
    .A2(n_14019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11507));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217328 (.A(n_14031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11505));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11502));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11500));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11498));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2124));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217334 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11495));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11493));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11491));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11488));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11486));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11485));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11484));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217342 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11414),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11401),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11394),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11482));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217343 (.A1(n_14014),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11481));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11501));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11464),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11499));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11497));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217347 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11147),
    .A2(n_14019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11496));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11464),
    .B(n_14029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11494));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217349 (.A1(n_14019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11492));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11452),
    .B(n_14493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11490));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217351 (.A(n_14021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11489));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217352 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11275),
    .A2(n_14019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11487));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11479));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11478));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11477));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217356 (.A1(n_14019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11476));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2123),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11475));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217358 (.A1(n_14014),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11474));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_346),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11473));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11472));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11354),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11471));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217362 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11470));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217363 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11469));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217364 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_347),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11468));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217365 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11400),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10905),
    .B2(n_14012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11467));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11466));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .B(u6_n_84),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11480));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11463));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11272),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11461));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217370 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11460));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217371 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11295),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11459));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217372 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11458));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217373 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11457));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11456));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_343),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11455));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11387),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11454));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11453));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11452));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11451));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2106),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11465));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217381 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11188),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11464));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11462));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11410),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11450));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11449));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11104),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11446));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .A2(n_14012),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11187),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11445));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .A2(n_14012),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_223),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11444));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217388 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .A2(n_14012),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11373),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11443));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217389 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11372),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10910),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11442));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217390 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11341),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11441));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217391 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .A2(n_14012),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11340),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11440));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217392 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11439));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217393 (.A1(n_14012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10915),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11438));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11382),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11437));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217395 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10982),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11386),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11436));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217396 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11366),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11435));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217397 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .A2(n_14012),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11308),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11434));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217398 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11305),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11433));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10897),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11273),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11432));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217400 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_344),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .B2(n_14012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11431));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11448));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2107),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11430));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_397),
    .B(n_14019),
    .Y(u6_n_84));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217405 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11229),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_477),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11428));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11427));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11420));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11414));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11413));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11412));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11409));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11147),
    .B(n_854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11406));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11141),
    .B(n_854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11405));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217427 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11214),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11410));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217428_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_423));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217429_dup (.A(n_14012),
    .B(n_854),
    .Y(n_14024));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11403));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11402));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11401));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11400));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11399));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217436 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11404));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217437 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2123));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11394));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217442 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2097),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11393));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11392));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217444 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11391));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217445 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11211),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11398));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217446 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11329),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11396));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11395));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11357),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11390));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11389));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11388));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11387));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11360),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11386));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11362),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11385));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11383));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .B(n_14012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11381));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .B(n_14012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11380));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217457 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11379));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11384));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11378));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2096),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11377));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217461 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11376));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217462 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11349),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11375));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11382));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11344),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11374));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11346),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11373));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11372));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11371));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11370));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11338),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11369));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11368));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11367));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11350),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11366));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11278),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11335),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11277),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11365));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11363));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11362));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11359));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217478 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10995),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11358));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217479 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10988),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11357));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11106),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11364));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11251),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2121));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11361));
 OAI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11312),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11224),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_11169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11360));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11355));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11354));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11353));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11352));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11351));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11356));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217494 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11300),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11110),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11348));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217495 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11017),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11015),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11347));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217496 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11314),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11346));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217497 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11311),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11345));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217498 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11224),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11350));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217499 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11239),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2119));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217500 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11311),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2118));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217501 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11098),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11349));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217502 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11344));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11343));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217504 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11342));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11341));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11055),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11340));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11339));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217509 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11338));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217510 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11337));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2106),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2110),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11191),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11336));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217513 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11335));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217514 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11306),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11334));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217515 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2107),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2109),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11194),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11333));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217516 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11008),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11332));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217517 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11300),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2117));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11330));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11328));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11298),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11327));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217523 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10990),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11326));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11297),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2086),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11325));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217525 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11297),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11331));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217526 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11209),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11329));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11324));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11320));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217530 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11077),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11318));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11317));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11316));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11315));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217535 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10993),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11004),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11107),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11323));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217536 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10987),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10996),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11109),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11322));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11174),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11321));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11312));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11311));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2116));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11280),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11309));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11308));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217545 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11139),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11307));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11245),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11306));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11305));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11281),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11304));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217549 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11303));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11097),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11314));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11287),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11208),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11313));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217552 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11207),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11310));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11299));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11298));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11257),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11296));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217558 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11269),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11302));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217559 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11100),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11301));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217560 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11267),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11300));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217561 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11297));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11295));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217563 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11140),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11233),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11026),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11294));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217564 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11261),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11293));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217565 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11143),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11292));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217567 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11269),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11290));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2115),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11288));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217570 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2115));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217571 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11007),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11286));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11285));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11082),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11284));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217574 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10937),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2068),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10944),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11283));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11181),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11219),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11282));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217576 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11281));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11011),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11289));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_342),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11280));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11137),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11117),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_11074),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11196),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11117),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11287));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11279));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11277));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_342),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11275));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11274));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11273));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11272));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217588 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2111),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11271));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217589 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11250),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2076),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11270));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217590 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11169),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11278));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11234),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_872),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11276));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11269));
 AOI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217593 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11118),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11075),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2100),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2103),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11118),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11268));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11266));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11267));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217596 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11265));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11264));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217598 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2097),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11263));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11262));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217600 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2094),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11261));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11260));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217602 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2098),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11259));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2111),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11258));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11257));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11191),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11212),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2106),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11256));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11255));
 NOR3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11192),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11254));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11210),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2107),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_11106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11253));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11106),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11248));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11247));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11246));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11245));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11244));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11243));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11242));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11241));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11240));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11252));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11251));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11239));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217625 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11074),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11250));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217626 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11075),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2100),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11249));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11238));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11236));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11234));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217635 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10995),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11233));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2105),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11232));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2104),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11231));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2100),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11230));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11229));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217640 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11228));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217641 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2084),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2114));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217642 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2089),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2113));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217643 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2100),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11227));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217644 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2101),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11226));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217645 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11237));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2071),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11225));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217647 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11235));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217648 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2092),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2112));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11068),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11131),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2111));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11224));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11222));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11220));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11214));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11212));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11210));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11139),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11209));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11208));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11207));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11223));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11221));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11219));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11206));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11205));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11218));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11204));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11217));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11216));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11175),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11203));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11202));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11215));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11213));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11211));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11200));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11193));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11076),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11190));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217676 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11189));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11201));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11188));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11187));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11186));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217682 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2081),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11185));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11184));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11183));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11199));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11198));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11197));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217688 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10960),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11196));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11195));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11194));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11192));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11191));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11182));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11180));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11178));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11174));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11172));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11171));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11168));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11167));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11166));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11162));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11160));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11181));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11159));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217711 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11158));
 AND4x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11013),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11003),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11179));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2094),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11157));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11156));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11155));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11177));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11176));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11175));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11154));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11153));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10939),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10957),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11173));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11152));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2110));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11170));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11169));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2109));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11165));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11164));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2108));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2107));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11163));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2106));
 AND3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10883),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11161));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11150));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11146));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11138));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2102));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2101));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11135));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11133));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11132));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217753 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10655),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10896),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10981),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11131));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217754 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10934),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10385),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11130));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2065),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10976),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11129));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217756 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2093),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11128));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217757 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2074),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10939),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11127));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217758 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11126));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217759 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10964),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11151));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217760 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2085),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2105));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11149));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217762 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2067),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11148));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217763 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11001),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_340),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2104));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217764 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10931),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2062),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11147));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11145));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217766 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10999),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11144));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10937),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10944),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11143));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217768 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10962),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2103));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11142));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217770 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10932),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2063),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11141));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10995),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11140));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10988),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11139));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10924),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10923),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11137));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2062),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10925),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11136));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217775 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2063),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2100));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10930),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10935),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2099));
 AO211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217777 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10772),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11134));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11125));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11123));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11121));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11115));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11113));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11111));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11108));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11104));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11102));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11124));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11101));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11122));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11100));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11120));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11099));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11098));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11097));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11119));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11118));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11117));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2082),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11096));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10912),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11095));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11116));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2085),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11094));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11093));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11114));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11034),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11092));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11091));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11090));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11112));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10997),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11089));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11088));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2084),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11087));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11086));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11085));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11007),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11084));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11083));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11110));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2098));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11109));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2097));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2096));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11107));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11106));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11105));
 AND3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10827),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11103));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11082));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11080));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11072));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11070));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11068));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11067));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217840 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11066));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11081));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10901),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11065));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11064));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11063));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11079));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11039),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11062));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11061));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11060));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10967),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11059));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11058));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11057));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11056));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2078),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11055));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11054));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11053));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2092),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11052));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11038),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11077));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10971),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11051));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11050));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10940),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11049));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11076));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11048));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217863 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10897),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_500),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11075));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11047));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11046));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11074));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10975),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11045));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_340),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11044));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217869 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11043));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_500),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11042));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_732),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11041));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11073));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217873 (.A(n_13849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10862),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2095));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11071));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2094));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11069));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11038));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11036));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11033));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11031));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11029));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11027));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11026));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11024));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11023));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11021));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11019));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11017));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11015));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11014));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11012));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11011));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217905 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11006));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11005));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11000));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10998));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10997));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10994));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10992));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10990));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10988));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10986));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217923 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10984));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10982));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10981));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11040));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10980));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217928 (.A(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10979));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11039));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11037));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10978));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_90),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11035));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11034));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11032));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11030));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11028));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2093));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11025));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2092));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2091));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2090));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11022));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2089));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11020));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11018));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2088));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2087));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11016));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2086));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2085));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11013));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2084));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11010));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2083));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11008));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11007));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2082));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2081));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11004));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11003));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10977));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11001));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2080));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10999));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2079));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10976));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10996));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10995));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10993));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10991));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10989));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10987));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10985));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g217975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10983));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10975));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10971));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10969));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10967));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10965));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10963));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10961));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10959));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10956));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10955));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g217991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10954));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10952));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10951));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g217998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10949));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10947));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10946));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10943));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10940));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10936));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218012 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10560),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10878),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10935));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10934));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218014 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10933));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10881),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10932));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218016 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10881),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10931));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_449),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10930));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218018 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10859),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10929));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218019 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10822),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10928));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218020 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10818),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10857),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10927));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10879),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10926));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10925));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10924));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10923));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10922));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10921));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10920));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10974));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10973));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10972));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10970));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10968));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10966));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2078));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10964));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10962));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2077));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2076));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2075));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10960));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10958));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10957));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2074));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10953));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2073));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2072));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10950));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2071));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2070));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10948));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2069));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2068));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2067));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2066));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10945));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10944));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10942));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2065));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10941));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2064));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10939));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10938));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10937));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10918));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10915));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10912));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10910));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10908));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10906));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10904));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10901));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10899));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10897));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218075 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10736),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10919));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10917));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218077 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10784),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10916));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218078 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10718),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10914));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10913));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218080 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10780),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10911));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218081 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10747),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10909));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218082 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10907));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10905));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218084 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_334),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10903));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218085 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10708),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10902));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218086 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10900));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10898));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10895));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2061));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10893));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10891));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218097 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10820),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10890));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218099 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10888));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218100 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10783),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10887));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218101 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10821),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10886));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218102 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10826),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10885));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10884));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10883));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218105 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2015),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10896));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218106 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10882));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2063));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2062));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218109 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10653),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10894));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218110 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_231),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10892));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10881));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2060));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218115 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10880));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10879));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10878));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218118 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10877));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218119 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10786),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10876));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218120 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10875));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218121 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10874));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218122 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10748),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10873));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218123 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10872));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10871));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218125 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10359),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_449),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10805),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10870));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218126 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10806),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10869));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218127 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10868));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218128 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10814),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_238));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218129 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10867));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218130 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10866));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218131 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10865));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218132 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10864));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .A2(n_14469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10863));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10862));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10819),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10861));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10860));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10859));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10858));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10857));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10809),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10856));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218141 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10769),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10855));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218142 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10809),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10854));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10852));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218144 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10337),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10663),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10850));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_449),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10767),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10849));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218146 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10785),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10848));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218147 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10847));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218148 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10351),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10754),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10788),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10846));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218149 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10749),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10353),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10845));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218150 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10746),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10844));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218151 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10778),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10843));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218152 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10842));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218153 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_336),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10841));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218154 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10734),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10840));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218155 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_335),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10839));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218156 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10710),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10838));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218158 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10836));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218159 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10587),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10853));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10851));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10835));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10754),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10834));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10833));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10799),
    .C(u6_n_87),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10832));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218165 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_337),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10831));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10830));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218167 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10829));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10763),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10828));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10827));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10826));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10825));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10824));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10823));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10822));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10821));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10820));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10819));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10818));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10816));
 INVx3_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10814));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10656),
    .B(u6_n_87),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10813));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10812));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10811));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2027),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10810));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .B(u6_n_87),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10817));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10815));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10808));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10806));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10805));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10804));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10411),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10803));
 AOI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10764),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10589),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10809));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218194 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10807));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10802),
    .Y(u6_n_87));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10799));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218197 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10738),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10593),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10798));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10797));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218200 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10481),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2032),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10796));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10795));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10794));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218203 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2022),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10764),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10793));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218204 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2056),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10792));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218205 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10791));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218206 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1997),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10790));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218207 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10690),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10802));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10800));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10788));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10787));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10786));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2059),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10785));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2056),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10784));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10783));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10782));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10758),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10781));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10780));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10779));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10778));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218220 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10756),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2037),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10789));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10776));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10775));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10774));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10773));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10772));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10777));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10729),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10682),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10768));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10767));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10733),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10766));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2054),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10765));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10738),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10771));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10739),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10770));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10769));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10763));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10762));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10740),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10761));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10760));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10459),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10759));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218247 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10723),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10758));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218248 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10398),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10757));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10756));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10605),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2059));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10721),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10764));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218252 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10722),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2058));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218253 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2057));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218254 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2056));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10754));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10753));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10752));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10751));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10716),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10750));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10749));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10748));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10747));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10746));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10745));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10744));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218266 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2025),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10743));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218267 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10416),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10742));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218268 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10741));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218269 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10693),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10755));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2055));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2054));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218274 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10740));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10738));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218276 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10702),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10739));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218277 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10737));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10736));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10735));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10734));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218281 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10666),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2052),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10733));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218283 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2006),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2035),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10729));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218284 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2015),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2017),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10551),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10728));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10494),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10547),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10727));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218286 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2016),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2050),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10726));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10700),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10725));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218288 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2050),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10732));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218289 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10699),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10731));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218290 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2050),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2053));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218291 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10700),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2046),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10730));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10721));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218293 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10683),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10649),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10703),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10720));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10719));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2050),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10718));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218297 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10650),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10717));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218298 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10699),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10716));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218299 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2038),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10724));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218300 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10701),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10723));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218301 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10722));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218304 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2029),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10478),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10715));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10714));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_333),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10713));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218307 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2045),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10490),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10479),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2052));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10695),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10712));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218309 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10420),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10711));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218310 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10446),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2044),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10488),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10477),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2051));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10710));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10709));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10708));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10688),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10707));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10706));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10705));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218319 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2030),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10582),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10704));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218320 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1998),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10425),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10703));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2050));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218324 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10702));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10700));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10701));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10699));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10698));
 AOI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2041),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_10559),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10602),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10637),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10697));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10696));
 NOR4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218334 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10616),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10603),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10693));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218335 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2007),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10557),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10692));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218336 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10691));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10651),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10690));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10555),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10689));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218339 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10404),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10688));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218340 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10399),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10687));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218341 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10559),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2041),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10695));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10694));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10686));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10684));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2041),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10681));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10680));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10679));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10609),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10678));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218352 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10608),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10677));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218353 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2041),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10676));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10611),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10685));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10636),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2049));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10632),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10683));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2048));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218358 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10627),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10682));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10675));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10672));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10671));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10670));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2042),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10669));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10668));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218365 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2028),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10587),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10674));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2023),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10673));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10667));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10663));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218371 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10418),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10549),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10662));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10589),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10449),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10661));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10586),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2015),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10666));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218374 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10665));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10658));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10654));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10652));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10648));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10647));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218383 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2039),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10646));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10645));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2038),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2047));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218386 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10463),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2046));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10660));
 AND4x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10476),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10472),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10659));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10644));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10643));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10642));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10657));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10641));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218394 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10339),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10656));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10640));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10655));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218397 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10383),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10653));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10617),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10639));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10651));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10447),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10650));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10605),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10649));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2032),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10486),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2045));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10631));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10629));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10626));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218415 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2008),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10408),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10624));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2018),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10623));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10436),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10622));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10464),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10621));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218419 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2002),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10620));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10397),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10619));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218421 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2011),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10618));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218422 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10638));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218423 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1999),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10637));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218424 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10474),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10636));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218425 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2033),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2044));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218426 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10367),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2043));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218427 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10450),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10454),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10635));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218428 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10392),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10634));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218429 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10401),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10633));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218430 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2004),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10632));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218431 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2009),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10630));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218432 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10628));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10627));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218434 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10340),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2042));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218435 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1996),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10374),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10625));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218436 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10340),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10372),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2041));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10617));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10615));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10613));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10607));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10604));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10594));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10592));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10590));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10589));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10586));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10585));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10584));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10616));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10583));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10614));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10582));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10581));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10612));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10580));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10611));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2040));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10610));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218466 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10609));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218467 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10608));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10579));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2039));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2000),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10606));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10417),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10605));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10603));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2038));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_196),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10602));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10578));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10577));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218477 (.A(u6_rem_96_22_Y_u6_div_90_17_n_677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10601));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10600));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218479 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10599));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10576));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218481 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10598));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10597));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10596));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10595));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218485 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10575));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10574));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10573));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218488 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10359),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2440),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10572));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10571));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10593));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10570));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10591));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10569));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10568));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10567));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10566));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10471),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10565));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10564));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218499 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10563));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10562));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10561));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2037));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10588));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10587));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10558));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10552));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10550));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10548));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10546));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218513 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10545));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10325),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10544));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218515 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10543));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218516 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10542));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218517 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10541));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10540));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10539));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10538));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10435),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10537));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10536));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10535));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10426),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10534));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10533));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218526 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10532));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218527 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10531));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10530));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10560));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2014),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10529));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10423),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10528));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10428),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10527));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10526));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218534 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10525));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218535 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10524));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218536 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10523));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10559));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10522));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218539 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_35),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10521));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10557));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10556));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2011),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10520));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2036));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10555));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10554));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10519));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10518));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10517));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10516));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10553));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10514));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218553 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10513));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218554 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_732),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10337),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10512));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218555 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10511));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10510));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10509));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10508));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10551));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2035));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10549));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10547));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10506));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10503));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10500));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10495));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10493));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10491));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218570 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10489));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10487));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10485));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10483));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10482));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10481));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10480));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10475));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10473));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10471));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10470));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10468));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10467));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10465));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10463));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10462));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10461));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2021));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10458));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10456));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10455));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10452));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10451));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10448));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10445));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10443));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10441));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10440));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10507));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10505));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10504));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_90),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10502));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10439));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10501));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10499));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10498));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10438));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10497));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2034));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10496));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10437));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10494));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10492));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10490));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10488));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10486));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10484));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2033));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2032));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2031));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10436));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10479));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10478));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10477));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10476));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2030));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10474));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2029));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10472));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2028));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10469));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2027));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2026));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10466));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2025));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2024));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_90),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10464));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2023));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10460));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2022));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2020));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2019));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10459));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_61),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2018));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10457));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2017));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10454));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10453));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2016));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10450));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10449));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10447));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2015));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10446));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10444));
 AND3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218676 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10271),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10442));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10435));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10433));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10431));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10429));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10428));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10426));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10424));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10423));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10421));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10419));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10418));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10416));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10415));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10412));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10411));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10409));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10408));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10403));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10402));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10400));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10398));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10396));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10394));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1998));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10389));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10387));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10385));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218724 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10384));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218725 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10383));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218726 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10382));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10381));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_35),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10380));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2014));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10434));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10379));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10432));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10378));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10377));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10376));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10430));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10375));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10374));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10373));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218740 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10372));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10371));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2013));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10427));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10425));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2012));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10422));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10420));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2011));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2010));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2009));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2008));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2007));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2006));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10370));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10417));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2005));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2004));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10369));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10414));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10413));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10368));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10367));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2003));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10410));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2002));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10407));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10406));
 NAND2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10405));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10404));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2001));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10401));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10399));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2000));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10397));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1999));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10395));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10393));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10392));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10391));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1997));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10390));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10388));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10386));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10365));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10363));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10361));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10359));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10357));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10355));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10353));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10351));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10349));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10347));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10345));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10343));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10341));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10226),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10366));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10364));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10362));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10360));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10358));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10223),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10356));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10354));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10352));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10153),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10350));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10175),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10348));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10346));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10203),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10344));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10342));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10339));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10337));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10335));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10333));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10331));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10329));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10327));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10015),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10259),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10326));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10279),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10325));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218821 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10324));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10323));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10280),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10322));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10281),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10321));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1996));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10340));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218827 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10338));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10275),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10336));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218829 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10127),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10334));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10332));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218831 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10042),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10330));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218832 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10130),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10328));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10319));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10240),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10318));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10317));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218836 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_420),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10316));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10315));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10314));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10313));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218840 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10312));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218841 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10311));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10310));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10309));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218844 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10320));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10308));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218846 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10307));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218847 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10285),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10306));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218848 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10305));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218849 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10304));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218850 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10303));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218851 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10302));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218852 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10301));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218853 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10046),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10300));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10299));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10298));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218856 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10255),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10297));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218857 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_329),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10296));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218858 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9821),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_471),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10295));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_471),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10225),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10294));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10190),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_471),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10293));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9754),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10217),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10248),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10292));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218862 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10208),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_468),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10291));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218863 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9935),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10222),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10290));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10205),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10289));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10209),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10288));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218866 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10129),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10287));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218867 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_331),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_472),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10286));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218868 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10176),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9743),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10285));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218869 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_327),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10284));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10156),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10283));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_326),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10282));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10242),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10281));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218873 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10243),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10280));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218874 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10250),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10279));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10277));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218877 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10217),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10045),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10276));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218878 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .A2(n_14473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10275));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218879 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9972),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_473),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9724),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10274));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218880 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10026),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10246),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10273));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218881 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10100),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10247),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10272));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218882 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10244),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10271));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218883 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10215),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10270));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10269));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218885 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10072),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10268));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218886 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10039),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10267));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218887 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10135),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10266));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218888 (.A1(n_14472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10265));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10264));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218890 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10263));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10262));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10261));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10260));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10259));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10257));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10258));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10255));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10249),
    .B(u6_n_89),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10256));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10254));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10253));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218901 (.A(u6_n_89),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10251));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10248));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9944),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10199),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1972),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10247));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9846),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10246));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10027),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10245));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218906 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9832),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9857),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10244));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218907 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10160),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10224),
    .Y(u6_n_89));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218908 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10102),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10250));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10249));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10241));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10240));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10239));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218913 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10000),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10220),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9999),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10238));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218914 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10219),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1966),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10237));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218915 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1982),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10243));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218916 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1983),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10242));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10236));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10235));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10234));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218920 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10123),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1988),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10182),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10110),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10233));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218921 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10232));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218922 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10231));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218923 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9795),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10230));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218924 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10229));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10228));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10227));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10199),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10226));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218928 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10225));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218929 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10064),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10224));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10191),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10223));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10222));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10221));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10219));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10217));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10216));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9947),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10215));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10214));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9829),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10213));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218939 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9826),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10212));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218940 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10211));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10210));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10178),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10220));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10133),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10157),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10218));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10209));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10208));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10207));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10206));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10205));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10204));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10203));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10202));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10201));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10199));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10198));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10195));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10194));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218957 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1952),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10191));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218958 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_324),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10200));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218959 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10099),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10197));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218960 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1991),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1986),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10196));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218961 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10065),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10193));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218962 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10192));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1992),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10190));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218964 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9948),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10159),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9949),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10189));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218965 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10188));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10187));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10186));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218968 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9783),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10185));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218969 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1963),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10184));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10183));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218974 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10182));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218975 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1971),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10058),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10181));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218976 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1969),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10106),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1970),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10060),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10180));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218977 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1955),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10179));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10178));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1935),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10177));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218980 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9963),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1995));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9970),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1994));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218982 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1976),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1993));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10176));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10175));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10174));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218990 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9851),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10173));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218991 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1942),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10172));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g218992 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10171));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218993 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1959),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10170));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218995 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9921),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10166));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10165));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g218997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10164));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218998 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10085),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9847),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9939),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10169));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g218999 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1948),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10078),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9858),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9943),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10168));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1992));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10162));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10159));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1990));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1991));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10158));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10156));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10155));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10154));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10153));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219014 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10056),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10161));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10054),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10160));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219016 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10055),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10157));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10150));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10025),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10147));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219023 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9834),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10145));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219024 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10121),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10144));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219025 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9960),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10152));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219026 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10151));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219027 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10149));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219028 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10148));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219031 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1987),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10113),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10142));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219032 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10080),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10114),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10141));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219033 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10111),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10140));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219034 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10084),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10139));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10138));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219037 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9967),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10143));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219038 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1989));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219039 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10137));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10136));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10135));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10109),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10134));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1986),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10035),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10092),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_10094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10133));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219044 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9779),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10132));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219045 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9776),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10096),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10131));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10130));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10129));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10128));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10127));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219053 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10082),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1988));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219054 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1944),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10126));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10125));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10123));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10121));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10120));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10117));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10115));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219062 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1961),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10114));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219063 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9827),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9859),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10113));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219064 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1974),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10124));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10093),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10122));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219066 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10013),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10119));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219067 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10118));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219068 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10011),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10116));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10112));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10109));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10107));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219072 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10044),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10105));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1980),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_10019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10104));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219074 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1967),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10111));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10060),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1969),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10103));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219076 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1980),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10110));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10058),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1973),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10108));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219078 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1972),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1982),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10106));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10102));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10099));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10094));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10093));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10092));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1966),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10101));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10091));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10063),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10100));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10090));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10089));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10088));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10049),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10087));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10098));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219095 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9954),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10097));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219096 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1977),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10096));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219097 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9983),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10095));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10086));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10083));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10081));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10079));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219103 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9984),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10077));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219104 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10076));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219105 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9996),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10075));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219106 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9991),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9965),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10074));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219107 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10073));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10072));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10071));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219110 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1951),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10085));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219111 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1940),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10070));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219112 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9995),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10084));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219113 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10001),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9977),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1987));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219114 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9787),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9982),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10069));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219115 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10003),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10082));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219116 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9988),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10080));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219117 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1957),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_10020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10078));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219118 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1978),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10068));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10067));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10063));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219126 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10059));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10057));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1981));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219133 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10056));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10055));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10054));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10066));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10065));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1986));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1985));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10064));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10062));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10061));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219143 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9935),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1984));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10060));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10058));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1983));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1982));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10053));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10051));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10047));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10046));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219153 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9920),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9774),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9919),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10045));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10044));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10043));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219156 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9913),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9774),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9914),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10042));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219157 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9867),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10041));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9918),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10040));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10039));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10038));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10037));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10052));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10050));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10029),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10036));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10049));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10048));
 AOI221x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219167 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9769),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_466),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1980));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10032));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10028));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10025));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10023));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10021));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10018));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10016));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10014));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10013));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10012));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10011));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10035));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10010));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9937),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10009));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9848),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10033));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10031));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10008));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10007));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10030));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10029));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9966),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1979));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10006));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10005));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9951),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10027));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10004));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1975),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10026));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10024));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10022));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10020));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10003));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9768),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10019));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10017));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219203 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9699),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10015));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10000));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9997));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9992));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9990));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9987));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9982));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9981));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219217 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1934),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9980));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219218 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9766),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9979));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219219 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9278),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9978));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219220 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9845),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9977));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219221 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9976));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219222 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9849),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9975));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219223 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9862),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9974));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219224 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9798),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9973));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219225 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1930),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9972));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219226 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9835),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10001));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1967),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9999));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1976),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9865),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9998));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219229 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9793),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1941),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9996));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9822),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9971));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1949),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9995));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9970),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9863),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9994));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9794),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9993));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9991));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1947),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9989));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9988));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1960),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9986));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219238 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9985));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219239 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9791),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9984));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219240 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1930),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9983));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219241 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1930),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1978));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219242 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1931),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1977));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9967));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9963));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9958));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9956));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9953));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9951));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9949));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9947));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9944));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9942));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9941));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9940));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9938));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9937));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9935));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219267 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9934));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9970));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9933));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9969));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9968));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219272 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9966));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9965));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9964));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1942),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9962));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1935),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9961));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9960));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9959));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9957));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9955));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1976));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9954));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9932));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9931));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9930));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9952));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219287 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9929));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9928));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9927));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9926));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9950));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9875),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9925));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1975));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1951),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9948));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9946));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9924));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9923));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9945));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9943));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1974));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1973));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1972));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9939));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1971));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1970));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1969));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1968));
 AO221x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9670),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9669),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9936));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9920));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9918));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9916));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9914));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9912));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219317 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9910));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9909));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219321 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9698),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9618),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9192),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_9697),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9906));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219322 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9700),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_9618),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_9275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9905));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219323 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9904));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219324 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9903));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219325 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9902));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219326 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9901));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_18),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9900));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9899));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9898));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9921));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219331 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_732),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9734),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9919));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9897));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9896));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219334 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9895));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9894));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9893));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9802),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9892));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9891));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9890));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9889));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9888));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9778),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9887));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9806),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9886));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9885));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9884));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219347 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9883));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9815),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9882));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9881));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9880));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9879));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9917));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9878));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9877));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9915));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9734),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9876));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9913));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1967));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9911));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1966));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1965));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9908));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9873));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9871));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9868));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9866));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9860));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9857));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9856));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219374 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9853));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9852));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9851));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9848));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9846));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9844));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1956));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9843));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9842));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9839));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9837));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9836));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9834));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9833));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9832));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9830));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9828));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9826));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9824));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9822));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9820));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_18),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9819));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9818));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9875));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1964));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9874));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9817));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9872));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9816));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_61),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9870));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9869));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1963));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9867));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9865));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_18),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9864));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9863));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9862));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9861));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9859));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1962));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9858));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9855));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1961));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9854));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1960));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1959));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1958));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_90),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9850));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9849));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9847));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9845));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1957));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1955));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_21),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1954));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1953));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9841));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1952));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9840));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9838));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1951));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9835));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1950));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1949));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1948));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9831));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9829));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9827));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9825));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219457 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9654),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9823));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9821));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9815));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9813));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9810));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9808));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9806));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9804));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9802));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9801));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9795));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9792));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219479 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9790));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219481 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9789));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9787));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9786));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9784));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9782));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9781));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9779));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9778));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9776));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9773));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9771));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9770));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9769));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219503 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9710),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9768));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219505 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9766));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219506 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9765));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9764));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9814));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9812));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9811));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9763));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9762));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9761));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219514 (.A(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9809));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9760));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9807));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9805));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_196),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9803));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9759));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1947));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1946));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9799));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_196),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9798));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9797));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9796));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1945));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9794));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9793));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1944));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1943));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9791));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1942));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1941));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1940));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9788));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1939));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1938));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1937));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9785));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1936));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9783));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1935));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1934));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9780));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_18),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1933));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9777));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1932));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9775));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9774));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9772));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9757));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9754));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9752));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9750));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9748));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9746));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9743));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9740));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219559 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9758));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219560 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9616),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9756));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219561 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9634),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9755));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219562 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9631),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9753));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219563 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9751));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219564 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9635),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9749));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219565 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9747));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219566 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9575),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9745));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9744));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9742));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219569 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9561),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9741));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219570 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9739));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9734));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9732));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9731));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9693),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9730));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9729));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9728));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219581 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9681),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9727));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219582 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9726));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1931));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1930));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9531),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9737));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9736));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219587 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9735));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9733));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9724));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219590 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9199),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9655),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9723));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9722));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219592 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9721));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219593 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9652),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9195),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9720));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219594 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9719));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219595 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9718));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219596 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9717));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9716));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219598 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9715));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219599 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9714));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219600 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9664),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9713));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219601 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9223),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9712));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219602 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9711));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219603 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9725));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9710));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219605 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9709));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219606 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9708));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219607 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9707));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219608 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9706));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219609 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9705));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219610 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9704));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219611 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9703));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9702));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9701));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9700));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9699));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9698));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9697));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219618 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9696));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219619 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9587),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9695));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219620 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1905),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9502),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9694));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219621 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9316),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1928),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1901),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9693));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9426),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9692));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9691));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9615),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9690));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219625 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9632),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9689));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219626 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9186),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9688));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219627 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9601),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9687));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219628 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9686));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219629 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9180),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9685));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219630 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9684));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219631 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9683));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9681));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219634 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9557),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9680));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219635 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9679));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9678));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9677));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9676));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219639 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9640),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9642),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9675));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9674));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9673));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9672));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219643 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9159),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9493),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9671));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9670));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9669));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9559),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9668));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9666));
 INVx5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9662));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9660));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1929),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1887),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9659));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9628),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9658));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9231),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9657));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9289),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9656));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219654 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9622),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9667));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1927),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9665));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219656 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1916),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1928),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9664));
 OR2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9663));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9620),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9661));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219659 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9388),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9623),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9387),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9655));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9654));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9653));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9652));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9651));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9650));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9649));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219666 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1927),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9424),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9648));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219667 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9228),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9647));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9645),
    .Y(u6_n_91));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9643));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9420),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9642));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9641));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9421),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9640));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219673 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9609),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9639));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219674 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9638));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219675 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9637));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219676 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9543),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9645));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219677 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9644));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9636));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9635));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9634));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9633));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9632));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9605),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9631));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9630));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9629));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9626));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1927));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219692 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9590),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9625));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219693 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9624));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219694 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9417),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1929));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219695 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9592),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1910),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9628));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219696 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9441),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9627));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219697 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9591),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1922),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1928));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219698 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9590),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1926));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9622));
 BUFx6f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9621));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9618));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9619));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219706 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9580),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9532),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9617));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9616));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9615));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9614));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219710 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9579),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9382),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9613));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219711 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1879),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9612));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219712 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9623));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219713 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9544),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9620));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9611));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219716 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9583),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9608));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219717 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9306),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9607));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219718 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9606));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219719 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9605));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219720 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9260),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9604));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219721 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9299),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9603));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219722 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1925));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219723 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9610));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219724 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9437),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9609));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9602));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9601));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9600));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9599));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9598));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9597));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9570),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9596));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9594));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219735 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9521),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9552),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9595));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219736 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9568),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9593));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9591));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219738 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9522),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9592));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9589));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219740 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9550),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9590));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9588));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9587));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9586));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9583));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9224),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1861),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9379),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9580));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9415),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9579));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9549),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9578));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1921),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9585));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219753 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9551),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9584));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219754 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9435),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1924));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9582));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219756 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9551),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1923));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219757 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9486),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9581));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219758 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9533),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9477),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9577));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9576));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9575));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9536),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9574));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219762 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9573));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219764 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9551),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1891),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9572));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1921),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9571));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219766 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9570));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9569));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219769 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9567));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219770 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1884),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9464),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9311),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1902),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9566));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219771 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9283),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9313),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9317),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9565));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9525),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9564));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9250),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1918),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9563));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9295),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1922));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219775 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1887),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1892),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9307),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9568));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1918),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9562));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9541),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9561));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9560));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9559));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9558));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9557));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219782 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9237),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9556));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219783 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1919),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9555));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9554));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9553));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9552));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1912),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9488),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9551));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1921));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9461),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9445),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_9432),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9466),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9445),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9550));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9549));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9548));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9547));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9473),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9546));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9471),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9545));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9452),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9417),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_9509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9544));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9504),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9543));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9542));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219804 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1912),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9541));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1863),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9540));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1913),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1920));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9432),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1919));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9431),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1918));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9539));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9537));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9534));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9531));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9530));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9529));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9528));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219816 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9444),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9527));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9475),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9526));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9538));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9536));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9470),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9535));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219821 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9436),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9533));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9494),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_872),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9532));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9525));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9522));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9521));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9450),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9520));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9510),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9519));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9378),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9524));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9523));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9518));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9516));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219833 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9380),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9221),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9381),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9514));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9513));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9385),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9222),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9221),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9512));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9511));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9416),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9517));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1862),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1917));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1901),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9515));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9510));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9506));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9503));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9501));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9498));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9497));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9495));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219849 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9175),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9493));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9492));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9491));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9281),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9509));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9490));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219854 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9215),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9489));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9488));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9434),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9507));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9505));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1905),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1916));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9487));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9486));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9504));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219862 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9276),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9275),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9485));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9429),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9484));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9502));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9483));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9482));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9481));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9500));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9499));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1882),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1872),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9496));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9452),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9480));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1860),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9163),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9494));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9476));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9474));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9472));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9468));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9465));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9463));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9460));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219887 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1895),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9459));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1894),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9458));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219889 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9246),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9457));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219890 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9257),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9456));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219891 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9236),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9455));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219892 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9286),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9454));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219893 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9453));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219894 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9288),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9479));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9478));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9409),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9477));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219897 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9475));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219898 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1880),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9473));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219899 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1904),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9471));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219900 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9245),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1878),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9470));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9469));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219902 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1869),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9467));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9466));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1899),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1915));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1888),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1914));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219906 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1898),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9464));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219907 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1907),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9462));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219908 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9205),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9461));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219909 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9175),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1913));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219910 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9176),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1912));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9450));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9447));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9443));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9441));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9439));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9435));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9431));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9429));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9427));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9424));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219923 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9421));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9419));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9415));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9412));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9452));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219928 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9410));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9409));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9408));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9407));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9451));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219933 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9449));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9298),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9448));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1911));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9446));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9445));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1875),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9444));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9442));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1879),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9440));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9438));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9437));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g219943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9436));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9434));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9433));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9432));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9430));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9406));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1910));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9428));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1897),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9426));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9405));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9425));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9423));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9422));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1905),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9420));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9404));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219958 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_565),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9403));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9402));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9401));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1907),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9400));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9399));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9398));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9397));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1903),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9395));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9394));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9418));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9393));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9392));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9391));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9417));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9276),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9416));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9414));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9413));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9411));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9390));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9388));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9386));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9384));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9381));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9377));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9376));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9375));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g219985 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9374));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219986 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9373));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9372));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9371));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219989 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9370));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9285),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9369));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9368));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9367));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219993 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9366));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9365));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9364));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9389));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9387));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9363));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g219999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9362));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9361));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220001 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9360));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_732),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9385));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9383));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9359));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220005 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_131),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_836),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9358));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1880),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9357));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1898),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9356));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220008 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9355));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220009 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9180),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9354));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9353));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9352));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9351));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9350));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220014 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9349));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220015 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9348));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1881),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9347));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9346));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9345));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9344));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9343));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9342));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9382));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9341));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9340));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9339));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9338));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220027 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9337));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220028 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9380));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220029 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9336));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9379));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9378));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9335));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9331));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9327));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9324));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9323));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9321));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9319));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9318));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9316));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9315));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9314));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9313),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9312));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9310));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9308));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9306));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9305));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9302));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9301));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9300));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9297));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9295));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9293));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9291));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9289));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9287));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9285));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9284));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9282));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9280));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9279));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9278));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9277));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9275));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9334));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9274));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9333));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9332));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1909));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9330));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9329));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9328));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9273));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9272));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9326));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_61),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9325));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9271));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1908));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1907));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9322));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9320));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1906));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9317));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9199),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1905));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1904));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1903));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1902));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1901));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9313));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9311));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1900));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1899));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9309));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220125 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9307));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220126 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9304));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220127 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1898));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9303));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220129 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1897));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9270));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1896));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9299));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220133 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1895));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9298));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1894));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9296));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9294));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9292));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9290));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1893));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9288));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1892));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9286));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1891));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1890));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1889));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1888));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9283));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1887));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9281));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1886));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1885));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1884));
 AOI211x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220154 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9094),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9115),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1883));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9276));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9268));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9266));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9264));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9262));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9260));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9259));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9256));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9254));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9253));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9252));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9250));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9248));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9247));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9243));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9241));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9239));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9237));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9234));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9233));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1865));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9230));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9229));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9226));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9223));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9221));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9220));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9219));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9216));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9215));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220210 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9214));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220211 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9159),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9213));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220212 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9138),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9212));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9211));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9269));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9210));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9209));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1882));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_18),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9208));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9267));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1881));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9265));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9207));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9206));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9205));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9204));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9203));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9263));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1880));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9261));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9258));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9257));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1879));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9255));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1878));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1877));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1876));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220237 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9251));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1875));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9249));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1874));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1873));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1872));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9246));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1871));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9245));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9244));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9242));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9240));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9238));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1870));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9236));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9235));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1869));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1868));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1867));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1866));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9231));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1864));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_30),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1863));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1862));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1861));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9228));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9227));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9225));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9224));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9222));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9218));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9217));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9201));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9199));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9197));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220272 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9194));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9192));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9190));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9188));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9186));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9184));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9182));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9180));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9178));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220281 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9051),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9202));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9200));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9198));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9157),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9196));
 AND3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9113),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_9132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9195));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220286 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9193));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9070),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9191));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9189));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9187));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220290 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8983),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9185));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220291 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9017),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9183));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220292 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9050),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9181));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220293 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8996),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9179));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9177));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9174));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9172));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9168));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9165));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9164));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9163));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220301 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9162));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9161));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220303 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9100),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9160));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9176));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9175));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8967),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9173));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9171));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8822),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9170));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9169));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9167));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220311 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9166));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9158));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220313 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9157));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220314 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9046),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9156));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220315 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1860),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9089),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9155));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220316 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9154));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9153));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220318 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9152));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220319 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9062),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9151));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220320 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9093),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9150));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220321 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9149));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220322 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9148));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220323 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9159));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220324 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9147));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220325 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9146));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220326 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9145));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9144));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220328 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8965),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9143));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9142));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9141));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220331 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9140));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220332 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9139));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9096),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9138));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9137));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220335 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8589),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9136));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220336 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9135));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220337 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8595),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9134));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8593),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9133));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220339 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1860),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9081),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8592),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9132));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220340 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8751),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9131));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220341 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8669),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9130));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220342 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1859),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8588),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9129));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1859),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9014),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9128));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220344 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9127));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220345 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9126));
 AOI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220346 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9058),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_9048),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9125));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220347 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8995),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9124));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1859),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8966),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9123));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220349 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8963),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9122));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8753),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9084),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9120));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220352 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8780),
    .A2(n_14474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9119));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220353 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9041),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9118));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9117));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9116));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220356 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9115));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9114));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9082),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9113));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9112));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9111));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9025),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9024),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9110));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220362 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8924),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9109));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9108));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9107));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9106));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9105));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220367 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8883),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9104));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8855),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9103));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8823),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8560),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9102));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220370 (.A(n_14474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9101));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9084),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9100));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220372_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_413));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9099));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220374 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9097));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220375 (.A(u6_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9098));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9080),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9096));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9095));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9094));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9093));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9074),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9092));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9091));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9090));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220383 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9076),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9089));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9087),
    .Y(u6_n_93));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8975),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9071),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9087));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9002),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9086));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220389 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8893),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9084));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9056),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8769),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9083));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9082));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9054),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9081));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220393 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9038),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8970),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9079));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9078));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220395 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9077));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220396 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1858),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9076));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220397 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9044),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8792),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9075));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220398 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9043),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9074));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9073));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220400 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9072));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220401 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1845),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9080));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8951),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9023),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8897),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9071));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9044),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9070));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220404 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8875),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9043),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8876),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_9042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9069));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9039),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9068));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9067));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9066));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9065));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9064));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9034),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9063));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9062));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9060));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9059));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9061));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1859));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9058));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220421 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8673),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9028),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9056));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220422 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8675),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9055));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220423 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8617),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_9029),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9054));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9053));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220426 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8974),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9057));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9007),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9051));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9050));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9049));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9048));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9047));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9046));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9045));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9042));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9041));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9040));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220440 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1853),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8930),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9044));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220441 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1858));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220442 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9000),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1857));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220443 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8998),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1856));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220444 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8997),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9043));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220445 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8949),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9038));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9037));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220447 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8795),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8998),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8796),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9036));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220448 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8961),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9035));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220449 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9004),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9034));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220450 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_9001),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1819),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9033));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220451 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1821),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9032));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220452 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1854),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9039));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9030));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9027));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220456 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8987),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9026));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9025));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9024));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1841),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8986),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9023));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220460 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8753),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1831),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8894),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9022));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220461 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9021));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220462 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9020));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220463 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_318),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9019));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1851),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9031));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220465 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1850),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9029));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220466 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8812),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9028));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9018));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9017));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9016));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9015));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9014));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9013));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8730),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9012));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220474 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9011));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9010));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1825),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8992),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9009));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1797),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9008));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220478 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1823),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9007));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220480 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8935),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8707),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8790),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1855));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220481 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9006));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8787),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9005));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9004));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1854));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220486 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8901),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9003));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8947),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8950),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9002));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9001));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1853));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9000));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220492 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8999));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8997));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220494 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8957),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8998));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8971),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8996));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8995));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8994));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8992));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1850));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220504 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8957),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8990));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220505 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8989));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220506 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1847),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8993));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220508 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1837),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1852));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220509 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_317),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1851));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220510 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1847),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8991));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220511 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1849));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8835),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8931),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8988));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220513 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8783),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8987));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1846),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8986));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8985));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8984));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8983));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220518 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8845),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8928),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8982));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220519 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8832),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8977),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8981));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220520 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8980));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8910),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8979));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220522 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8674),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8691),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8704),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8978));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220523 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1812),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8705),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8680),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8977));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8618),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8623),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8646),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8976));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8951),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8975));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8942),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1845),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8913),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8974));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220527 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8641),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8973));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220528 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8972));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220529 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8632),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8944),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8971));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220531 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8969));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8887),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8968));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8944),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8967));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8966));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8965));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8964));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8963));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8962));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220539 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8943),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8970));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220540 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1848));
 NAND4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8907),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8909),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8782),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8961));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1847));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220545 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8802),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1836),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8833),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8802),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8959));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220547 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8958));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8956));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220549 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8828),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8807),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_8801),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8840),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8807),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8957));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8955));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220552 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1834),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8905),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1846));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220553 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8907),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8954));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8953));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220555 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8952));
 AND4x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8904),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8781),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8951));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8950));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8894),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8753),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8892),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8949));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8948));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8942));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8947));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8907),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1845));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8941));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8918),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8940));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8939));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8906),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8938));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8905),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8937));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8894),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8936));
 OA21x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8946));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220571 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8945));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220572 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8944));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8943));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8934));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8932));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8930));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8927));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8925));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8924));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220581 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8806),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8923));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220582 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1822),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8935));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220583 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8933));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220584 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8827),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8922));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8921));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220586 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8829),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1802),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8920));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220587 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8804),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8931));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8929));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220589 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8928));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220590 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8809),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8926));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1820),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1844));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8919));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8918));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8916));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8914));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8912));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1841));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8906));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8904));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8903));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8810),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8902));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8901));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8917));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8915));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1843));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8900));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8913));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8911));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8910));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1842));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8909));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8908));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8907));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8905));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8899));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8896));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8892));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220621 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8764),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8620),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8891));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220622 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8758),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8619),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8890));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220623 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8702),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8889));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8888));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8887));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8886));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_872),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8885));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8884));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8761),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8883));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8882));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8898));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8897));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8895));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8881));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8894));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8893));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8880));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8878));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8876));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8874));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8869));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8867));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8865));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8863));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8860));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8858));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8857));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8856));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8879));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8855));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8854));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_838),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8877));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8853));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8783),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8852));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_565),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8851));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8850));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8875));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1834),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8849));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8873));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8872));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8871));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1830),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8848));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8847));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8870));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8846));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8868));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8866));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8864));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8862));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220671 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8861));
 AND3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8566),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8859));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8842));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8839));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8837));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8831));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8829));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8827));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8825));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8655),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8824));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220687 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8823));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220688 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8822));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220689 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8666),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8821));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1806),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8820));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220691 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1799),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8819));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220692 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8608),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8818));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220693 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8682),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8817));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220694 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8693),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1818),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8816));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220695 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1816),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8815));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220696 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8694),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8814));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8845));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220698 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1826),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1840));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220699 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1815),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8844));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220700 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1814),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8690),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8843));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220701 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1824),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8841));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220702 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8648),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8840));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220703 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1839));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220704 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8645),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8838));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220705 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1798),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8836));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8618),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8835));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220707 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8642),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8833));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1812),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8832));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220709 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1838));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220710 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8830));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220711 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8607),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8828));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8826));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8812));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8800));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8798));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8796));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8794));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8792));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8791));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8789));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8787));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8785));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8782));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8780));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8779));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8813));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8811));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8810));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220739 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_528),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8809));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220740 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1837));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220741 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8808));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8807));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8806));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8805));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220745 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8804));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8803));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8802));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8801));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8799));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8778));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8777));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8776));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8642),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1836));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1820),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8797));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8775));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8774));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8795));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8773));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8684),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8772));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8701),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8771));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8770));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8706),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8793));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8769));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8768));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8767));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8685),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8766));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1835));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1834));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1833));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1832));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8790));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8788));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8786));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8667),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8784));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8783));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8781));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8765));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8763));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8761));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8759));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8757));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8754));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8752));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8750));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8749));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8748));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8747));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8746));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8745));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8764));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8744));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8743));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8742));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8762));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_132),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8741));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8740));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220799 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8739));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8738));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8737));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8736));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1815),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8735));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220804 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8734));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8733));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8732));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8731));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2842),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8730));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8729));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8649),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8728));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8727));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8726));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8725));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8724));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8760));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8723));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_745),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8722));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1813),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8721));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8720));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8719));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220821 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8758));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8718));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8717));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8756));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1831));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8755));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1830));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8753));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8751));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8716));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8714));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8712));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8710));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8708));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8706));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8704));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8701));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8700));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8699));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8698));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8697));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8696));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8692));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8688));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8686));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8684));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8681));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8678));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8676));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8674));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8673));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8671));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8669));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8667));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8666));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8715));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1829));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8713));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1828));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8665));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8711));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8664));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8709));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8663));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8662));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8661));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8707));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8705));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1827));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8703));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8702));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1826));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1825));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1824));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1823));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1822));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1821));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1820));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1819));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1818));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1817));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1816));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8695));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8694));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8693));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220905 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8691));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8690));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220907 (.A(u6_rem_96_22_Y_u6_div_90_17_n_119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8689));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1815));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8687));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1814));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1813));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8660));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8685));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8659));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8683));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8682));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8680));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8679));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8677));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8675));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1812));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8672));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220923 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8670));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220924 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8486),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8668));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8658));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8655));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8653));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8651));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8647));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8644));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8643));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8641));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8640));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8639));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8638));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8635));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8632));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8629));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8628));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8627));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8625));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8622));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8621));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8619));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8617));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220961 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8616));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8615));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220963 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8614));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220964 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8613));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220965 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8536),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8612));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8611));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220967 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8610));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220968 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8537),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8545),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8609));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8608));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8657));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8607));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8606));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8656));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8654));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1811));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1810));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8652));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8650));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8605));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8604));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1809));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8649));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1808));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8648));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8646));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8645));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8603));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1807));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1806));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8642));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1805));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1804));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1803));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8637));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8636));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8634));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g220997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1802));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g220998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8633));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g220999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8631));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8630));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1801));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1800));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1799));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8626));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1798));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8624));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8602));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8623));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1797));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8601));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8620));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8618));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8599));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8597));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221015 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8595));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8593));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8591));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8589));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8587));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8585));
 INVx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8583));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8581));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8579));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8577));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8600));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8598));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221027 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8436),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8596));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221028 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8594));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221029 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8466),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8592));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8510),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8590));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8588));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221032 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_309),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8586));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8584));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8582));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8580));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221036 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8578));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1796),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8575));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8573));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8570));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8568));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221043 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8488),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8567));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221044 (.A1(n_14476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8566));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221045 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8565));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221046 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8564));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8563));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_316),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8562));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8561));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221050 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8576));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1796));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8574));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221053 (.A(n_14520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8572));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8571));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221055 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8569));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8560));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8559));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221061 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8558));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221062 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8464),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8557));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221063 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8014),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8483),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8556));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221064 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8555));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221065 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8554));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221066 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8553));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221067 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8552));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221068 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8487),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8551));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221069 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8550));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221070 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8549));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221071 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8405),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8548));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221072 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8547));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221073 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8499),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8546));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221074 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1795));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8545));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221076 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8544));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221077 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8543));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221078 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8542));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221079 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_429),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8541));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8540));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221081 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8539));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221082 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_430),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8417),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8538));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8537));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8536));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8535));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8534));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8533));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8532));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221089 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8531));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221090 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8529));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221091 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8332),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8528));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221092 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8387),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8527));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221093 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8470),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8526));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221094 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8012),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_314),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8525));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221095 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8010),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8524));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221096 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8008),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8452),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8432),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8523));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221098 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_428),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_446),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8521));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221099 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8520));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221100 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8519));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221101 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8518));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221102 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8517));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221104 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8530));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8515));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221106 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8334),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8514));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221107 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .A2(n_14477),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8513));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221108 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8475),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8512));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221109 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8444),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8511));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8510));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8509));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8508));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221113 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8391),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8507));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8506));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8504));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221117 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8317),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7991),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8503));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8471),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8502));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8501));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221120 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8351),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8500));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8496));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221122_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_429));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1794),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8106),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8493));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221125 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8066),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8492));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221126 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1756),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8491));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221127 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1750),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8490));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221128 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8306),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8499));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221129 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8498));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221130 (.A(u6_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8497));
 OR2x6_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221131 (.A(u6_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8495));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8489));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8457),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8243),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_8456),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8488));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8487));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8486));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8485));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8484));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8483));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221140 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8457),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8482));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8479));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8478));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8477));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8476));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1762),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8475));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221146 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8249),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8474));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221147 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1731),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8473));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8472));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221149 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8471));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221150 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8420),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8367),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8449),
    .Y(u6_n_95));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8480));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8470));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8469));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8429),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8468));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8467));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8466));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8465));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8441),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8464));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8463));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221161 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1793),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8462));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8460));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8456));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221166 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8124),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8455));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221167 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1790),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8461));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8233),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8426),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8459));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8252),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8423),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1794));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1791),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8458));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221171 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8325),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8457));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8454));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8451));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221175 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8335),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8357),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8408),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8354),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8450));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221176 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8424),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8449));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8448));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221178 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8427),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8447));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221179 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8427),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8453));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221180 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8368),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8452));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8445));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8444));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8443));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8137),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8442));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8414),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8441));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221189 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8440));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221190 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8439));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8272),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1793));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8267),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1792));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_312),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8446));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8438));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8437));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8436));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8435));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8434));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8402),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8433));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8432));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8431));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221203 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8430));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221204 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8429));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221205 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8347),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8428));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8427));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8426));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8342),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8380),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8425));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221210 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8424));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8423));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8422));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1791));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8421));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221216 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8420));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8419));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1790));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221220 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8344),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8418));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8417));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8416));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8415));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8413));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8412));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8411));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8237),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8410));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1755),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8336),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1774),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8238),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8409));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8209),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8372),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8408));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8262),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8414));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8261),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1789));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1786),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1788));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8376),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1787));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221239 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8361),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8379),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8406));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1786),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8405));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221242 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8297),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8404));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8403));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1786),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8044),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8402));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8376),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8401));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1747),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8400));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221247 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8381),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8407));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8399));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8397));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8111),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8114),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8395));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8394));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8393));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221253 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1757),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8108),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8112),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8392));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8391));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221255 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8106),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1761),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8120),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8398));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221256 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8370),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8390));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221257 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8122),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8396));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8363),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8389));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8388));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8362),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8387));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8386));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221264 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8371),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8385));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221265 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8369),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8384));
 NAND2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8354),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8383));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8382));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8381));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221271 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8282),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8380));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221272 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1731),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1749),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8379));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8378));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1786));
 OAI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221277 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8259),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1780),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1783),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8259),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8377));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8375));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221279 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8376));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221280 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8374));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221281 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8337),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8373));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221282 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8339),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8372));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8368));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8346),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8322),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8367));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1784),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8366));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221288 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8319),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8365));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1777),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8364));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221290 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1740),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8363));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221291 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8362));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221292 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1778),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8371));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221293 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8370));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221294 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1779),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8281),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8369));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8360));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8358));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8356));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8353));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8352));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8351));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221302 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8299),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8350));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221303 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8349));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221304 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8348));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221305 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8294),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8361));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8270),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8359));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221307 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8289),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8357));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8302),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8271),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8355));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221309 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1753),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8354));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8346));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8271),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8344));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8343));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8342));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221314 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8341));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8347));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8238),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1755),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_8126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8345));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221317 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8340));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8338));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8334));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221321 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8339));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221322 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1770),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8337));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221323 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1765),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8336));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8207),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8335));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8329));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8327));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8325));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8323));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8319));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8318));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8317));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221337 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8037),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1729),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8314));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1778),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8313));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8312));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8236),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8311));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8310));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8309));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8332));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8308));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8307));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8306));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8305));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8331));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1785));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8330));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8116),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1750),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8328));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8326));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8122),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8324));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8322));
 NAND3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8103),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8321));
 AOI211x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7970),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8320));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8304));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8301));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8295));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8293));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8291));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8288));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8285),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8286));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8285));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8283));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1782));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8281));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1781));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1732),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8279));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8109),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8278));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8277));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221377 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8048),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8276));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8275));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221379 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1767),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8274));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8061),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8273));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221381 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8043),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8303));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8302));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1764),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1784));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221384 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1762),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8300));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8299));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1739),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8052),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8298));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1741),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1783));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8297));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1731),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_8047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8296));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221390 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1748),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8294));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221391 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8073),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8292));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221392 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1773),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8139),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8290));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221393 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8116),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8289));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221394 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8287));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221395 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8033),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1729),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8032),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8284));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221396 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1728),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8034),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8282));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221397 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1730),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8280));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8269));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8267));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8264));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8261));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8257));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8250));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8248));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8246));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8244));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8242));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8239));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8237));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8235));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8234));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8272));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8271));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8009),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8270));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8268));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8266));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8233));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1772),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8265));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8263));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8262));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8260));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8259));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8258));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8232));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1747),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8256));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8255));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1780));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1779));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8254));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8253));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8252));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8251));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8049),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1778));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221438 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8014),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_559),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8231));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8249));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8230));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8247));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8245));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8229));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8228));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8227));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8226));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8225));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8224));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1777));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221450 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8223));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8222));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8243));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1769),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8221));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1767),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8220));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8219));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221456 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8218));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8241));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8240));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8238));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8236));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8217));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8215));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8209));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221469 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8205));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221470 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8204));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8157),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8203));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8202));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8201));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221474 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8200));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8216));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8199));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221477 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8198));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8197));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221479 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8196));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8195));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8194));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8045),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8214));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8193));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8192));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8046),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8191));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8190));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8189));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8188));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8213));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8187));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8186));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8185));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8184));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8183));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8182));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221496 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_8005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8181));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8180));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8179));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8092),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8178));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8063),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8177));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8062),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8176));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221502 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8175));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1752),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8174));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8173));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8055),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8172));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8085),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8171));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8170));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221508 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8211));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1761),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8169));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221510 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8210));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8168));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8167));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1776));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221514 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8207));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8164));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8161));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8159));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8157));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8155));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8152));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8149));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8148));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8146));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8145));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8143));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8140));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8139));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8137));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8136));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8134));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8132));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8130));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8129));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8128));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8127));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8125));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8124));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8121));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8119));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8118));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8117));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8115));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8113));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8110));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8107));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8105));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1756));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8102));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8101));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8099));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8097));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8096));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8166));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8165));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8163));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8095));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8162));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8094));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1775));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8160));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8158));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8156));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8093));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8154));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8153));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8151));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8150));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1774));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8147));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8144));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8142));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8141));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1773));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8138));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1772));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8135));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8133));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1771));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1770));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8131));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1769));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1768));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1767));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1766));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1765));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8126));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8123));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8122));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8120));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1764));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1763));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1762));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8116));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1761));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1760));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8114));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1759));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8112));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8111));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1758));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8109));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8108));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1757));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8106));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8104));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8103));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1755));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1754));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7987),
    .C(n_14478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1753));
 AND3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7986),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8100));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221638 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7947),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8098));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8092));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8087));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8085));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8083));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8081));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8079));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8077));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8075));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8074));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8071));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8070));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8066));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8063));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8062));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8060));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8058));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8056));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8055));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8053));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8051));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8046));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8045));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8042));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_102),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8039));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221692 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8037));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221693 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_459),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_462),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8036));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8091));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8035));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8034));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8033));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8032));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8090));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8031));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8088));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8086));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8084));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8082));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1752));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8030));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8080));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221708 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8078));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8029));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8076));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1751));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1750));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8073));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8072));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1749));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8069));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8068));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8024),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8067));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8065));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8064));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1748));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1747));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1746));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1745));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8061));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1744));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8059));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8057));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1743));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1742));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1741));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1740));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8054));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8052));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1739));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8049));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1738));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8048));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8047));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221740 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1737));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1736));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1735));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1734));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8044));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8043));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1733));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1732));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8041));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8040));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1731));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8027));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8025));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8023));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8021));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8018));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8016));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8014));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8012));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8010));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8008));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7851),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8028));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221762 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7890),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_305),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8026));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8024));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221764 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7879),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8022));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7849),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8020));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221766 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7878),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8019));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8017));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221768 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7910),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8015));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221769 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8013));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8011));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7978),
    .B(n_14575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8009));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1728));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8005));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8000));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7996));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7994));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221783 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7913),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7993));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7992));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1730));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1729));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8006));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7971),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8004));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8003));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7965),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8001));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7974),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7999));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7998));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7973),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7997));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7995));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7990));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7932),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7989));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7881),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7988));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221798 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_462),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_307),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7987));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7986));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7985));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7915),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7984));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7983));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7982));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221804 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7981));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7911),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7980));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7880),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7979));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_462),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7991));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7819),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7978));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7977));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221810 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7976));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221811 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7975));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221812 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7974));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221813 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7973));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221814 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7834),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7972));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7971));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221816 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7755),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7942),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7970));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7969));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7968));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7967));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7966));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7965));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7912),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7964));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221824 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7622),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7962));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221826 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7760),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7905),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7960));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7959));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_462),
    .Y(u6_n_96));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221829 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7529),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7957));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7956));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7955));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7954));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7953));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7952));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7951));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221836 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7693),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7950));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7949));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7948));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7947));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7945));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7901),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_462),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7627),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7944));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7943));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7942));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_419),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7941));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221846 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7899),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_461),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7455),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7940));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221847 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_419),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7939));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221848 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7938));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221849 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7450),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_461),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7937));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221850 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7448),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7936));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221851 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7882),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_304),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7935));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221852_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_463));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7883),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7921),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7946));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221854 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_416),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7934));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7875),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7933));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7897),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7932));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221857 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_418),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7931));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221858 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7776),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_419),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7930));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_416),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7929));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_418),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7928));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7753),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_416),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7425),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7927));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221862 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1665),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_416),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7926));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7896),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7925));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7924));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7921));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7918));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221869 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7917));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7537),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7923));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7916));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7853),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7806),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7920));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221873 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7894),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7919));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7887),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7915));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7914));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7913));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7912));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7911));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7910));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7908));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7907));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7906));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221884 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7555),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7562),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7905));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7904));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7903));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7828),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7909));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7901));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7900));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7899));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221893 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7869),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7898));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221894 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7897));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221895 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7896));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221896 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7902));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7894));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7892));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221902 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7788),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7839),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7793),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7891));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7673),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7862),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7674),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7890));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1725),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7889));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1693),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7888));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221906 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7887));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221907 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7886));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221908 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1668),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7885));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221909 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1724),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7884));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221910 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7764),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1726));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221911 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7854),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7895));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221912 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7854),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7893));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7882));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7649),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7881));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7880));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7879));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7878));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7877));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7656),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7876));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7875));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221923 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7874));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7873));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221925 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7798),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7883));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221926 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7782),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7872));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221927 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7871));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7836),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7870));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221929 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7869));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7868));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221931 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7836),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7867));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7866));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7862));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221937 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7861));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7476),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7860));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221939 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7540),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7859));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221940 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7482),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7858));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221941 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7822),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7857));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7824),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7856));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7541),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7855));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221944 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7865));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221945 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7682),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7864));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221946 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1725));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221947 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_300),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7863));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7854));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7826),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7852));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7851));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7850));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221953 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7669),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7821),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7668),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7849));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7664),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7830),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7665),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7848));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7847));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7846));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7845));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7823),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7844));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7843));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221960 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7662),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1724));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221961 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7758),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7853));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221963 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7786),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1703),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7542),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1723));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7842));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221965 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1682),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7574),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7579),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7841));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1700),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7729),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7840));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221967 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7722),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7839));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221968 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7807),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7838));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7836));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221970 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1721),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7837));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7698),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7835));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7834));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7833));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7809),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7832));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7829));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7792),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7828));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221978 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7827));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7795),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7826));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221980 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7825));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7737),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7831));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221982 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7830));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221983 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7795),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1722));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7821));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221986 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7820));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221987 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7819));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7818));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221989 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7658),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7824));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g221991 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7823));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221992 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7813),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7822));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7817));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221994 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1667),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1672),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7495),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7815));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221995 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1683),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1694),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1696),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7814));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221997 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7699),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7813));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g221998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7812));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g221999 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1685),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7546),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7545),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7816));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222000 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7811));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222001 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7512),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7810));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7491),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7809));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222003 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7536),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7778),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7807));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7791),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7806));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222005 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1716),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7805));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7804));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7785),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7803));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7802));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7801));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7767),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7800));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7799));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222012 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7777),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7808));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7764),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7683),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7798));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7696),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7797));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7796),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7795));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7719),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7796));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222022 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7697),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1721));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222023 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7794));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222024 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7754),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7793));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7790));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7787));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222031 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7784));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7754),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7783));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7792));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222034 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1686),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1720));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222035 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1697),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1719));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7791));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7729),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7789));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7731),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7537),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7782));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7722),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7788));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222041 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1699),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7786));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222042 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1708),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1718));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222043 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7785));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222044 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1706),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1717));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7780));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7776));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7702),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7775));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222049 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7707),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7774));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222050 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7687),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7773));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222051 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7709),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7772));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1706),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7771));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7770));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222054 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1708),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7769));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222055 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1706),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7768));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222056 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7659),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7781));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222057 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7779));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222058 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7577),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1716));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222059 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1707),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7767));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222060 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7731),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7778));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222061 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7723),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7777));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7766));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7762));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7759));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7758));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7537),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7757));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7756));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7765));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7764));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1715));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7763));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1714));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7761));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7730),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7760));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7475),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7753));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7729),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7752));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7755));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222083 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7751));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7740),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7750));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7749));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7748));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7747));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7746));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222089 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7471),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7623),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_454),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7754));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7744));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7742));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7739));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7737));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7733));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7730));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7728));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7726));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7724));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7719));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7666),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7718));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7717));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222105 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7534),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7716));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7715));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7714));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7745));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7743));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1713));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7741));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7713));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7740));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2438),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7738));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7736));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7735));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7734));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7732));
 AND4x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7543),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7556),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1712));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7731));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7729));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7727));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7725));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2438),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1711));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222125 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7723));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222126 (.A(u6_rem_96_22_Y_u6_div_90_17_n_865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7722));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222127 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7721));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7720));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7710));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7708));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7706));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7703));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7701));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1708));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1706));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7695));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7519),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7522),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7694));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7693));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222148 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7474),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1666),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7692));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222149 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7565),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7691));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222150 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7690));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222151 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7486),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7689));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222152 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7549),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7688));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1701),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7687));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222154 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7686));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222155 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7510),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7685));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222156 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7684));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7712));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222158 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1670),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7711));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222159 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7478),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1710));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1669),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7709));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222161 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7707));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222162 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1690),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1709));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222163 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1688),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7705));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222164 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7556),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7704));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222165 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7489),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7702));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7552),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7559),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1685),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7700));
 AND4x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7534),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1684),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7699));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222168 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7698));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1666),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7697));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1666),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7468),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1707));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222171 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7457),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7696));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7674));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7671));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7669));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7667));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7665));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7663));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1684),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7662));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7661));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7660));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7683));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7682));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7659));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7658));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7657));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7681));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_123),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7680));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7656));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7679));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222194 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7678));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7677));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7676));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7675));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7655));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7673));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7672));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7452),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7654));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7653));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7652));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7651));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7650));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7649));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7670));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1699),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7668));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7648));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7647));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7666));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7646));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7645));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7557),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7644));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7643));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7642));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7641));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7640));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7639));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1688),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7664));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7638));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7637));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7635));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7630));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7628));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7626));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7624));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7623));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7622));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7621));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7620));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7619));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7618));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7617));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222238 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7452),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7616));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7615));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222240 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7614));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7613));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7612));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7611));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7610));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7609));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7608));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222247 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7428),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7636));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7607));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7634));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7606));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7605));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7604));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7603));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7602));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7601));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7600));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222257 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7423),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7599));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7494),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7598));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7597));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7596));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222262 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7595));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222263 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7594));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7593));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222265 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7633));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1690),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7632));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222267 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7592));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7631));
 AND3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7416),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7399),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7629));
 OA211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222270 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7417),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7627));
 AND3x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7420),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7398),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7625));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7590));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7588));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7585));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7583));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7581));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7580));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7578));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7576));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7575));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7572));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7571));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7570));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7569));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7568));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7566));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7562));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7560));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7558));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7557));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7555));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7554));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7552));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7551));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7550));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222317 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7548));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7547));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7544));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7541));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7540));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7538));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7537));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7535));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7532));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7531));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7529));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7528));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1705));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7527));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_92),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7591));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7589));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7587));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7586));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7584));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7526));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1704));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1703));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7582));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1702));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7579));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1701));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7577));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7574));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7525));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7573));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1700));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222356 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1699));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1698));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1697));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7567));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7565));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7564));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1696));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7563));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7561));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1695));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7559));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1694));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7556));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1693));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1692));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7553));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1691));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1690));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222374 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1689));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222375 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7549));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222376 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7546));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7545));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1688));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1687));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7543));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1686));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7542));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222383 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1685));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1684));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1683));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222386 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7539));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7536));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1682));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7534));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7533));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1681));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7530));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7524));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7521));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7519));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7517));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7514));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7512));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7511));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7509));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7508));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7507));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7502));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7495));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7494));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7492));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7488));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7484));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7483));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7481));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7479));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7477));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1667));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222432 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_102),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7474));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7473));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222434 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7472));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7471));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222436 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7470));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_454),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7469));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7468));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7523));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7467));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1680));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7466));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1679));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7522));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7520));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7518));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7465));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7516));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7464));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7515));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7463));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7462));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1678));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1677));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7513));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7510));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1676));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1675));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1674));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7506));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7505));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7503));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7500));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7499));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7461));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7498));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7497));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7496));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1673));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7493));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7491));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7490));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7489));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222474 (.A(u6_rem_96_22_Y_u6_div_90_17_n_189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7487));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7486));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7460));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222477 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7485));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1672));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222479 (.A(u6_rem_96_22_Y_u6_div_90_17_n_796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1671));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7482));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222481 (.A(u6_rem_96_22_Y_u6_div_90_17_n_782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1670));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7480));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222483 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1669));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7478));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7459));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7476));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7475));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1668));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7458));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7455));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7452));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7450));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7448));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7446));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7444));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7442));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7440));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7438));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7436));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7434));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7432));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7457));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222504 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7456));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7454));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222506 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7453));
 NAND3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7369),
    .B(n_14479),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7451));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222508 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7449));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7367),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7447));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7404),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7445));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222511 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7443));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7441));
 AO221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222513 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7283),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7287),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7439));
 AO221x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7278),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7280),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7437));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7435));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7433));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7431));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7428));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7425));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7423));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7356),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7422));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7421));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7420));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222527 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7359),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7419));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7418));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222529 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7417));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7416));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222531 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7355),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7415));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6976),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7414));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1666));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7380),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7430));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222535 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7199),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7429));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7427));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7426));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7424));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1665));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222544 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7412));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222545 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7411));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222546 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7410));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222547 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_296),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7409));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222548 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7408));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222549 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7407));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7271),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7406));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7405));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222552 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7281),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7404));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222553 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7403));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222554 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1664));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7402));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222556 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7401));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222557 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7400));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7399));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7398));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222560 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7397));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222561 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7351),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7396));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222562 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .A2(n_14524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7395));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222563 (.A(n_14522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7394));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7346),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7393));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7392));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222566 (.A1(n_14522),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7391));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222567 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6870),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7389));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222569 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_293),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6886),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7387));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6883),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7291),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_294),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7386));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222571 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6881),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7285),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7385));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222572 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7329),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7384));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222573 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6877),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1658),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7327),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7383));
 AOI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222574 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7279),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7338),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6875),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7382));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6873),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7381));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222576 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7380));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7379));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1659),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7253),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7378));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7377));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1586),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7144),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7376));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222581 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6888),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7375));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222582 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6865),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7374));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222583 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6909),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7342),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7373));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1634),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7390));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222586 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7215),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7371));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7370));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7369));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7344),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7368));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7367));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7366));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7365));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7364));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7363));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7362));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222596 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7242),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7361));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7168),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7360));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7342),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7359));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7335),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7358));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7357));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7356));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7355));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7354));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7353));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7336),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7352));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7351));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222607_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_442));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7349));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222609 (.A(u6_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7350));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222610 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6995),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7348));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222612 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6971),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7346));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7345));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7344));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7343));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7340),
    .Y(u6_n_99));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7338));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222620 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6921),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7337));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222621 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7336));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222622 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6975),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7335));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222623 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6906),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7334));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7333));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222625 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6977),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7332));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222626 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7305),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7331));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222627 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7163),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7342));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222628 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1657),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7340));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7339));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7330));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7295),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7329));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7299),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7328));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7327));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7326));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7325));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7324));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7298),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7323));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7322));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7321));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7320));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7319));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7318));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7317));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7316));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7313));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7312));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7251),
    .B(n_13851),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7204),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_7200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7311));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6899),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7310));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7075),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7274),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7309));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222654 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7273),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7308));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1657),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7314));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222656 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1657),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1663));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222665 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1618),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7300));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222666 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7010),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7299));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222667 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1615),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7298));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222668 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6982),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7297));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222669 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1654),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7296));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222670 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7260),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7295));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222671 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6973),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7294));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222672 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7307));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222673 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1662));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222674 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1661));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222675 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7127),
    .A2(n_14480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7305));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222676 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1652),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7304));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222677 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7267),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7302));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222678 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7193),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7301));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7291));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1660));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1659));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1658));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7289));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7288));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7287));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7097),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7286));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7285));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7284));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7283));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7282));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7281));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7280));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7279));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7278));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222703 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6944),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7277));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222704 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7259),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7208),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7293));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222705 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7276));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7275));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222707 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7176),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7274));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7273));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222711 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1657));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7240),
    .B(n_14481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7271));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222714 (.A(n_14480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7270));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222717 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7265));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222718 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7264));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222719 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7263));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222720 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6938),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7262));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222721 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7232),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7261));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222722 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7231),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1656));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222724 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7267));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222725 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1644),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7266));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7260));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1653));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7258));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1649),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7257));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7256));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7255));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7254));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7253));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222738 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1655));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222739 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1638),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1654));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222740 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1652));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7259));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7252));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222744 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7247));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222745 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7246));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6920),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7251));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7016),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7249));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6989),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7248));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7162),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7244));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7202),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7243));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7242));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7241));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7219),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7240));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7239));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222757 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6922),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7237));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222758 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7162),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7236));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222759 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7005),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7235));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222760 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1648),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7234));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6915),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7238));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7232));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7231));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1650));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1649));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7228));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7227));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6907),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7138),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1651));
 AOI211x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7211),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6957),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7233));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222775 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7201),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6991),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7230));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222776 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7073),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7229));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222777 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7182),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6974),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7226));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222778 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7225));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7177),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7224));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7193),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7223));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222781 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7178),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7222));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222782 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7189),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7221));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7220));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6929),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7079),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6905),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7217));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1646),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7216));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7215));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7214));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6913),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7213));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7173),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7219));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7212));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1641),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6904),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7210));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7209));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7208));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1642),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7207));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1640),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7206));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222799 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7211));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7204));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1648));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6901),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_7160),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_7062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7200));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7199));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7147),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7198));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7145),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7197));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_871),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7203));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7078),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7202));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7060),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7201));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7195));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7192));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7188));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222816 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7196));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222817 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7187));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1631),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_7063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7186));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7123),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7185));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7184));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6989),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1647));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7194));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7193));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7191));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222825 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6996),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7189));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1646));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7181));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7177));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7173));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7171));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6893),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7170));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7169));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7168));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7157),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7120),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7183));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6928),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7167));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7182));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1597),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7028),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7180));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222840 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7178));
 AND4x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1634),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1610),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7176));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1584),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6891),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7174));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6950),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7172));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7165));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7160));
 NOR3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6937),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7159));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222850 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7158));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7157));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222852 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1604),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7156));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222853 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7155));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1645));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7166));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222856 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6967),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7164));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222857 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7163));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7162));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7161));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7078),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1644));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7154));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222863 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6967),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7153));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6967),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7152));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7151));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222866 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1643));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7150));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7145));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222873 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6960),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7144));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222875 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1605),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7142));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222876 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7008),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7141));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222877 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6910),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7140));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222878 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1596),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7139));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222879 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1594),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7138));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7149));
 AND4x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6904),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6945),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7148));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7074),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7137));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222883 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1614),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_7003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1642));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7136));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222885 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1617),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7147));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222886 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1641));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222887 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6899),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7135));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1616),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1640));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222889 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6970),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7134));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7146));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222891 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1587),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1639));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7133));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7131));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7126));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7119));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7118));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222902 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_531),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6887),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7117));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7116));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6906),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7115));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6887),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_795),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7114));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6971),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7113));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222907 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7132));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7112));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7130));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7129));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7128));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1620),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7111));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7127));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7110));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7109));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7108));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1638));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7125));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7107));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7106));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7124));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7105));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222923 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7007),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7104));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7024),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7103));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7123));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222926 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6876),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7122));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7102));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1588),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7101));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222929 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1588),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_564),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7100));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7099));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7098));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7097));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7096));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7095));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7094));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7004),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7121));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7093));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7023),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7092));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7091));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1617),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7089));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7088));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7087));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6986),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7086));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7085));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7084));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7083));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7082));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7120));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1637));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7080));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7077));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7071));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1635));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1634));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7067));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222963 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6826),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6850),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7066));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6896),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7065));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222965 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6856),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7064));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6852),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7063));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7062));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6951),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7061));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7060));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222970 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7059));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g222971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6843),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6856),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_687),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7058));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7081));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222973 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1588),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7057));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7056));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7055));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6928),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7054));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7053));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7079));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g222979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7078));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7052));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7051));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7050));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6942),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7049));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7048));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7076));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6939),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7047));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_796),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7046));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1605),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7045));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7044));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7043));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7042));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7075));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7041));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7040));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7074));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222996 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6860),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7039));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6935),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7038));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222998 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_74),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6856),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2418),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7073));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g222999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7037));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7036));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7034));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7033));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6932),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7032));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6911),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7031));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7030));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7072));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7028));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1636));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7069));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7068));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7027));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7023));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7017));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7014));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7013));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7012));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7010));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7009));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7007));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7005));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7004));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1622));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7000));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6999));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6995));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6993));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6992));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6991));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6988));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6986));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6983));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6982));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6980));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6977));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6976));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6975));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6973));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6971));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6969));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6967));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6966));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6965));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7026));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7025));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7024));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7022));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7021));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7019));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7018));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1633));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7016));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7015));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1632));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1631));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7011));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1630));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1629));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1628));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1627));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7008));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7006));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1626));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1625));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1624));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1623));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7003));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7001));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1621));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1620));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6998));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6996));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1619));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6994));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1618));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1617));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1616));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1615));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6990));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6989));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1614));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1613));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1612));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6987));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6985));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6984));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1611));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6981));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223125 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6979));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223126 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6978));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223127 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1610));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6974));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223129 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1609));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1608));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6972));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6970));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223133 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6968));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6963));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6960));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6958));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6956));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6953));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6948),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6949));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6947));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6945));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6943));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6942));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6940));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6937));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6935));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6932));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6930));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6928));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6926));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6925));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6922));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6921));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6919));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6917));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6915));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6914));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6913));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6911));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6909));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6907));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6906));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6903));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6901));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6899));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6898));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1590));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_381));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1591));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223208 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6896));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6895));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1607));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6894));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6962));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6961));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223214 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6959));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6957));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223216 (.A(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1606));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6955));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6863),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6893));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6954));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6952));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6892));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6891));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6890));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6951));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6950));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6948));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_74),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1605));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6946));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6944));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6941));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1604));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1603));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6939));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6938));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6936));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6934));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223237 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6933));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6889));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6931));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1602));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6929));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6927));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6881),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1601));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6799),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6828),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1600));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6924));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6923));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1599));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1598));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6920));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6918));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1597));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1596));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1595));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6916));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1594));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6912));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6910));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1593));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6908));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6905));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6904));
 AO221x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223262 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6783),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6782),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6902));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223263 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6773),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6900));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223264 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1582),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_734),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1592));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6887));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6885));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1588));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6883));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6881));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6879));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6877));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6875));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6873));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6870));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6868));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6866));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6864));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6888));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6886));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223287 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1589));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223288 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6884));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6882));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6880));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6878));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6784),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6876));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6786),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6874));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6842),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6872));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6785),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6871));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223296 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6665),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6869));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223297 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6645),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6867));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6865));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6863));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6860));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6858));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6856));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6854));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6853));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6802),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6852));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6850));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223309 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6764),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6849));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223310 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6800),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6848));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223312 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6742),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_6765),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6846));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223313 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1587));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6862));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6824),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6861));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6859));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6597),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6857));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6806),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6855));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1586));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1583));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223326 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6845));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6809),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6844));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6779),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6566),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6843));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6842));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6841));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223331 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6775),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6840));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223332 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6839));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223333 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6838));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6761),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6813),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6837));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223335 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6836));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223336 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1585));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223337 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1584));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6835));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223339 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6699),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6834));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223340 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6833));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223341 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6832));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223342 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_451),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6831));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6830));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223344 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6829));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223345 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6596),
    .A2(u6_n_101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6828));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223346 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6774),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6827));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6826));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6825));
 AOI32xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223349 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .A2(u6_n_101),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6824));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223350 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6823));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6822));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223352 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6667),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1474),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6821));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223353 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6644),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6820));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223354 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6664),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6819));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1472),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6818));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1494),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6817));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6816));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223358 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6750),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6531),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6815));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6814));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6729),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6813));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6723),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6812));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223362 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6811));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223363 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6694),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6810));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223364 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6660),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6809));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223365 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6808));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6807));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6806));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1577),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6805));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6767),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6804));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6802));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6800));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1470),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6801));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223375 (.A(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6799));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_480),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6798));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223377 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6740),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6797));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6748),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6796));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6795));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6738),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6741),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6794));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6793));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6792));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223383 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6791));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6790));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6789));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223386 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6788));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6787));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6786));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6785));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6784));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6767),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6783));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6782));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1582));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6781));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6779));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6780));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6597),
    .B(u6_n_101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6778));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6777));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6776));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6775));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6774));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6747),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6773));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6755),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6772));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6771));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6770));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1579),
    .Y(u6_n_101));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1579));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223413 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6768));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223415 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6718),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6433),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1577));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6734),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6767));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6766));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6765));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6764));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6763));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6762));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6761));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223423 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6625),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6688),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6595),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6760));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6759));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6758));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6757));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6756));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223428 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6719),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6432),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6755));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223429 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6754));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223430 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6537),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6718),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6536),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6752));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6751));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6750));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6716),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6749));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6748));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223435 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6722),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6747));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223436 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1575),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6746));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223437 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6711),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1523),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6753));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6743));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6742));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1576));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223443 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1570),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6615),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6741));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6535),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6740));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6739));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223446 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1526),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6616),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6738));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223447 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6711),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6737));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223448 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6362),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6736));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223449 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1477),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6735));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6734));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223451 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6364),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6733));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223452 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6745));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223453 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6647),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6675),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6744));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6732));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6731));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6706),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6730));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6729));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6728));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6727));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6726));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6725));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6724));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6723));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223465 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6617),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6722));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6720));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223467 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1571),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6721));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223469 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1575));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6718));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223471 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6719));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223472 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6717));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6684),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6716));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6715));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6714));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6533),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1571),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6532),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6713));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6709));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6708));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6707));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1565),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6706));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223484 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6371),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6705));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223485 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1564),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6367),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6704));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223486 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6677),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6703));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223487 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6542),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6712));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223488 (.A1(n_14482),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1574));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223489 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6711));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223490 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1541),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6710));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1573));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6702));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6701));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6700));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6699));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223496 (.A(n_14482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6698));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6697));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6696));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6695));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6694));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6693));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6692));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6691));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6690));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223505 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1527),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6576),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6689));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223506 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6556),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6688));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223508 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1559),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6375),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6431),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6686));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223510 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1507),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6430),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6684));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6683));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6428),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6682));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6681));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1572));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223516 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6611),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6680));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223517 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1518),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6470),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6573),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6679));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1571));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1570));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1561),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6678));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6676));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1565));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6674));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223533 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6652),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6673));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223534 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1488),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6672));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223535 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1504),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6671));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223536 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1562),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6670));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1560),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6374),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6669));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223538 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6480),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1535),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6677));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223539 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1560),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1569));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223541 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1561),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6599),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1567));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223542 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1562),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1566));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223543 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6614),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6675));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6668));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6667));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6666));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6665));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6653),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6664));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1556),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6642),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6663));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6662));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6661));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6660));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223555 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6561),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6659));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223556 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6482),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6649),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1564));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223557 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6363),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1510),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6462),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6658));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223558 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1544),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1478),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6657));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223559 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6656));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6626),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6655));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6624),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6654));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1562),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6651));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1562));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6649));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1560));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6543),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6618),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6647));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1533),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1563));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223576 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6593),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6653));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1534),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6652));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6592),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6650));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1561));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1554),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6648));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223581 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6549),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6646));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6645));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6644));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6643));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1476),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1490),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6642));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223586 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1487),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6641));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223587 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1483),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6640));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223588 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1553),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6639));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6638));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6636));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6634));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223594 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6538),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6630));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6629));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6637));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1526),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6635));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223598 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6633));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1514),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1542),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6631));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223600 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6472),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1559));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6628));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6626));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6624));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223605 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6622));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223606 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6567),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6627));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223607 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6621));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6424),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6433),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6625));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1519),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1522),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6623));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1518),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1523),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6620));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223611 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6569),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1558));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6619));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6616));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6539),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6548),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6614));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6484),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6613));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6612));
 NAND4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6540),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6546),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6611));
 NAND2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6610));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6609));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6618));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6617));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6608));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6607));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6606));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6568),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6605));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1549),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6604));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6615));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1552),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6603));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6602));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6601));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6599));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6595));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6593));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1555));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6591));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1553));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6589));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1536),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6587));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223647 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6586));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223648 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6585));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6600));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1537),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6584));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1538),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6583));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6508),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6582));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6509),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6477),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1557));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223654 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6483),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6598));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6581));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6597));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6494),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6596));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223658 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1556));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223659 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6178),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_871),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6594));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223660 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6504),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6592));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223661 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1554));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223662 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6552),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6588));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6577));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6575));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6572));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6570));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1546));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223676 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1545));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6568));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223678 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1552));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6580));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6579));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1551));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1550));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1549));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6578));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6576));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6574));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6573));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6571));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6567));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1548));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1547));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6569));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6566));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6564));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6562));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6559));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6557));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6396),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6565));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223703 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6377),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1529),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6555));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223704 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6422),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6563));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223705 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_287),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6554));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223706 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1475),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6553));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223707 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6552));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223708 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6305),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6551));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1544));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223710 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1543));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6550));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6549));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6561));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6560));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223715 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6558));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1542));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6556));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6548));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6546));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6544));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6542));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6540));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223724 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6539));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6537));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6535));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6533));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1540));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6530));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6528));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6547));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6340),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6527));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6332),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6526));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223737 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6525));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1484),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6524));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6545));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223740 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6543));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6523));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6522));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223743 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6541));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1541));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6538));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6536));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6521));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6474),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6520));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6519));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6471),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6518));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6467),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6517));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6516));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6534));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6515));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6532));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223757 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6359),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6514));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6513));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6279),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1539));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6420),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6531));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6278),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6529));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6512));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6510));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6507));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223769 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1501),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6506));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223770 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6505));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223771 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6504));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6328),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1502),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6503));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6339),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6502));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6349),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6501));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223775 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6331),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6500));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223776 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6499));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223777 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6498));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223778 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6497));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6437),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6496));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223780 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6327),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6495));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223781 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6494));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223782 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6493));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6492));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6491));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223785 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1481),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1538));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1517),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6490));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1506),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6511));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1479),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1537));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6489));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6488));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1486),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6509));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6341),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1536));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1535));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6487));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223795 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6486));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_803),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6485));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6508));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6484));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6481));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6480));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6478));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6476));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6473));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6471));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6469));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6467));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6466));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6465));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6464));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6463));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6461));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6460));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6483));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1534));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1533));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1532));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1504),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6482));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223840 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6293),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6459));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6458));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_795),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1531));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6341),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1530));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223844 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6479));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6298),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6293),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6457));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6456));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6455));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6454));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6453));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223850 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6477));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6452));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6451));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6450));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6475));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1510),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6449));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6448));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6474));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6447));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6446));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6445));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6444));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6387),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6443));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6442));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6391),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6441));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6440));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6472));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6470));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1529));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6468));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1528));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1527));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1526));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1525));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1524));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1523));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1522));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223877 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6462));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1521));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1520));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1519));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1518));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6438));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6437));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6435));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6432));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6429));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6428));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6426));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6425));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6424));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223902 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6214),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6273),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6423));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_686),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6422));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6214),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6285),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6421));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6420));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g223906 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6272),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6419));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223907 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6418));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6417));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223909 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1472),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_795),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6416));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6415));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6414));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6413));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223913 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6293),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6412));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6411));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6439));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6410));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6409));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6436));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6434));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6344),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6408));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6347),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6407));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223923 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6406));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223924 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2840),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6302),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6405));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6404));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6335),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6403));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6402));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6401));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6400));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6399));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6398));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223933 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6397));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223934 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1470),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6396));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6433));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6431));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6395));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6394));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6430));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1517));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1516));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6427));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1515));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1514));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1513));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6393));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1512));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1511));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6391));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6389));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6387));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6384));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6382));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6380));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6379));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6378));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6376));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6372));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6370));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6369));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6366));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6365));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1497));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6364));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6362));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6361));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6359));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6357));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6355));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1494));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6352));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6392));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6390));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6388));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g223997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6386));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6351));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g223999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6385));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6383));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6381));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1510));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1509));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6377));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6350));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1508));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6349));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6375));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6348));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6374));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6373));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1507));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1506));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1505));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224015 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1504));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6371));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1503));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6368));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1502));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6367));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1501));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1500));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1499));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1498));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6363));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1496));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1495));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224028 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6193),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6360));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6358));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224030 (.A(n_14526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6356));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224031 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6203),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6354));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6353));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6347));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6345));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6344));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6342));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6340));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6338));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6336));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6335));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6333));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6332));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6330));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1484));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6327));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6326));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6325));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6324));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1476));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6323),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6322));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6320));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224072 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1463),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6319));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224073 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1463),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6318));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6274),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6317));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224075 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6316));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1493));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6315));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6314));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6313));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6312));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6311));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6346));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1492));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1491));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6343));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1490));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6341));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6310));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1489));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6309));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6339));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6308));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6337));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1488));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6334));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1487));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1486));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6331));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1485));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6329));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6328));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1483));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6307));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1482));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1481));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1480));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1479));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1478));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1477));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6323));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224111 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2736),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6321));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6306));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1474));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6304));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6302));
 INVx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6301));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224128 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1472));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6298));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6295));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6293));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6290));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6286));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224142 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1432),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6075),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6285));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224143 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6305));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224144 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2518),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1475));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1473));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6303));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224147 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_283),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6300));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6299));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1471));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6296));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6294));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6292));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6291));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224154 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6151),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1466),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6288));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6287));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1470));
 AOI322xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224161 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6180),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2641),
    .B1(n_3627),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6154),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_1462),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_2823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6284));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224162 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6283));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224163 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6282));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224164 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6281));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224165 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6280));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6279));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6278));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224168 (.A(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6277));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6214),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6276));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6275));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6274));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6273));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6272));
 AO22x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224174 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2651),
    .A2(u6_n_102),
    .B1(n_3626),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1469));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224175 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6271));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224176 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6270));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224177 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6269));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224178 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6268));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224179 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6202),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6267));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224180 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6199),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6266));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224181 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_285),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6265));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224182 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6264));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224183 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1354),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6194),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6263));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6262));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224185 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6074),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6261));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6260));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6259));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6258));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224189 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6257));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224190 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6256));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6255));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6254));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6200),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6253));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6208),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6252));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6251));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6250));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6249));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6248));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6247));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6056),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6246));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224203 (.A(u6_n_102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1468));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224204 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6071),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6245));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224205 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6109),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6244));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224206 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6243));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224207 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6050),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6242));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224208 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6149),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1463),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6241));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224209 (.A1(n_14282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1356),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6240));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224210 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1455),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6150),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6239));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224211 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6085),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6238));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224212 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1340),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6237));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224213 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6152),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6236));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224214 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_284),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6235));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224215 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6173),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6044),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_1406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6234));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224216 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6183),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6233));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224217 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5902),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6232));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .Y(u6_n_102));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6231));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6230));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224221 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6107),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6229));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224223 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6227));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224224 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6190),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6226));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6225));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224226 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6139),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6224));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6137),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6223));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224228 (.A1(n_14484),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6222));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6221));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6220));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6219));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6218));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224233 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6217));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6216));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1466));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6214));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6213));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6212));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5856),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6211));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1406),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6210));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5812),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6209));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6170),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6208));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224247 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5864),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6207));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224248 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6206));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5825),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6205));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224250_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_412));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224251_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_448));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6204));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6203));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6202));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6201));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6200));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6199));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6198));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6197));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6196));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6195));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6194));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6193));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224265 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5885),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1402),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6190));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224266 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6131),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5886),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5992),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6189));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6188));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5785),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6187));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6186));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6192));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6185));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6181));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6178));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1463));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1462));
 BUFx6f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1464));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6176));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224284 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6133),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6174));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6047),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6184));
 AOI21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224286 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6133),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6183));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6132),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6180));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5678),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6179));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224289 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6078),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6177));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6172));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224296 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6098),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6125),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6168));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224297 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6066),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6104),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6167));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224298 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5896),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6166));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224299 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1382),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1454),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6165));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224300 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5863),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6164));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224301 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5859),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6163));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224302 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6118),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6162));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224303 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6173));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224304 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5997),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1461));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224305 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5970),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1460));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1418),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1459));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224307 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6126),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6171));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6116),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6170));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224309 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5987),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1452),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1458));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6155));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1456));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1457));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1455));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6154));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224327 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6153));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6152));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6151));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1454),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6150));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6149));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6148));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6146));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6145));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6144));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6126),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5818),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5815),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6143));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224339 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5880),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6142));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224340 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6118),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6156));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6141));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224342 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5829),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1374),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6140));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6096),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5954),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6139));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6138));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224345 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5869),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6137));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224346 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1446),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1397),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5956),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6136));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6133));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6132));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6131));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1453));
 A2O1A1O1Ixp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5952),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5945),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5697),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6125));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5872),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6124));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5817),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6123));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224362 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6092),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6122));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224363 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1449),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1372),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6121));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224364 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1446),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6130));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224365 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6129));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5979),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6093),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1454));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224367 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1447),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6128));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1434),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6093),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6126));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6034),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1452));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6120));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6116));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6115));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224375 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6114));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6068),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1451),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5698),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_6087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6113));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6112));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6031),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6099),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6111));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6110));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6083),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6109));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6089),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6118));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6092),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6117));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6108));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5951),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6107));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224387 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5948),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6105));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224388 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5947),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1417),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6104));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224389 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6027),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1444),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6103));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6100));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6095));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6093));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224400 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5898),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1409),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6091));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224401 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1408),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5901),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6090));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5857),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1425),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1403),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5900),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1451));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224403 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5888),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6101));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224404 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1395),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5883),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5847),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5851),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6099));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224406 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5978),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6096));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224407 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1441),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1421),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1450));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224408 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6007),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1449));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224409 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1440),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6092));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1448));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1446));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1445));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6088));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1407),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1433),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1436),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5946),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_6041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6087));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6086));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1441),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6085));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224423 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6045),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6084));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224424 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1441),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6083));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224426 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5837),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6081));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224427 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6037),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1447));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224428 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1438),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6035),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6089));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6080));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224430 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6079));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6067),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6078));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6047),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6077));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6074));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6073));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224439 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1412),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1386),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1393),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6072));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6071));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6014),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6070));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224442 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6002),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1428),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1444));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224443 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6042),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6075));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224444 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6069));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224445 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6036),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1443));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1441));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1439));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224456 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5981),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1426),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6064));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224457 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6025),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6063));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224458 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5977),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1429),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6062));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5985),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6068));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224460 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5982),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_6023),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1442));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5944),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6028),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6067));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1432),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5947),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6066));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224463 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6038),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1440));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1375),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1438));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6045),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6061));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1423),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5988),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6060));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224467 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1365),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1370),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6059));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6003),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_6004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6058));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1437),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6057));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6046),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6056));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6055));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224472 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6054));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5911),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1362),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5928),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6053));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5910),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6052));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6051));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6050));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6049));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1436),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6046));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6044));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1432));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224489 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6041));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1421),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5832),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6040));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6039));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224492 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6038));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5874),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6037));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224494 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6036));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5827),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1379),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6035));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1437));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6047));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1436));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1364),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5857),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1435));
 NAND4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5893),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5886),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6034));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5809),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6045));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224502 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1391),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6033));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224503 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1391),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6032));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5901),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6031));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224505 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1391),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6030));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1381),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1382),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1434));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224507 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6029));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6028));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1433));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6042));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6024));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6022));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224522 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5840),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6020));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224523 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1368),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6019));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224524 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5874),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6018));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224525 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1374),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5875),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6017));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224526 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6016));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1431));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1418),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1430));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224529 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5819),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5796),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1429));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224530 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1365),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6015));
 NAND4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1409),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1396),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5861),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6027));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5869),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5881),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1428));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224533 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5835),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6025));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224534 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1405),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1427));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224535 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1384),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5801),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6023));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224536 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1380),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1426));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1404),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5848),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6021));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224538 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1375),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5813),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6014));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224539 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2762),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6013));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6012));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224541 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1413),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1363),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1425));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224542 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1412),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6011));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1424));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6010));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6008));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6007));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6005));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6003));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6001));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5997));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5994),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5995));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5993));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1419));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5989));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5988));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5987));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5699),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5986));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5985));
 AO22x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224568 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6009));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224569 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5984));
 AO22x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1352),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1423));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224571 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5983));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224572 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1354),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1422));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224573 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5982));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224574 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5981));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5766),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5980));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5979));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5978));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6006));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5977));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224580 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1421));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1401),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6004));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5976));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224583 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6002));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5891),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5975));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224585 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5787),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5974));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5856),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5973));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5972));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5878),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5971));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5970));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5969));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5968));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1366),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6000));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5967));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5906),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5966));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1396),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5998));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1408),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5965));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224597 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1354),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_390),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5996));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1416),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5964));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5994));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5896),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5963));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224601 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_226),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1354),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5962));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5992));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224603 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5961));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5887),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5960));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5959));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5958));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5990));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5957));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5955));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5950),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5951));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5945));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224616 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5944));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5943));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5956));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224619 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_610),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1340),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5942));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224620 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5954));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224621 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5941));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5940));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5953));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224624 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1418));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5939));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5938));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5937));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224628 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_852),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5936));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224629 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5935));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224630 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5934));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224631 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5933));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5932));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224633 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5931));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5930));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224635 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_795),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5929));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5952));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5928));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5927));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5836),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5926));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1380),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5925));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224641 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5924));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1384),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5923));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5922));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224644 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5776),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5921));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1374),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5950));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5920));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5948));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224648 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2418),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5919));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5918));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5917));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5916));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5915));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_831),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5914));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1385),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1364),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5913));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5947));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1417));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5912));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5946));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5911));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5910));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5908));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5906));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5904));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5903));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5902));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5899));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5897));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5895));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5894));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224693 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5893));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5891));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224695 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5889));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5887));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5885));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5884));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224704 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1401));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5880));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5878));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224707 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5876));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1399));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5873));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5871));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5868));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5865),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5866));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5864));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224723 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5863));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5861));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5860),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5859));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5858));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5856));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5855));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1390),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1391));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1390));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5853));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5909));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5907));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5905));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_94),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1416));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5852));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1415));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224748 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5851));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1414));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5850));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5849));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1413));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1412));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1411));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1410));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1409));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5901));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5900));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5898));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1408));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1407));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224762 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1406));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1405));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5896));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1404));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5848));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1403));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5892));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5890));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5847));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5888));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1402));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5886));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5883));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5881));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5879));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5877));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5875));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1400));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5874));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5872));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1398));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5869));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1397));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5865));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1395));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_94),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5862));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5860));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1394));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5857));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1393));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2733),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5854));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5846));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5845));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5843));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224803 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5842));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5841));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5838));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5835),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5836));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5834));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1378));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5832));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5829));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5826));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5825));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1371));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5820));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5817));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5815));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1364));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5814));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5813));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5812));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1359));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5810));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5809));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5808));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5807));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1389));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1388));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5806));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1387));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5804));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5803));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1386));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1385));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5844));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1384));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1383));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1382));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224876 (.A(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5840));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2840),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5801));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1381));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5837));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5835));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1380));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1379));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1377));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5831));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5800));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1376));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1375));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5799));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5827));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1374));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1373));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1372));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5824));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5821));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5798));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1370));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5819));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5797));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1369));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1356),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5818));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1368));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1367));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5796));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224905 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1366));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1365));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224907 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1363));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5795));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5794));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1362));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224911 (.A1(n_3628),
    .A2(u6_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5759),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1361));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1360));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224913 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5309),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5811));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224916 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1358));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1357));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224923 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5787));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5785));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5783));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1356));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1355));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1354));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224949 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5736),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5777));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5793));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5789));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5704),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5788));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5786));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5784));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5782));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5706),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5781));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5779));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5778));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g224961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5776));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1352));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1350));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1348));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g224991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1345));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g224998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1343));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1341));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1340));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1339));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225020 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5761));
 AOI221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5685),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1332),
    .B2(n_3629),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5760));
 OA22x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225022 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2653),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5736),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2461),
    .B2(u6_n_104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1353));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5775));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5773));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5771));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1346));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5746),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5757),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5768));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5766));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5763));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1338));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225031 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5684),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5758));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225032 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5688),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5686),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5757));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225033 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5756));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225034 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5755));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225035 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5650),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5754));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225036 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5753));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225037 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5730),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5752));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225038 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5751));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225039 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5617),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5750));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225040 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5622),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5749));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225041 (.A(u6_n_104),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5759));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225042 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5587),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5748));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225043 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5644),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5747));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225044 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1334),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5746));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225045 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5745));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225046 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5744));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225047 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5618),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5743));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5742));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225049 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5741));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225050 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5740));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5701),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5739));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5502),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5738));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225053 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5619),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5735));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5734));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225055 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5651),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5733));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225056 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5638),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5732));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225057 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_282),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5731));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225058 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5669),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5730));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225059 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5646),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1331),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5729));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225060 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5653),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5624),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5728));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225061 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5621),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5727));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225062 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5726));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225063 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5649),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5725));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225064 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5583),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5724));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225065 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5614),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5723));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225066 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5589),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5722));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225067 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_281),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5721));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225068 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_258),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1252),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5720));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225069 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5567),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5719));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1332),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .Y(u6_n_104));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5736));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5718));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5717));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225074 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5660),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5716));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5623),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5715));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5548),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5714));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5590),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5713));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5564),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5712));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5711));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5710));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225081 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5632),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5709));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5708));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5586),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5707));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5706));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5705));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225086 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5663),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5704));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225087 (.A(n_14283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5703));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5702));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5666),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5701));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5700));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5697));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5695));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5694));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5692));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5691));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5679),
    .B(n_14164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5699));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5698));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5690));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225104 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1332),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5696));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225105_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .B(u6_n_105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_235));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5680),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5693));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5689));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5688));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225109 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5687));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5658),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5686));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5685));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5684));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5683));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225114 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5344),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5682));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225115 (.A(u6_n_105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5680));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225116 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5678));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225117 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5552),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1327),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5677));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5676));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5675));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225120 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5565),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5661),
    .Y(u6_n_105));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5679));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5674));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1335));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225129 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1334));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5669));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5444),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5668));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5642),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1282),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5667));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225134 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5666));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225135 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5607),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5670));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225136 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5558),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5612),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5664));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225137 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5364),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1287),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5663));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225138 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5539),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5662));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225139 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5470),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1327),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5534),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5661));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225140 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5559),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5610),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5660));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225141 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5659));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225142 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1280),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5658));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225143 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5637),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5343),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5657));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225144 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5656));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5655));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225146 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1328),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5665));
 BUFx6f_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5654));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1331));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5653));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1332));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5652));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5651));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1328),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5650));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5649));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5431),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5648));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5646));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5645));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5644));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1330),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5643));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1333));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1316),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5642));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225171 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5641));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225172 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5640));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225173 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5609),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5337),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1297),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5639));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5414),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5638));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5634));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225178 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5403),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5633));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5452),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5632));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225180 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5631));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225181 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1270),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5319),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5630));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225182 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5629));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225183 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5601),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5628));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5603),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1293),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5627));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225185 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5376),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5626));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5465),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1330));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5601),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5637));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1307),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5635));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1329));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5624));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225195 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5623));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5622));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5621));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1324),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5620));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5619));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5618));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225201 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5617));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5616));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5615));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5614));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5593),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5613));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225206 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5537),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1328));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5612));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1283),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1290),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1306),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5610));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225211 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1279),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5369),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5422),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1327));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5609));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5608));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225214 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5536),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5607));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5606));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225219 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1326));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225220 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1322),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5499),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5604));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5600));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5577),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5329),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5597));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225228 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1276),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5596));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225229 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5335),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5595));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5323),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5594));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5368),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5593));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1273),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5592));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5603));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225234 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5458),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5602));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5574),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1325));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1317),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5601));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1324));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225238 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1321),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5498),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1323));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5429),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5591));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5590));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5589));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5588));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5587));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5586));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1281),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1295),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5585));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5584));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5583));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1317),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5582));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5550),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5581));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5580));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225252 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5384),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5579));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225254 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1286),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1322));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225255 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5324),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5545),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5578));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5574));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1321));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1320));
 NOR4xp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1315),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5450),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5568));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225265 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5528),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5577));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225266 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1304),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5576));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225267 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5575));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225268 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5573));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225269 (.A1(n_13869),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5571));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225270 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1312),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5569));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5567));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225272 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1316),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5566));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5541),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5565));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5564));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5563));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225276 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1312),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5562));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225277 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1313),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5316),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5561));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225278 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1314),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5560));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5559));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225283 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1280),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5555));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225284 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5483),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5554));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5518),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5553));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1319));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225287 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1315),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5558));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225288 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1311),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5556));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5552));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1318));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225293 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5489),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5436),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5549));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5471),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5548));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5472),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5547));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5473),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5546));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225297 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5509),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1278),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5545));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225298 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5493),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5544));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225299 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5543));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225300 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5491),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5453),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1317));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225301 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5487),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5550));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225302 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5542));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5540));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1315),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5538));
 NAND5xp2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5466),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5458),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_5361),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_5349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5537));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5454),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5536));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5512),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5464),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5535));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225311 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5223),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5196),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5534));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225312 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5420),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1285),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5541));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225313 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5420),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5539));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225314 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5420),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5533));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225315 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_829),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5420),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1316));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5532));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5420),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1315));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1314));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5531));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225322 (.A(n_13869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1313));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5528));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5221),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5195),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5526));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225328 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_576),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5525));
 OAI221xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5278),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_835),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2990),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5524));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5197),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5523));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5522));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5419),
    .B(n_13857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5530));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5476),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1312));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5521));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5517));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5514));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5508));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5422),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5520));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5358),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5507));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5423),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5351),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5506));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5295),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5505));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5320),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5504));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225349 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5366),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5518));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225350 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5503));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_563),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5502));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225352 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5516));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225353 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5515));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5462),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5501));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5513));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5500));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5448),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5512));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5499));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1286),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5498));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5511));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5509));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5321),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5497));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1311));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5496));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5494));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5492));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5488));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5486));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5484));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225373 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5336),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5481));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5357),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1274),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5480));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5296),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1271),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5479));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225376 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5313),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5478));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5291),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5304),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5476));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5474));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225381 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1268),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1310));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225382 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5309),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5495));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225383 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1275),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5316),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5493));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5473));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225385 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1276),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5491));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1267),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5489));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5472));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225388 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1289),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5334),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5487));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5381),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5485));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5471));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225391 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5470));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5483));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5469));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5466));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5464));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5462));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5459));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5457));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5455));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5454));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5452));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5450));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5468));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1272),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5449));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5448));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225413 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5465));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225414 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1309));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225415 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5461));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5458));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5447));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5456));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225419 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1308));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5269),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5453));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225421 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5446));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225422 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5445));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1284),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5444));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5370),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5443));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5451));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225426 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5442));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5352),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1303),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5441));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225428 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_94),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1307));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1296),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5440));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5439));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225431 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_94),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5438));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225432 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5437));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5436));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5381),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5435));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5434));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5433));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5348),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5432));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225438 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5431));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5365),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5430));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225440 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5429));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225441 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_533),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5428));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225442 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5427));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1301),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5426));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5425));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1306));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5424));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5420));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225450 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5419));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5418));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225452 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5417));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225453 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5416));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1278),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5415));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225455 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_829),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5414));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1295),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5413));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1272),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5412));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225458 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1259),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5411));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5272),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5410));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225460 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5409));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225461 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5408));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225462 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2840),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5407));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225463 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_36),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5406));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1250),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5405));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225465 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5404));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5403));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225467 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_114),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5402));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225468 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1250),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5401));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5400));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1277),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1305));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5399));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1275),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5423));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225473 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5398));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225474 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5326),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5397));
 AO22x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225475 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1304));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5396));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1252),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5395));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225478 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5394));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225479 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5393));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225480 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1250),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5392));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_5263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5391));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5390));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225483 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5314),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5389));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5388));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225485 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5422));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5421));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5387));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1298),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5386));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5385));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5384));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5383));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5376));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1292),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1293));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5374));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5372));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225514 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5371));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5370));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5367));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5365));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1288),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5364));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1287),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5362));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5361));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5360));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5358));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5356));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5353));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5351));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1284));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5349),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5348));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5347));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1282));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5344));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5343));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_58),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5342));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1303));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1302));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5341));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5340));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5339));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1301));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5338));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1300));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1299));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5337));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1298));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1297));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1296));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1295));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1294));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5381));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5379));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5377));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225570 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5375));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1292));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5373));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1291));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1290));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5336));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5369));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5368));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5366));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5335));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1289));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5334));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1288));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1287));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1286));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5359));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1285));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5357));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5355));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5352));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_58),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5350));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1283));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5349));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5345));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1281));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1280));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1279));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1278));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5333));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5331));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5329));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5327));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5326));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5324));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5322),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5323));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5320),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5321));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5318),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5319));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5312));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5310),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5311));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1266));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1265));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225635 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5206),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5307));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5306));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5305));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5304));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5332));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5330));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5301));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5300));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5299));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5298));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5297));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5296));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5295));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1277));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1276));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1275));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5294));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5328));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_58),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1274));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1273));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5325));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225658 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1272));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5293));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225660 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5292));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5291));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5322));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1271));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5290));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5320));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1270));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5318));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1269));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5316));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5314));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5313));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1268));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5288));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225676 (.A(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1267));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5287));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5285));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5310));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225681 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4804),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5309));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5308));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1264));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225701 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1262));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5278));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1261),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5277));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1259));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5272));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5269));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1256));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225743 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5282));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1263));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5279));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1261));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1260));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225748 (.A1(n_14284),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1258));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5238),
    .B(n_14485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_408));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_277),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1255));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5265));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5263));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5260));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1252));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5258),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1253));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225774 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1250));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1249));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5253));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5251));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5250));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5207),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5249));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5262));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1254));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5258));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2728),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5203),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1251));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_395));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225793 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5254));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5252));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225795 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5158),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5248));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5247));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5246));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225798 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5199),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5245));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5125),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5244));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5243));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5242));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5160),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5241));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .B(n_3630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5240));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225804 (.A1(n_14285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5239));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_275),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5238));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_278),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5237));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5236));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5235));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4897),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5234));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225810 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5233));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225811 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5232));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5231));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225813 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1248),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5230));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1174),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5225));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225816 (.A(n_14286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5224));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5223));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_846),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5222));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5221));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5220));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225821 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5229));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5219));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5218));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225825 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5228));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5226));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225827 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5072),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5216));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5215));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5214));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225830 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5031),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5213));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5212));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5211));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5210));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225834 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5175),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5209));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5208));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_274),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5207));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5206));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5205));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5204));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5203));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1248));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225848 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1244),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1238),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5199));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225849 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .B(n_14528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5198));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5197));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5196));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5195));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225853 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(n_14486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5194));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225854 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5193));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2454),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5192));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225856 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4773),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5191));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225857_0 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_410));
 OR2x6_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5200));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225859 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5018),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5190));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4785),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5189));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5188));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225862 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_279),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5187));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225863 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5053),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5186));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5185));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5184));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225866 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5149),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5183));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225867 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5151),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5182));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5181));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5180));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5179));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1247));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225876 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5034),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5051),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5175));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225877 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5074),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5076),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5174));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225878 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5110),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5036),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5049),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5173));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225880 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5083),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5084),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5171));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225881 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5115),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5170));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225882 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1246),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5169));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225883 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1199),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5168));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225884 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4956),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5167));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225885 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4805),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5166));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225886 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5056),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5177));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5176));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5082),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5165));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225889 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5118),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5164));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225890 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2799),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2802),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5163));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225892 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5001),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5000),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5161));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5160));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5159));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5158));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5157));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5156));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5155));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5154));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5153));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225901 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4820),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4926),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5152));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5151));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225903 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4820),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4816),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5150));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225904 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1194),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1178),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5149));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225905 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1193),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4928),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5148));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5146));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225907 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5045),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5147));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225908 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5112),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4903),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5145));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225909 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5110),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5144));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225911 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5136));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5140));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225917 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5048),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5137));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5110),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5135));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5014),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5133));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225923 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4697),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4699),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5132));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225924 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5131));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225925 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4836),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5130));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225926 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4871),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5129));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225927 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5098),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5128));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4948),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5134));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225929 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4944),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5094),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1246));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225930 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4947),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5098),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1245));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1244));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225935 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1243));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5126));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5125));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5085),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5124));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5086),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5120));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5088),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5119));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225945 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5032),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5127));
 OAI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225946 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5070),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4821),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5118));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225947 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5097),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5117));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225948 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4823),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1195),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5116));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4930),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5115));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5112));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5029),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5111));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5110));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1242));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225959 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5028),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5109));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225960 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5078),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5108));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5097));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5095));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5010),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5033),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4983),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4971),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2996),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5093));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225972 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4982),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4970),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5092));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225973 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4826),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5107));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225974 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1240),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5105));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225975 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1224),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5103));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225976 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4961),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5102));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225977 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4995),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5098));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225978 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5064),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1241));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5094));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5052),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5091));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225984 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5041),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5062),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5090));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225985 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5043),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5054),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5089));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225986 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5071),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5088));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5087));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g225988 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1204),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5086));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225989 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4855),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5085));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5084));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5083));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5082));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5081));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5080));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225997 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5077));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g225998 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4910),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5076));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g225999 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4866),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5046),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5075));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226000 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5026),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4807),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5074));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226001 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1234),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4914),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5073));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4810),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4809),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5072));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226003 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5078));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5070),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5069));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1240));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5064));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226016 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1216),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1199),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1201),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5062));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1221),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5071));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226018 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5070));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226019 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1234),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5068));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226020 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5021),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5066));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4999),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5023),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1239));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5059));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5057));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4982),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1229),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4956),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5056));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226028 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1236),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4906),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1237),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5055));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226029 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1197),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1177),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1180),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5054));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5024),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5053));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226031 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1236),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4812),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5052));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226032 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_5022),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5058));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5051));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4983),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_5006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5048));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226037 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4991),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5047));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226038 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4980),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5046));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5034),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4902),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5045));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226040 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1222),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_5004),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5049));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226041 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1230),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1238));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5042));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5040));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226045 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4984),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5039));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226046 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1228),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4977),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5038));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226047 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4988),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5037));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1227),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5043));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226049 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4966),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5041));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5036));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4899),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5033));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5013),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5032));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226054 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2783),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_140),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5031));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226055 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2782),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4846),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5030));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4990),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4964),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5029));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4967),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5028));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5034));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5027));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5026));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5024));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1237));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1236));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1235));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5021),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1234));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4946),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5020));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4945),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5019));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5018));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5017));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5016));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5015));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226077 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1165),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5023));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226078 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4979),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4796),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5022));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226079 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4788),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4972),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5021));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5012));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5008));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5006));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1229));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5005));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4916),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4850),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5003));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1221),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4858),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5002));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226094 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4771),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5001));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1165),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5000));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4999));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226097 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_14),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4802),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4998));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1233));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4997));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4996));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4995));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4901),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5014));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4994));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226104 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1232));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1209),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4866),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5013));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5011));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5010));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1199),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1207),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4848),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5009));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5007));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4993));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1231));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1230));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5004));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4992));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4989));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4987));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4985));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4981));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226121 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4979));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226122 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4978));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226123 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4857),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4977));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4862),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4976));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226125 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4849),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1203),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4975));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226126 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4793),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4974));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226127 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4798),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4973));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226128 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4972));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226129 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4803),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4971));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226130 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4710),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4970));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226131 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1215),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4991));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4790),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4814),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4990));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226133 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4988));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4969));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226135 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1190),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1228));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226136 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1205),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4986));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226137 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4799),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1227));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226138 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1189),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4984));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226139 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_835),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4983));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226140 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4803),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4982));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226141 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4872),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1209),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4980));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226142 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4968));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226144 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4967));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4964));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4961));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4957),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4958));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4955));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4954));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4953));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4952));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226159 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1226));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1173),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4966));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4951));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226162 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1225));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226163 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4950));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1224));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226165 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4949));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4948));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4947));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226168 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1173),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4963));
 AO22x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226169 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4962));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226170 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4960));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226171 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4946));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4945));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4944));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4959));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1215),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1206),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4943));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4942));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4941));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4940));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4939));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4938));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4875),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4937));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4936));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226184 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4935));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226185 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1171),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4934));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4933));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1168),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4932));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1223));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4957));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4956));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1222));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4930));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4927),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4928));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4922),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4923));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4921));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4919));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4917));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226201 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4915));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4913));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4911));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4909));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4907));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4905));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4902));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4901));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4896));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4897));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226214 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4894));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226215 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4893));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226216 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4892));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226217 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_58),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4891));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4818),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4890));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226219 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1166),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4931));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4929));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4889));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226222 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2766),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4888));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226223 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4887));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1197),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1188),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4927));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4926));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4924));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4922));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4920));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1160),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4918));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226231 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1191),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4916));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4851),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4886));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4762),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1221));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4828),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4914));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4885));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1160),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4884));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1166),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4883));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1189),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4912));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4834),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4910));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4908));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4882));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4906));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4881));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4904));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4808),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4880));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4903));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1220));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4899));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4761),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4895));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4878));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4876));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4875));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1212));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4872),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4874));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226270 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4870),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4871));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226274 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1210));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4869));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4867));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4865));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4863));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4861));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226281 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4858));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1207));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4856));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4854));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4852),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4853));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4851));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4850));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4846));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4845));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4844));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1219));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_56),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4843));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4842));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4841));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4879));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4840));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226311 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4839));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226312 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1218));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1217));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2500),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1216));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1215));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1214));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226317 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1213));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1211));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4872));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4870));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226321 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1209));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226322 (.A(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4868));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4838));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_68),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4866));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4837));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4864));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226327 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4862));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4836));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4859));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226330 (.A(u6_rem_96_22_Y_u6_div_90_17_n_56),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4857));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1208));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226332 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1206));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1205));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226334 (.A(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4855));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1204));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226336 (.A(u6_rem_96_22_Y_u6_div_90_17_n_56),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1203));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226337 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4852));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1202));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1201));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4849));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4835));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4848));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_140));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226344 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1200));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1199));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1198));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4833),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4834));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4831));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4829));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4827),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4828));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4825));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4822));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226359 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4821));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1194));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4819),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4820));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4817),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4818));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4816));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4813));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226380 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4811));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4810));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4809));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4808));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4807));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1181));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1179));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4805));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4803));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4802),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4801));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226409 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4800));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4799));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4798));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4797));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4796));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226414 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4833));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4832));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4830));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1197));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226418 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4827));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4795));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226420 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4794));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4826));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1196));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4823));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1195));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1193));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4793));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4819));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4792));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4817));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1192));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1191));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4791));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1190));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2816),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1189));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1188));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4790));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226437 (.A(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4814));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4789));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226439 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1187));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4812));
 AOI221xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226441 (.A1(u6_n_108),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2648),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1159),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2463),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1186));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4788));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226443 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1185));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1184));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1183));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1182));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4787));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1180));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1178));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1177));
 OA21x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226451 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4804));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4802));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4785));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1176));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4783));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1174));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1173));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1171));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226474 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1172));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226479 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1170));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4778));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1168));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1169));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1166));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1167));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4775));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4773),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4772));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4750),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4786));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4751),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4784));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226501 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4683),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1175));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4782));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226503 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4654),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4781));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226504 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_270),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4779));
 NOR2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4747),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4777));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226506 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4650),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4774));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226507 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_272),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4714),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4773));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4771));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1163),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1164));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1162));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1160));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4766),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1161));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4764));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4762));
 XNOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226528 (.B(u6_rem_96_22_Y_u6_div_90_17_n_4559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4761),
    .A(u6_rem_96_22_Y_u6_div_90_17_n_4730));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226529 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1101),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1155),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4760));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226530 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(n_14287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4759));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226531 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1159),
    .A2(n_3632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1165));
 AO22x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226532 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2647),
    .A2(u6_n_108),
    .B1(n_3632),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1163));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4768));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4766));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4754),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4765));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4735),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4763));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226537 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4651),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4758));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226538 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4679),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4757));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226539 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4756));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226540 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4755));
 AOI32xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226541 (.A1(u6_n_109),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2632),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4691),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4754));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226542 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4583),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4753));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226543 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4752));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226544 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4751));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226545 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4750));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226546 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4749));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226547 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4748));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226548 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4732),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4747));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226549 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4686),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4746));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226550 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4624),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4745));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226551 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4744));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226552 (.A1(n_3633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1154),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4743));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226554 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1090),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4741));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226555 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4371),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4740));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226556 (.A1(n_14288),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1156),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1097),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4739));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226557 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1095),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .B(n_14487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4738));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226558 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4684),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4737));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226559 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4680),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4736));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226560 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4563),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4735));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226561 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4653),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4734));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226562 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4733));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226563 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_221),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4732));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226564 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1079),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4731));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226565 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1127),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4455),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4730));
 OR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226566 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1159));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_n_108));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4728));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226570 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4644),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4645),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4727));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4726));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4725));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4724));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4625),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4723));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226575 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_273),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4649),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4722));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4721));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226577 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1156),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1076),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4720));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4576),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4391),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4719));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4718));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4717));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226581 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4623),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4716));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4714));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4715));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226584 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2685),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4713));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4711));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4659),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4712));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226587 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4710));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226588 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4709));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4605),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4707));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226591 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4646),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4706));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226592 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4618),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4705));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226593 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4674),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1142),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2734),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4704));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4701));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4700));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4699));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4698));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4697));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4696));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226601 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1117),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4669),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4443),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4695));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226602 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1105),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4694));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226603 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4702));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4693),
    .Y(u6_n_109));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4693));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1157));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4691));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1156));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4690));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226619 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4689));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226620 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4664),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4687));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4686));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4666),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4685));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4476),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4684));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4667),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4683));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4670),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4682));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4665),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4681));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4663),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4680));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226628 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1133),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4692));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226629 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4668),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4688));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4679));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4678));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4677),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4676));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4677));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4675));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4674));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4670));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4599),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4668));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226638 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4667));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226639 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4636),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4666));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226640 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4638),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4665));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226641 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4639),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4664));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226642 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4663));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226643 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4598),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4673));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226644 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4672));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226645 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4466),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4671));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4635),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4565),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4669));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1155));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226650 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1154));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226651 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4662));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4660));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226654 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4661));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4659));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4657));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4656));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4622),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4654));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4653));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226662 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4620),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4652));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4651));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4650));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226665 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4640),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4491),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4658));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4649));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226669 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4612),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4575),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1148),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4500),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4648));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226670 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4615),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4498),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4647));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226671 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1112),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4614),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1113),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4499),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4646));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4645));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4644));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226674 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1152),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4643));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226675 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4584),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4642));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226677 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4641));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4634));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226683 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1104),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1147),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1109),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4496),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4632));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226684 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4495),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4631));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226685 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4612),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4630));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226686 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4444),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4629));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226687 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4607),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4640));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226688 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1149),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1153));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226689 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4608),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4639));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4638));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226691 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4636));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226692 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4635));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226693 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4633));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4513),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4628));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4505),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4627));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4626));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4625));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4624));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4623));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226702 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4457),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4622));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226703 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4616),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4445),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4621));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226704 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4450),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4620));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226705 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1113),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4619));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4615),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1112),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4618));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226708 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4454),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1152));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226709 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4590),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4617));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4614));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4613));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4612));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4610));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1150));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226719 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4608));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226722 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1149));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226723 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4557),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4478),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4606));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226724 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1151));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226725 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4519),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4616));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226726 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4525),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4615));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226727 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4567),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4611));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226728 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4578),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4568),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4609));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226729 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1143),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4607));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4605));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226731 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1118),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4604));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4603));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226734 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4581),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4398),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4418),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4602));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226735 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1145),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4601));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226736 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4600));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4599));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4598));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4597));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226740 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4549),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4437),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4596));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4536),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4595));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4535),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4594));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4593));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1148));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4591));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4537),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4474),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4589));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1139),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4521),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4588));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4522),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4587));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4518),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4586));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4592));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4547),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4515),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4590));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4472),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4583));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1147));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4566),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4479),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4585));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4496),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4469),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4584));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226759 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4464),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1146));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4581));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4580));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1145));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1144));
 AOI221x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226769 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1093),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4502),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4438),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4577));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4576));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4495),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1117),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1134),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4582));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4579));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4540),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4578));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1106),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1143));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4575));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4574));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4572));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226779 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4332),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1142));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226780 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4353),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4333),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4570));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4429),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1110),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1115),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4569));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1122),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4568));
 NAND3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4422),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4567));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4566));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4565));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4350),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4331),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4564));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1106),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4374),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4563));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4391),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4375),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4562));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226789 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4420),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4573));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1100),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2500),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4561));
 NOR3x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4458),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4571));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1099),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4560));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1101),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_660),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4559));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1101),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4558));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226795 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1093),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4557));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1100),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4556));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1137),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4555));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226798 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4554));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226799 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4552));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226800 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4550));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226802 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4548));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4546));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4419),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4545));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4446),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4430),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4433),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4544));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226808 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1128),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4543));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4440),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4542));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226810 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4394),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4541));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226811 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .A2(n_14488),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4540));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226812 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4401),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4539));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226813 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1114),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4400),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4553));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226814 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1101),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_820),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4538));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4551));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226816 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4451),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4549));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4417),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4397),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1141));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2779),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4537));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4431),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4547));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2770),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4536));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4535));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4454),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1140));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226823 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4427),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4399),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1139));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4534));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4532));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4530));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4528));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4524));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226835 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1078),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4523));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226836 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4533));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4531));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_619),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4522));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1081),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4379),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4521));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226840 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4389),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4520));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226841 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4529));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1083),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4519));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1082),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1138));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226844 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4518));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4517));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4443),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4516));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226847 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1096),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4515));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226848 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1079),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4514));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4513));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4512));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4436),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4465),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4527));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1137));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4511));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226854 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1097),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4510));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4509));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4468),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4508));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1090),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4507));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226858 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4525));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4450),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4506));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226860 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4456),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4505));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1088),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4504));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226862 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1088),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4503));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1136));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1135));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4502));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4501));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1134));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4499));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1078),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4494));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226873 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1078),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_26),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4493));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226874 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_14),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4361),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4492));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226875 (.A1(n_14150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4355),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1133));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226876 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4354),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4491));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226877 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_807),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1090),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4490));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4489));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226879 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1085),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4488));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226880 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1096),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1097),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4487));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1115),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4486));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226882 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_778),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1088),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4485));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4484));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4500));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226885 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1082),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4483));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226886 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_113),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1080),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4498));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226887 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4371),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4482));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1080),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_56),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4481));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4376),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4480));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4479));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4478));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4477));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4476));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226894 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1077),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4475));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226895 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1076),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4474));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4473));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226897 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4361),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4497));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226898 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_407),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .B2(n_14488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4472));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226899 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1076),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_731),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1077),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4471));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226900 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1083),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4470));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4496));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4495));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4469));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4468));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4466));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4465));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226910 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4462),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4463));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4461));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4459));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4458));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4457));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4453));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4449));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1125));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1124));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4445));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4444));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4443));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4440),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4441));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4439));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226942 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1120));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4436));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4435));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4434));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4467));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4433));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4432));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1132));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1131));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4464));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4462));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226957 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1130));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_34),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4460));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1129));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1128));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4456));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4455));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4454));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1127));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4451));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_167),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4450));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1126));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226968 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4447));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4431));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4446));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1123));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226972 (.A(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1122));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226973 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1121));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226974 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4442));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226975 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4430));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4429));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4440));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4438));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g226979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4389),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4437));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g226980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1119));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226981 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1118));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1117));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4427),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4428));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4426));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4425));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1113));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1112));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g226999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4423));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4421),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4422));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4419),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4420));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4417),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4418));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4416));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4414));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1105));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1101));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1102));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4411),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1103));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4410));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1099));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1100));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_380));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4408));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1116));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4407));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_113),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4406));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4405));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4404));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4403));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4402));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4427));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1115));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1114));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4424));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1111));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4401));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1110));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4400));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4399));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1109));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4421));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4419));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4417));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_40),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4398));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1108));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4397));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4383),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1107));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4415));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_26),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1106));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4395));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4394));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .B(n_14488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4393));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4412));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4392));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1104));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227065 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4295),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4360),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4411));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4359),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4311),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4409));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4391));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4389));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1097));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1096));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4385),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1095));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4385));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4386));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1093));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1090));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4384),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1091));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4382));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1089));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1088));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1087));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4380),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4379));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4335),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4358),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_407));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4388));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227116 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4304),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4351),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4387));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4312),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1094));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4315),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4345),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4384));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4383));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4316),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4381));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4310),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4380));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4378));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4374),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4375));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227125 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4374));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227127 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4371));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1086),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1085));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1086));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1083));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1082));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1084));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1080));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1079));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1081));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1078));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1077));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1076));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1075));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227173 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4289),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4360));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227174 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4292),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4346),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4359));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4335),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4376));
 NAND3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4335),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4373));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4372));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4368));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227179 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4365));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4349),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4363));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227181 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4319),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4336),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4361));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227183 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4308),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4356));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4355));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227185 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4354));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227186 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4353));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227187 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4352));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227188 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4254),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4329),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4351));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227189 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4350));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227190 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4275),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4349));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227191 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1028),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4274),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4290),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4348));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4330),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4347));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227193 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1072),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1074),
    .B(n_3634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4358));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227194 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4288),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4346));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227195 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4268),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4345));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227196 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4226),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4344));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227197 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4324),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4343));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227198 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4204),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4342));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227199 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4341));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227200 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4326),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4340));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4339));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227202 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4303),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4232),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4309),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4338));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227203 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4291),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4296),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4337));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227204 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1073),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4278),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4336));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227205 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1045),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4256),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4334));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_24),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4333));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4332));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4331));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4271),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4228),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4330));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227210 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4252),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4329));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227211 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_266),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4328));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227212 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1041),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4255),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4327));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227213 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4196),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4326));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227214 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_268),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4325));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227215 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4257),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4274),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4324));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4298),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4335));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227219 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4321));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227220 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4194),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4320));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4294),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4319));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4231),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4318));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227223 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4167),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4166),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4317));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4316));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227225 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4270),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4315));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4227),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4314));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227227 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4225),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4313));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4312));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4311));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227230 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4203),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4306),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4310));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4230),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4272),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4309));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4308),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4307));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4304));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227236 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1074));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4302),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1073));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3984),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4301));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227240 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4300));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227241 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4299));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227242 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2656),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4298));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4297));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227244 (.A(n_3635),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4296));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227245 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3898),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4308));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4281),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4306));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227247 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4305));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4271),
    .B(u6_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4303));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4271),
    .B(u6_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4302));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4088),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4295));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4294));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4262),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4293));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4292));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227254 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2729),
    .B(u6_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4291));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4290));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4266),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4289));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4261),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4288));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4287));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1072));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4283));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4286),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4282));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4286));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227267 (.A(u6_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4281));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227268 (.A(u6_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4279));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227269 (.A(u6_rem_96_22_Y_u6_div_90_17_n_182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4250),
    .Y(u6_n_111));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227270 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1065),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4278));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227271 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2807),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4277));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227273 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4275),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4274));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4275));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4272));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4271));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4236),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4270));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4237),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4269));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4238),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4268));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227281 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4239),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4267));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227282 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4180),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4222),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4058),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4266));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227283 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4052),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4243),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4265));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227284 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4036),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4245),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4264));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4136),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4161),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4263));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227286 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1055),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4262));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227287 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4261));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4273));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4121),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4260));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4233),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4259));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227291 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1070),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4258));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227292 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4235),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4257));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4246),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4256));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227294 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4234),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4255));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4244),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4254));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227296 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4253));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4242),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4252));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227298 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4205),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4251));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227299 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4174),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4250));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227300 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4187),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4229),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4249));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227301 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4223),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4163),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4248));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227302 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4221),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4173),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4247));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4246));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4243),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4244));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4242));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4240));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227308 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4216),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4079),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4075),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4238));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227309 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4217),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1057),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4237));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227310 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4206),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4236));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227311 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4235));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227312 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4234));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227313 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4219),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1056),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4233));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227314 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1067),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4211),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4245));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227315 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4215),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4138),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4243));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227316 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4210),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4241));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227317 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4206),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4176),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4239));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227318 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4216),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1071));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227321 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4093),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4232));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4201),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4095),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4231));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4091),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4230));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227325 (.A1(n_14530),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3921),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_4156),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_4190),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4229));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4213),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4228));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227327 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4115),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4227));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227328 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4226));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227329 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4217),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4097),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4225));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4140),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4206),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1070));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227331 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4224));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227332 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4078),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4199),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4223));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4222));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227334 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4070),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4221));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4220));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227338 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4216));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227339 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4215));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4213));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227341 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4211),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4212));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4211));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4041),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4161),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4109),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4209));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227344 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4049),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1065),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4108),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4208));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227345 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1068),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4219));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227346 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4182),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4218));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227347 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1069),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4217));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4181),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4214));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227349 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4182),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4210));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4206));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227352 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4204));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227353 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1069),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4203));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4202));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1069),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4020),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4201));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227357 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4182),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4030),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1054),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4200));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227358 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4184),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4205));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4171),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1055),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4199));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227360 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1066),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4198));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4196));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227363 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4195));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4165),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4194));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227365 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4124),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4193));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4130),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4159),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4192));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4191));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227368 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4157),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4190));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227369 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4177),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4189));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227370 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4175),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4135),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4188));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1067),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4187));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4086),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4186));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4092),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4185));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1069));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4129),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4184));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227381 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4034),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4182));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1068));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3994),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4181));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4180));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4178));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4176));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4173),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4174));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4172));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4056),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1057),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4019),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4170));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227394 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1056),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4022),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4169));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4032),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1049),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4029),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_4018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4168));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227396 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4021),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4037),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4167));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4038),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4166));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4133),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4179));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1054),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4017),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4177));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4165));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227401 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4132),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4175));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4164));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3996),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4163));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227404 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4025),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4173));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227405 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4076),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4066),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4171));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1067));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4160));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4158));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227412 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4155));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227413 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4031),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4011),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4153));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227414 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4033),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3992),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4152));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227415 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4009),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4151));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1051),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4150));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4059),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4149));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1062),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4148));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227419 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4055),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4147));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1060),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4064),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1066));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1029),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4161));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1029),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1065));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227423 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1053),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4159));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227424 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_4053),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3993),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4157));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_44),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4146));
 AND3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3997),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_4035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4156));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227427 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1050),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_4027),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4154));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227428 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4145));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227429 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4142));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4140));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4137),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4138));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4135),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4136));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3922),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4134));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227434 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4144));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4051),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4133));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4077),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1055),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4132));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227437 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1030),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_814),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4131));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227438 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4130));
 AO22x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227439 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4143));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227440 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1036),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_778),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4141));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227441 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2494),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4129));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227442 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3975),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4139));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227443 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_113),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4128));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227444 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4127));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4126));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227446 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1030),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4125));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227447 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1036),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4137));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227448 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4124));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227449 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4123));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4068),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4122));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227451 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3969),
    .A2(n_14146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4135));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4121));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4058),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4120));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227454 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_546),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4119));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227455 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4118));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227456 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3984),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4117));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4116));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4115));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3984),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4114));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4067),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4113));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1064),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4065),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4112));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3915),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4109));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227465 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4108));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227466 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1037),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4107));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227467 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2857),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1046),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4106));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227468 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3989),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4105));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227469 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1045),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4104));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227470 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_113),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4103));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227471 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4102));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4101));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1053),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4100));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4099));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227475 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1041),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_778),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4098));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227476 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4111));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227477 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4097));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227478 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3967),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4096));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227479 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1032),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4095));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227480 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1028),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4094));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227481 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4093));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227482 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3964),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4092));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227483 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1032),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4091));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227484 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3970),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4090));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227485 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_26),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4089));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227486 (.A1(n_14146),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1028),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4088));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227487 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_507),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4087));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227488 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3964),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4086));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227489 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_730),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4085));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227490 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4084));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227491 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3989),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_619),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4083));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4081));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4078));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1061));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4075));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4073),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4074));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4072),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4071));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4069),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4070));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4068));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4066),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4067));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4065));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1058),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4063));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4061),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4062));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4060));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4058));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4055),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4056));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4053),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4054));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4052));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4050));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4049));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4048));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4047));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4046));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4045));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4082));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1064));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4044));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4043));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4042));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1063));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1062));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4080));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4079));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4077));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4076));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3975),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1060));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4073));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4041));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4072));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4069));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1059));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4066));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4064));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1058));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1057));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4061));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4059));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1056));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4057));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4055));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4053));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4040));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4039));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4051));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1055));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4038));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4036));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227559 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4033),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4034));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4032));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4030));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4028));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4026));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4024));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4021));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4020));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4018));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4016));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227575 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4014));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4012));
 AOI31xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227578 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1023),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1024),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4010));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3961),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4009));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4008));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4007));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227582 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4006));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4004));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_26),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4037));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4003));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4002));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4001));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4000));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3999));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227591 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4035));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4033));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4031));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4029));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1054));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4027));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3998));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3997));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4025));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1029),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3996));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227601 (.A(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1053));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3995));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1052));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4022));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1051));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4019));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227607 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3994));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1050));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4017));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3993));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4015));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227612 (.A(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3992));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4013));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1049));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4011));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3991));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1048),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3989));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1046));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3988),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1047));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1044));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1045));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3984));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1043),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1042));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1043));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227644 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1041));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227646 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1040));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3981));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227648 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3982));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227656 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1039),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1038));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3976));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1037));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1036));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3951),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1048));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3988));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227669 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3934),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3891),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3987));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3985));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227671 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3980));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1039));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3975));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1035));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3973));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1033));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1032));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227699 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1031));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3970));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1028));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227709 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1029));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3966),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3968));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3967));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1027));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227720 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3964));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227727 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1025));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227728 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1026),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3963));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1026));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1023),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1024),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3962));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1034));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3972));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227733 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3906),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3934),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1030));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227735 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3950),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3966));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227736 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3942),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2521),
    .B2(u6_n_112),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3965));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3961),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1024));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227739 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3961));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227741 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3958));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227742 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3926),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3876),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3957));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227743 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3956));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227744 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3861),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3955));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227745 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2634),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3960));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227746 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3871),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_977),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3954));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3896),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3953));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3952));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227749 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3860),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3951));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3816),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3950));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227751 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3828),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3949));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3948));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227753 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3946));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3815),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3945));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3827),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3944));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227756 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3943));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227757 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .Y(u6_n_112));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227758 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3942));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3941));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227762 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3858),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3940));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227763 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3886),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3939));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227764 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3832),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3831),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3938));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3862),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3936));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2731),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1023));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3934));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3883),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3935));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3932));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3875),
    .B(u6_n_113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3933));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3894),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3876),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3931));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3876),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3897),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3930));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3929));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3901),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3928));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3899),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3753),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3927));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3926));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3925));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3922),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3923));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3921));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3918),
    .Y(u6_n_113));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227782 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2806),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3876),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2509),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3917));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3916));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .C(n_14150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3915));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227785 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3914));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(n_14150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3924));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227787 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3922));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3884),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3920));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3848),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3872),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3918));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227790 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3913));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3876),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3863),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3912));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3640),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3911));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3910));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227794 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3905),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3909));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227795 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3887),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3908));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227796 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3907));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3906));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227798 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3856),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3905));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3819),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3820),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3904));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3903));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3851),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3854),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3902));
 A2O1A1O1Ixp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3774),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3806),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3690),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1003),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3901));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3870),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_996),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3900));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227804 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1002),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3899));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3898));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3867),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3897));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3896));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3895));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3894));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227810 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3796),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3795),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3893));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3892));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3866),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3891));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3859),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3890));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227814 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3762),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3889));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3725),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3888));
 O2A1O1Ixp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227816 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3845),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_995),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3724),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3887));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3711),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1008),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3886));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3884));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3885));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3881));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3882));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227829 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3817),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3847),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3883));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3874),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3876));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3874));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227836 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3850),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3849),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3875));
 AOI31xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227837 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1019),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3761),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_3774),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3873));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227838 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3734),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3852),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3872));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227839 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3791),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3852),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3871));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227841 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1021),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3869));
 A2O1A1O1Ixp25_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227842 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3768),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1017),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3790),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3705),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3868));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227843 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3867));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227844 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3841),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1022));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227845 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3866));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227846 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3838),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1013),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3870));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1021),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3865));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3864));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3838),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3863));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3834),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3862));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3861));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3860));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227853 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3712),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3843),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1010),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3859));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3858));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227855 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3810),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3802),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3857));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3739),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3856));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3764),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3855));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227858 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3810),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_409),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3740),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3854));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227860 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_998),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3851));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227861 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1013),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3756),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3792),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3732),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3850));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3818),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3849));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3848));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227864 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3825),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3847));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227865 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1002),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3803),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1011),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3703),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3697),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3852));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227867 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3755),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3813),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1021));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227868 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1017),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3846));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3845));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227870 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3766),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3844));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3842),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3843));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3842));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3841));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227875 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3811),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3840));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227877 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3798),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3822),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3838));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3837));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1019));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227883 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3814),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3797),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1020));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227884 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1016),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3687),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1001),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3835));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227885 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3666),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1017),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3834));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1016),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3833));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3745),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3832));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3744),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1017),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3831));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3830));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3742),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3829));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3716),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3828));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3778),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3827));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227894 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3805),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3760),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3787),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3825));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227895 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3789),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3758),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3783),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3824));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227896 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1014),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3757),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3823));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227897 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3769),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3822));
 NAND5xp2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1002),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3733),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_1004),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_1009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3821));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227899 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2769),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3735),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3820));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227900 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2768),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_982),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3819));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227901 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3713),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_996),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3818));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3761),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3737),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3817));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227903 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3816));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2761),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3815));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227908 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1017));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227909 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1018));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227910 (.A(n_14489),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3779),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3814));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1016));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3812),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3813));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227914 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3812));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227915 (.A(n_14490),
    .B(n_13859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3811));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1015),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3810));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227919 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1015));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227920 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3808));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3806));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3804));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3801),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3802));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3801));
 NOR4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227927 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3707),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3685),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3799));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227928 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3769),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3798));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3767),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3702),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3797));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227930 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3676),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_982),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3796));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227931 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3643),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3645),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2769),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3795));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227932 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3635),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3616),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3794));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227933 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3699),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1005),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3793));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227934 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_997),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3792));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227935 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3691),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1007),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3696),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3805));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227936 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1001),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1014));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3803));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3662),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3800));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227939 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3773),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3703),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_1002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3791));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227941 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3790));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3610),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3788));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1003),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3787));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227945 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_195),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3785));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227946 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3617),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3784));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227947 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3701),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1006),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3783));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_982),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3781));
 AOI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227951 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3642),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3659),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3671),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3779));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1013));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3778));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_981),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_44),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3777));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227955 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3665),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1000),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3667),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3789));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3776));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3773));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227959 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3771));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3768));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1012),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3766));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3765));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3763));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3761));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227967 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3759));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227968 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3774));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1004),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3772));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227970 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_991),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3758));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_991),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3757));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227972 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3756));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227973 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_984),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3770));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227974 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3769));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227975 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3767));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227976 (.A(u6_rem_96_22_Y_u6_div_90_17_n_999),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3755));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227977 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_975),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1012));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227978 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3754));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3753));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227980 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3752));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3751));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3750));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1008),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3764));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3749));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227985 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3748));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227986 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_984),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3762));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3747));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227988 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3746));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g227989 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3760));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3745));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3743));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3741));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227993 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3739));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3735),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3736));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3733),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3734));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g227996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3731),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3732));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g227999 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2768),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3728));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228000 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2857),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3727));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228001 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_984),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3726));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_195),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3725));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228003 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_195),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_983),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3724));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228004 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3640),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3723));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228005 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3744));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228006 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_37),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3722));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228007 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_596),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_973),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3721));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228008 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3689),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3720));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_998),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3742));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228010 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_981),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3719));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228011 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_981),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3718));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228012 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_973),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3740));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3738));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228014 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3717));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228015 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_979),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3716));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228016 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_979),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3715));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3737));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228018 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_977),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3714));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228019 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_979),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3735));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228020 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3733));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228021 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3731));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228024 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1009),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3712));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1007),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1008));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3711));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3709));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3708));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3706));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3705));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3702));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3700));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3698));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3697));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3696));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3695));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3694));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3693));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_993),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3713));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1011));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1010));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1009));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1007));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3710));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3692));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1006));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3707));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228057 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1005));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228058 (.A(u6_rem_96_22_Y_u6_div_90_17_n_63),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3691));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3704));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1004));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3703));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228062 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3701));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3699));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228064 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3690));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1003));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1002));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3689));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3687));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_999),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3685));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3683));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3681));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_998),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3680));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228078 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3679),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_998));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3676),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3678));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3675));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_995),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3673));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_995));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3688));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3671));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_28),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_977),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3670));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3668));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3667));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228094 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1001));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228095 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3666));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1000));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228097 (.A(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3686));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3665));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228099 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_999));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3682));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228103 (.A(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3679));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228106 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3662));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228107 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2857),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_997));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3676));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228110 (.A(u6_rem_96_22_Y_u6_div_90_17_n_799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_996));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228111 (.A(u6_rem_96_22_Y_u6_div_90_17_n_784),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3660));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3674));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3659));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228114 (.A(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3672));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_993));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228129 (.A(u6_rem_96_22_Y_u6_div_90_17_n_992),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_991));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_989),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3651));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228139 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_989));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_987),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_986));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_985),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_984));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228169 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_983));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228171 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3602),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_139));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_992));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228173 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3605),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3652));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3601),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_987));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228175 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3626),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_985));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3646));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3645));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228182 (.A(u6_rem_96_22_Y_u6_div_90_17_n_981),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3643));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_981));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3642));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_979));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_977));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_976),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3640));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_976));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_973));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228224 (.A1(n_3638),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_982));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228225 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2460),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3619),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3644));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3622),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_980));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228227 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3568),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_978));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3599),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_975));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228229 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3600),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_974));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228230 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3581),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3637));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228231 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3636));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228232 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_200),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3635));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228233 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3594),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3634));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3594),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3579),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2654),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3633));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228235 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3632));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228236 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3631));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228237 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_260),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3630));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228238 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3629));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228239 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3582),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3626));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228240 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3625));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228241 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3624));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228242 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_264),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3611),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3623));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3578),
    .A2(n_3639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3593),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3622));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3570),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_930),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3621));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3628));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228246 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3627));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228248 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_939),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3618));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_971),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3617));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228250 (.A(u6_rem_96_22_Y_u6_div_90_17_n_200),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3616));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2595),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3615));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228252 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3614));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228253 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3613));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228254 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_944),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3577),
    .B(n_14534),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3612));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228255 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3611));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228256 (.A(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3610));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3619));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3569),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3609));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228259 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_932),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3608));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228260 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_935),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3607));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3526),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3606));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3605));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228263 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_937),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3604));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228264 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3549),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3603));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3567),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3602));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228266 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3601));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228267 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3600));
 NAND2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3513),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3599));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_972),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_971));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3598));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228282 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3594));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3576),
    .B(u6_n_115),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3593));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3592));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228285 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3525),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3591));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228286 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3502),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3503),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3590));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228287 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2654),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3589));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228288 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3338),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_972));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228289 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3596));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228290 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3571),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3595));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228291 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3544),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3543),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3588));
 OA21x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228292 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2803),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2800),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3587));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3586));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228294 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3515),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3516),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3585));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228296 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3546),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3583));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3582));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3472),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3581));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3579));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228300 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3578));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228304 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3577));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228305 (.A(u6_rem_96_22_Y_u6_div_90_17_n_738),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3580));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228306 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3499),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3532),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3558),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2792),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3576));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3575));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228308 (.A(u6_rem_96_22_Y_u6_div_90_17_n_876),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3574));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228309 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3572),
    .Y(u6_n_115));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3572));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228311 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3541),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3514),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3538),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2796),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3571));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228312 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3485),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_970),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3495),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3428),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3570));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228313 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3451),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3569));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228314 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3568));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228315 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3554),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3473),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3567));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3556),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3453),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3566));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228317 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3552),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3452),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3565));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228318 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3498),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3530),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3564));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228319 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3488),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3563));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228320 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3542),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3419),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_960),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3562));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228321 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3421),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_970),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3561));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3450),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3560));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228325 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3339),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3537),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3559));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3558));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228327 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3349),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3534),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3557));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228328 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3402),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3529),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3556));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228329 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3474),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3555));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228330 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3532),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_955),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3554));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228331 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3422),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3438),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3553));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228332 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3387),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3408),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3552));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3533),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3551));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228334 (.A(u6_rem_96_22_Y_u6_div_90_17_n_969),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3550));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228335 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3527),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3549));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228337 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_965),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3518),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3547));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228338 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3509),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3519),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3546));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228340 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3414),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3411),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3459),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3544));
 AOI211xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228341 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_965),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3413),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3458),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3543));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228343 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_961),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3542));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228346 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_970));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228347 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_967),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3505),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3541));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228348 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3433),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3434),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3540));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_968),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3539));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228350 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3443),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3494),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3487),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2686),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3538));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228351 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3476),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3439),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3429),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3347),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3537));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228353 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_965),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3478),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3535));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228355 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_966),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3481),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_969));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228356 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3435),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_962),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3427),
    .C(n_13863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3534));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3533));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228358 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3532));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3531));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228361 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3512),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3506),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3530));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3529));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228363 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3510),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3528));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228364 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_966),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_958),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3527));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_966),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3468),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3526));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228366 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3464),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3525));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3465),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3524));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228369 (.A(u6_rem_96_22_Y_u6_div_90_17_n_967),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_968));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228371 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3396),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3395),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_967));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3486),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3523));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3522));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228374 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3483),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3496),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3491),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3521));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_963),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3482),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3520));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228376 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3519));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228377 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3518));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228378 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3507),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3479),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3517));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228379 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3406),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3444),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3516));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228380 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3417),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_948),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_950),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3456),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3515));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3484),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3504),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3514));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228382 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3447),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2595),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3513));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228385 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3512),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_966));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228386 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3390),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3457),
    .B(n_13861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3512));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3511));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_965));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228391 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_951),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3455),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3510));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_964),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3509));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3508));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3480),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3506));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3477),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3479),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_964));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228398 (.A(u6_rem_96_22_Y_u6_div_90_17_n_961),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3505));
 AOI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228399 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_929),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(n_13864),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3504));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_949),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_951),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3503));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228401 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_950),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3406),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3502));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228402 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3418),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_960),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3501));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228404 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_959),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3392),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_963));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228405 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3409),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3388),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3397),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3507));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3498),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3499));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228407 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3496),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3497));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3495));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228411 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3420),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3437),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3425),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3491));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228412 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3385),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3407),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3490));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228413 (.A(u6_rem_96_22_Y_u6_div_90_17_n_953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3436),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_955),
    .D(n_13862),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3498));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228414 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3405),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_948),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3489));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3440),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3401),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3359),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3488));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228416 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_929),
    .A2(n_13864),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3348),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3487));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228417 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3415),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3496));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228418 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_953),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_956),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_962));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228419 (.A(u6_rem_96_22_Y_u6_div_90_17_n_931),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3486));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228420 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3426),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3494));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228421 (.A(u6_rem_96_22_Y_u6_div_90_17_n_933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3492));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3485));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3481));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228425 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3478));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228426 (.A(u6_rem_96_22_Y_u6_div_90_17_n_952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3476));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228427 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_946),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3484));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228428 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3374),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3382),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3483));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228429 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3374),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3382),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3482));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3480));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228431 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_43),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_938),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_961));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228432 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_930),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3475));
 AO22x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228433 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3479));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228434 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3412),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3389),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3477));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228435 (.A(u6_rem_96_22_Y_u6_div_90_17_n_953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3474));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3442),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3473));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228437 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_946),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3472));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228438 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_944),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3471));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228439 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_602),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_944),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3470));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3434),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3469));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228441 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_941),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3468));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3431),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_955),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3467));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228443 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_943),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3466));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228444 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3465));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228446 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3461));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228447 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3458),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3459));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228448 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3457));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228449 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2765),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3456));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228450 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3455));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228451 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_938),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_602),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3454));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228452 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_946),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3453));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228453 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_941),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3464));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228454 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3462));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228455 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_943),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_784),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3460));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228456 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3375),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3452));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228457 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_939),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3375),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3451));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228458 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_938),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3450));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_931),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_932),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3449));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228460 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3375),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3448));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228461 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_931),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3447));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228462 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_938),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_937),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3458));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228463 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_934),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3446));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228464 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_934),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_935),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3445));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228465 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_934),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_935),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3444));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228466 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_929),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(n_13864),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3443));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3441),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3442));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3439),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3440));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3437),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3438));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3435),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3436));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_959),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3434));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3432),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3433));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3431));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3429));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3428));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3441));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3439));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3427));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3426));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3425));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3424));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3423));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3422));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3437));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_960));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3435));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_959));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_941),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3432));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_958));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_957));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_956));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3421));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_955));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_954));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_953));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3420));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3419));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3418));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3416),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3417));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3414));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3412),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3413));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228514 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3410),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3411));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3409),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3410));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3407),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3408));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3406));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_949),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_950));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3405),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_949));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3404));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3402));
 NOR2x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3416));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3400));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3399));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3398));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3397));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3396));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3395));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228538 (.A(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3393));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3392));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3415));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3412));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3409));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_952));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228545 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3390));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3407));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228547 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3389));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_759),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3388));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_951));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3405));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228551 (.A(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3387));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_784),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3403));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_784),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3401));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_948));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3385));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_947),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_946));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3383),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_947));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228566 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3331),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3368),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3383));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_944));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3382),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_945));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3381),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3382));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228579 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3301),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3367),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3381));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_942));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3379),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_943));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228589 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3316),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_927),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3366),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3379));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_941));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3378),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_940));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3378));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3355),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3365),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3377));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228600 (.A(u6_rem_96_22_Y_u6_div_90_17_n_939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3375));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228605 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_939));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3376),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3374));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3364),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3356),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3376));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_937));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3373),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_938));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3354),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3362),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3373));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_934),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_935));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228624 (.A(u6_rem_96_22_Y_u6_div_90_17_n_936),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_934));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3372),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_936));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228627 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3358),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3363),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3372));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_932));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_931));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3371),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_933));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228636 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2464),
    .A2(u6_n_116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3369),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3371));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228640 (.A(u6_rem_96_22_Y_u6_div_90_17_n_929),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_930));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3370),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_929));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228643 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3319),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3370));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228644 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2579),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2562),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3350),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3369));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228645 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3345),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3357),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3368));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_263),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3328),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3302),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_3323),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3367));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228647 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3321),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3344),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3366));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228648 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3343),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3365));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3320),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3342),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3364));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2727),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3341),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3363));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3352),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3297),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3362));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3176),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_927),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3312),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3361));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3323),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .Y(u6_n_116));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228656 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_234),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_806),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3359));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228657 (.A(n_14535),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3358));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228658 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3329),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3330),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3194),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3357));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3313),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3356));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228660 (.A(n_14292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3355));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228661 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3298),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3354));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3352),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_927));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3350));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3349));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3348));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228669 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_924),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3347));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3336),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3352));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3329),
    .B(u6_n_117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_926));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3271),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3345));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228675 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_906),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3334),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3344));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228676 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_900),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3335),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3343));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228677 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3332),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3342));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228678 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3329),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2804),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2507),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3341));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228679 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3333),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3340));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228680 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3325),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_806),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3339));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228681 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3338));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228682 (.A(u6_n_117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3336));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228683 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3310),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3241),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3286),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2796),
    .Y(u6_n_117));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228684 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3275),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3276),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3335));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3334));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228686 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3288),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3287),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3333));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3315),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3328),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3332));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228688 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3317),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3273),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3331));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3318),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3272),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3330));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228690 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3311),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3329));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228691 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3269),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3311),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3328));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3325),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_924));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3325));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_925),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3323));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3327),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_925));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228703 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3305),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3240),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3261),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3327));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228704 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_915),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3223),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3322));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228705 (.A(u6_rem_96_22_Y_u6_div_90_17_n_923),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3321));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3309),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3238),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3320));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228707 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_921),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3292),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3296),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3208),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3319));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228708 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3206),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_912),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3318));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228709 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3215),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3225),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3317));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228710 (.A(u6_rem_96_22_Y_u6_div_90_17_n_922),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3316));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3303),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3236),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3315));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228712 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3308),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3237),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3314));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3313));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3306),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3233),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3312));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228715 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3289),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3282),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3293),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3311));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228717 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3249),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3300),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_923));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228718 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3299),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3310));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228719 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_917),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3309));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228721 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3307),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3308));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228722 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3283),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3252),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_919),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3307));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228724 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_920),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3258),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3268),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_922));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3305),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3306));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228726 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3290),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3294),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3305));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228727 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_920),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3304));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228728 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_914),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3283),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3303));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3284),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3234),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3302));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228730 (.A(u6_rem_96_22_Y_u6_div_90_17_n_920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3301));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228733 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3300),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_921));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3299),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3300));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228735 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3192),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3263),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3299));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3264),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3235),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3298));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3239),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3260),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3297));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228738 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3295),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3296));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228739 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3270),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3265),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3278),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3295));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228740 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3277),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3267),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3280),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3294));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228741 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3274),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3279),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3293));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3292));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3277),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3290));
 NOR4xp75_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3256),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_915),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3219),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3291));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_914),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3205),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3228),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3289));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3259),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3200),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3288));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228747 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3211),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3254),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3287));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3162),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3207),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3163),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3286));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228750 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3285),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_920));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3283),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3284));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228752 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3282),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3283));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228754 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3243),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3224),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3280));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228755 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_912),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3229),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3231),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3279));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228757 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3255),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3222),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3278));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228758 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3213),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3253),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3262),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3285));
 AOI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228759 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3198),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3201),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2781),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3187),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_913),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3282));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3203),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3276));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228761 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3204),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3202),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3275));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228762 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_906),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_32),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3274));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228763 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3194),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3273));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228764 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3277));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_32),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3194),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3272));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228766 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3194),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3271));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3255),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3270));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3267),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3268));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3265),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3266));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3263),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3264));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3176),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3172),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3164),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3269));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228773 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3188),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3214),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3262));
 A2O1A1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228774 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3173),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3165),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2712),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3261));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228775 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_918),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3212),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3217),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3267));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228776 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3226),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3218),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3265));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228777 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3196),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_919));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228778 (.A(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3260));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_900),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_728),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2780),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3259));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .C(n_14536),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3263));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3258));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228782 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3256));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2781),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3254));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228784 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3180),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3253));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228785 (.A1(n_14291),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3252));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228786 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3251));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228787 (.A(n_14134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3250));
 OAI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228788 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_903),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_910),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_43),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3257));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228789 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3249));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228790 (.A(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3248));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228791 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3247));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228792 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_43),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3246));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228793 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_906),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3245));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3223),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3244));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3255));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228796 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .B(n_14134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3243));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228797 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3242));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228798 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3175),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3241));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228799 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3174),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3240));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228800 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3180),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3239));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228801 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_43),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_901),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3238));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228802 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_191),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_906),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3237));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228803 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_901),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_759),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3236));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228804 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3180),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3235));
 AOI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228805 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_31),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3234));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228806 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3176),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3233));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228807 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_901),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3232));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3231));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228809 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_900),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3230));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3229));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_32),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3228));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3226),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3227));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228814 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3224),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3225));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228815 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3222),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3223));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_916),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_915));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228821 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3221));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228822 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3219));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228823 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3217));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228824 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3226));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3216));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_918));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3224));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3215));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3222));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_917));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3214));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3213));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228833 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_916));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3212));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_914));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_31),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3220));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228837 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3218));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3211));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3207),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3208));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3205),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3206));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3204));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3203));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3202));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3200));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3197));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3194));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_911));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228861 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3209));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228862 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3193));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3192));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228864 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3191));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228865 (.A(n_14134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3207));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228866 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3190));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3189));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_191),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3205));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_913));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3188));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228871 (.A(u6_rem_96_22_Y_u6_div_90_17_n_728),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3201));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228872 (.A(u6_rem_96_22_Y_u6_div_90_17_n_730),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3198));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228873 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3187));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_912));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228875 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3196));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228876 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3137),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3195));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3185));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228883 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_908));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_907));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228888 (.A(u6_rem_96_22_Y_u6_div_90_17_n_910),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_909));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_910));
 OA211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228890 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_261),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3158),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3186));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_904),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_906));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_904));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228901 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3134),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3184));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_901),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_902));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228913 (.A(u6_rem_96_22_Y_u6_div_90_17_n_903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_901));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228915 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_903));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228916 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3119),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3167),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3182));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3180));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3160),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3181));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_900));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228926 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_899));
 OA22x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228927 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2639),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3161),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2520),
    .B2(u6_n_118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3179));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228928 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3145),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3178));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3177));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228936 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3130),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3153),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3176));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228937 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3175));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228938 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3174));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228939 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3173));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228940 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3151),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3172));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228941 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3150),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2907),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3171));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_897),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2732),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3170));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_897),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3127),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3169));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228944 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_886),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3168));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228945 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3167));
 AOI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228946 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3138),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_897),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_880),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3166));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228948 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3165));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_780),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3164));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228950 (.A(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3163));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3162));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228952 (.A(u6_rem_96_22_Y_u6_div_90_17_n_895),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .Y(u6_n_118));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228953 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3140),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3153),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3161));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228954 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2642),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3160));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228955 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2805),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3159));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228956 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_895),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3158));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228957 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3133),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_889),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3157));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228958 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3115),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3156));
 OAI22xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228959 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3118),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3155));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3153));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3154));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228963 (.A(u6_n_119),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_897));
 NAND2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3152));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3151));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228967 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3149));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228970 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3149),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_234));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228979 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3150));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3018),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3148));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3110),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3109),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3139),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3147));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228982 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3135),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3083),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3146));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228983 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3078),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3145));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228985 (.A(u6_n_119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3144));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3143),
    .Y(u6_n_119));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228987 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3121),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3086),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3100),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3143));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3141));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3140));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_895));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228993 (.A(n_14269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3142));
 AO21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228994 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3120),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3129),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3006),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3139));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g228995 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3131),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3080),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3138));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3079),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3137));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g228997 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3066),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3122),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_891),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3136));
 AOI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228998 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3125),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3075),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_890),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3135));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g228999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3123),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3134));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3092),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3133));
 OAI31xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229001 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3113),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_892),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_3097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3132));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229002 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_892),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_894),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3131));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229003 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_893),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3057),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3130));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3102),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3129));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229005 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3114),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3077),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3128));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229006 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3114),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3089),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3127));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229007 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3126));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229008 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3111),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3061),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3125));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229009 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3096),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3124));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229010 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3123));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229011 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2600),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3073),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3070),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3056),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3064),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3122));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229012 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3098),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3094),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3105),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3121));
 A2O1A1O1Ixp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229013 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3054),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3058),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3088),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_3085),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3120));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3108),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3082),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3119));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229015 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3112),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3084),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3118));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3107),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3081),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3117));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229017 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3099),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3095),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3116));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3091),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3115));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3114));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229023 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3113),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_894));
 AOI321xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229024 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3067),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3065),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2785),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3069),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3065),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3059),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3113));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3112));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229026 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3071),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3072),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3110));
 OAI221xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229027 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3046),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_100),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2744),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3109));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3043),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_631),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3108));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3047),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3111));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3107));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3106));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3104));
 NOR3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229034 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3087),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3055),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3102));
 AOI222xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229035 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_887),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_3051),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .C1(u6_rem_96_22_Y_u6_div_90_17_n_3041),
    .C2(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3105));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229036 (.A(u6_rem_96_22_Y_u6_div_90_17_n_891),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_893));
 O2A1O1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229037 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3033),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_3032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3101));
 AOI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229038 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_880),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3031),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3030),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3100));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229039 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3053),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3076),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3062),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3103));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3098),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3099));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3097));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3094),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3095));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229044 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3052),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_892));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229045 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3048),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3098));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229046 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_631),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3046),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3093));
 AOI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229047 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_889),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_31),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3092));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229048 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3046),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3091));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229049 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_889),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3090));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229050 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_889),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3089));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229051 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3032),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3096));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229052 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3048),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3094));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3087),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3088));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229054 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_880),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3031),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3086));
 OAI31xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229055 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3040),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3029),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_191),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3027),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3085));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229056 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_737),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_881),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_736),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3084));
 AOI22xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229057 (.A1(n_14291),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_886),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3083));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229058 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_881),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3082));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229059 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_631),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3081));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229060 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3038),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3080));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229061 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_886),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3079));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229062 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3039),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3087));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229063 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_885),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3078));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3076),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3077));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229066 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3074),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3075));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3045),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3073));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229068 (.A(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3072));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_100),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3071));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229070 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3070));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_41),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_891));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229072 (.A(u6_rem_96_22_Y_u6_div_90_17_n_86),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3069));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229073 (.A(u6_rem_96_22_Y_u6_div_90_17_n_889),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3068));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3076));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3067));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229076 (.A(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3066));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_31),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3074));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3063),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3064));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3062));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229081 (.A(u6_rem_96_22_Y_u6_div_90_17_n_737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3061));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_737),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3060));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229083 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3059));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229084 (.A(n_14291),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3058));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3038),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3057));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_890));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3056));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229088 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3041),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3065));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229089 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3055));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229090 (.A(u6_rem_96_22_Y_u6_div_90_17_n_887),
    .B(n_14291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3054));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2488),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_884),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3063));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3053));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_888),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_889));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3052),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_888));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3051),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3052));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3050),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3051));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229105 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3022),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2988),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3036),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3050));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_886));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_885));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_887));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229116 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3022),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2994),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3035),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3049));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229117 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3048));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3046));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229119 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3044),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3043));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229120 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3045),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3044));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3042),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3045));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229122 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3047),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3042));
 OAI22x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229123 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2633),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3026),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2468),
    .B2(u6_n_120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3047));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229132 (.A(u6_rem_96_22_Y_u6_div_90_17_n_883),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_881));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229133 (.A(u6_rem_96_22_Y_u6_div_90_17_n_882),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_883));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229134 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_882));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3041),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_884));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229136 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2730),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3022),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3037),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3041));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229137 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3039));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229138 (.A(u6_rem_96_22_Y_u6_div_90_17_n_880),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3038));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3040),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_880));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229144 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3021),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3009),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3034),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3040));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229145 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2636),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3025),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3037));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229146 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2987),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3024),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3036));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229147 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3020),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2995),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3023),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3035));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229148 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3007),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3019),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_853),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3034));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3033));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3018),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3032));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3031));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229152 (.A(u6_rem_96_22_Y_u6_div_90_17_n_877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_845),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3030));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229153 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3028),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3029));
 NAND2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_32),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3028));
 OR3x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_877),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_845),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_32),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3027));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3015),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3020),
    .Y(u6_n_120));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3014),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3019),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3026));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229159 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3010),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3025));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229160 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2986),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3010),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_857),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3024));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229161 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2993),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3010),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_856),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3023));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3022),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3021));
 NAND2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3012),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3022));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3020),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3019));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3010),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3020));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_878),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3018));
 OR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229172 (.A(u6_rem_96_22_Y_u6_div_90_17_n_845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_878));
 OAI32xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229173 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_3004),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_2985),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_494),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_788),
    .Y(u6_n_124));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229174 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3015));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3014),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_877));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3016),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3014));
 NOR2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2943),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3008),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3016));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229180 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3011),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3012));
 O2A1O1Ixp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229181 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2998),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2964),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2967),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3011));
 OAI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229182 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2992),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2983),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3010));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229183 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3001),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3009));
 AOI21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229184 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_3000),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2963),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2968),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3008));
 A2O1A1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229185 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_869),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2962),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3007));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3005),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3006));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229187 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2912),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3005));
 OR5x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229188 (.A(u6_rem_96_22_Y_u6_div_90_17_n_870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2966),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2849),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_733),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3004));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3002),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3003));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_835),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3002));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3000),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3001));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229192 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2961),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2980),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2956),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3000));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_876),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2999));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229196 (.A(u6_rem_96_22_Y_u6_div_90_17_n_218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_876));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_875),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_218));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229200 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2989),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_875));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229201 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_868),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2978),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_869),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2998));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2997),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2996));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229203 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2985),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2997));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2979),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2973),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2995));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229205 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2981),
    .B(n_14289),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2994));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2965),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2993));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229207 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2958),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2982),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2992));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2991),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2990));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_871),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2991));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229210 (.A(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_870),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_855),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2989));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2977),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2988));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2976),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2987));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2975),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2747),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2986));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2984),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2985));
 NOR2x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229215 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2984));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229216 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2955),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2941),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2937),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2983));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2957),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2969),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2982));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229218 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2980),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2981));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2980));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2954),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_874));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229222 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2978),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2979));
 MAJIxp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229223 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2952),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2978));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_872));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_220),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_871));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229241 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_857),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_86),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2953),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2977));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229242 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_857),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2953),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2976));
 OAI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229243 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2953),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_100),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2975));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229244 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_854),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2974));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229245 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_86),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_856),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2488),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2973));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2970),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2971));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229249 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2940),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2935),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2969));
 OAI21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229250 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2941),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2939),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2968));
 AOI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229251 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2942),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_41),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2938),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2967));
 OR3x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_855),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2912),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2559),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2966));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229253 (.A(u6_rem_96_22_Y_u6_div_90_17_n_126),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_870));
 OAI22xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229254 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_737),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_856),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2965));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229255 (.A(u6_rem_96_22_Y_u6_div_90_17_n_858),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2970));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229258 (.A(u6_rem_96_22_Y_u6_div_90_17_n_51),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2964));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2941),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2963));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229260 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2962));
 NOR2xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229261 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_869));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229262 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2487),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_868));
 NOR2xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_51),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2961));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_138));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229276 (.A(u6_rem_96_22_Y_u6_div_90_17_n_867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_866));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_15),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_867));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229283 (.A(u6_rem_96_22_Y_u6_div_90_17_n_248),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_15));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229297 (.A(u6_rem_96_22_Y_u6_div_90_17_n_863),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2960));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229306 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_863));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229310 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_864));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229324 (.A(u6_rem_96_22_Y_u6_div_90_17_n_216),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_865));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229343 (.A(u6_rem_96_22_Y_u6_div_90_17_n_215),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_860));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229345 (.A(u6_rem_96_22_Y_u6_div_90_17_n_136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_215));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_136));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229350 (.A(u6_rem_96_22_Y_u6_div_90_17_n_214),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_859));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_861),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_214));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_861));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229359 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_710),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2933),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2959));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229360 (.A(u6_rem_96_22_Y_u6_div_90_17_n_103),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2958));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229361 (.A(u6_rem_96_22_Y_u6_div_90_17_n_736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2957));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229362 (.A(u6_rem_96_22_Y_u6_div_90_17_n_51),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2956));
 OAI21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229363 (.A1(n_14164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2934),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_248));
 XNOR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2934),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_216));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2936),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2614),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_858));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229366 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_31),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2955));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_857),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2953));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2952),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_857));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229373 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2954),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2952));
 OAI22x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229374 (.A1(n_14492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2927),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_587),
    .B2(u6_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2954));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229375 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2951));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2945),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_856));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229383 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2944),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2945));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229384 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2929),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2931),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2944));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229385 (.A1(n_14130),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_845),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2943));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_846),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2930),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_855));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_853));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_854));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229392 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2942),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2941));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2940),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2942));
 AOI211x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229394 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2915),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2919),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2922),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2940));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2939));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229396 (.A(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2938));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229397 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2937));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229398 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2558),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2936));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2924),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2935));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2933),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2934));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_852));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229417 (.A(u6_rem_96_22_Y_u6_div_90_17_n_239),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_851));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_239));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_848));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_847));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_850),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_849));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_850));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229484 (.A(u6_rem_96_22_Y_u6_div_90_17_n_846),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2932));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229485 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2637),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2920),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_844),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2914),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2931));
 NOR3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2930));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229487 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2917),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2893),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2929));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229488 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2678),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2908),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2933));
 XOR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2913),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2667),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_247));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2909),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2668),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_846));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229491 (.A(u6_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2927));
 NOR2x1p5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2917),
    .Y(u6_n_122));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2926),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_845));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_791),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2924));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2918),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2926));
 NOR2xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_790),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2923));
 NOR2xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2882),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2921),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2922));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2920),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2921));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2889),
    .B(u6_n_123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2920));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2919));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2918));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2917),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_844));
 AO211x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229509 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_791),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2892),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2827),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2902),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2917));
 O2A1O1Ixp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229510 (.A1(n_13865),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2891),
    .C(u6_n_123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2915));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2735),
    .B(u6_n_123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2914));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229512 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2535),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2913));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2856),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2912));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_840),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2911));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2911),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_135));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_213),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_840));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229556 (.A(u6_rem_96_22_Y_u6_div_90_17_n_134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_213));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229573 (.A(u6_rem_96_22_Y_u6_div_90_17_n_394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_134));
 XNOR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2666),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_394));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2910));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_133),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_837));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_133));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229602 (.A(u6_rem_96_22_Y_u6_div_90_17_n_131),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_836));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229604 (.A(u6_rem_96_22_Y_u6_div_90_17_n_132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_131));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_132));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229610 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_838));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_835));
 XOR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2901),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_839));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2908),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2909));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229633 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2681),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_833),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2682),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2908));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229634 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2906),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2907));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229635 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2881),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2906));
 OA21x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229637 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2903),
    .Y(u6_n_123));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229638 (.A1(n_14491),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2872),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2903));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229639 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2890),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2873),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_51),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2902));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229640 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_695),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_826),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2901));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_834),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2900));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2894),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_834));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229645 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2680),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_826),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_833));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229659 (.A(u6_rem_96_22_Y_u6_div_90_17_n_129),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_830));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_129));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_130));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229679 (.A(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_8));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229691 (.A(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_831));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229694 (.A(u6_rem_96_22_Y_u6_div_90_17_n_127),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_9));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_832),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_127));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229698 (.A(u6_rem_96_22_Y_u6_div_90_17_n_126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_832));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229700 (.A(u6_rem_96_22_Y_u6_div_90_17_n_826),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2665),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_126));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229706 (.A(u6_rem_96_22_Y_u6_div_90_17_n_828),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_827));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_212),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_828));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229713 (.A(u6_rem_96_22_Y_u6_div_90_17_n_210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_212));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229717 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2897),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_210));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229718 (.A(u6_rem_96_22_Y_u6_div_90_17_n_125),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2897));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229732 (.A(u6_rem_96_22_Y_u6_div_90_17_n_829),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_125));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229736 (.A(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_829));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_246),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_14));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229744 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2888),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2617),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_246));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229745 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2895),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2896));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229746 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2895));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229747 (.A(u6_rem_96_22_Y_u6_div_90_17_n_805),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2894));
 AOI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229748 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_791),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_736),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2878),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2893));
 NAND3xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2890),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2873),
    .C(u5_mul_69_18_n_89),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2892));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229750 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2875),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2874),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2891));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2879),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2890));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229752 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_103),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_792),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2889));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229753 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_690),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2869),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2525),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2888));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229756 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_810),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2676),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_826));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229764 (.A(u6_rem_96_22_Y_u6_div_90_17_n_823),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_822));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229766 (.A(u6_rem_96_22_Y_u6_div_90_17_n_209),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_823));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229779 (.A(u6_rem_96_22_Y_u6_div_90_17_n_824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_209));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229780 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_824));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229781 (.A(u6_rem_96_22_Y_u6_div_90_17_n_825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2886));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_821),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_825));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_821));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_820),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_124));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_810),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2664),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_820));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_207));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229835 (.A(u6_rem_96_22_Y_u6_div_90_17_n_123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_816));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_123));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2885));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_122),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_11));
 XOR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229865 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2870),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_122));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229867 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_814));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_204),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_813));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229884 (.A(u6_rem_96_22_Y_u6_div_90_17_n_38),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_204));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_38));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_811),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_121));
 XNOR2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229920 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2871),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_811));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229921 (.A(u6_rem_96_22_Y_u6_div_90_17_n_789),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_712),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2882));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_799),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2881));
 AOI32xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229924 (.A1(n_3646),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2851),
    .A3(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .B1(n_3645),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2879));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229925 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2877),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2878));
 AOI221xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229926 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2853),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_100),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2757),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2718),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2849),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2877));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229928 (.A(n_14178),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_790),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2875));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2873),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2874));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229930 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2853),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2483),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2873));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229931 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2872));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229932 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2534),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2871));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229933 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_786),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_257),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2870));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229934 (.A(u6_rem_96_22_Y_u6_div_90_17_n_810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2869));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229937 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_810));
 INVxp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229938 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_37));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229943 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2865));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229944 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2864));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229956 (.A(u6_rem_96_22_Y_u6_div_90_17_n_808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_35));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229966 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_808));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g229969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_36));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229977 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2866));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2868),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_807));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g229992 (.A(u6_rem_96_22_Y_u6_div_90_17_n_203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2868));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_203),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_806));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g229996 (.A(u6_rem_96_22_Y_u6_div_90_17_n_786),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_203));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_202),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_801));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_800),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_202));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_120),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_800));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230029 (.A(u6_rem_96_22_Y_u6_div_90_17_n_119),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_120));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_119));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_201),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_803));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_256),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_201));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230065 (.A(u6_rem_96_22_Y_u6_div_90_17_n_804),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_256));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_804));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_805),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_200));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_787),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_805));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230077 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_797));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_141));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2859),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_796));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2859));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2858),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_795));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2858));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230098 (.A(u6_rem_96_22_Y_u6_div_90_17_n_794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_34));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_794));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230101 (.A(u6_rem_96_22_Y_u6_div_90_17_n_793),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2857));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230105 (.A(u6_rem_96_22_Y_u6_div_90_17_n_199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_793));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_199),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_799));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2850),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_199));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_792),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_791));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230114 (.A(n_3647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_788),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_792));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2856));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230118 (.A(u6_rem_96_22_Y_u6_div_90_17_n_789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_790));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2854),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_789));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2853),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2854));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230124 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2836),
    .B(n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2853));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230130 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2830),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2713),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_787));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230132 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .A2(n_3647),
    .B(n_13866),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2851));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230134 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2671),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_719),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_786));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230135 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2850));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230136 (.A(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2826),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2849));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2847),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2846));
 BUFx3_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2847));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2845),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_782));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2845));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_781));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230154 (.A(u6_rem_96_22_Y_u6_div_90_17_n_784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2844));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_784));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230161 (.A(u6_rem_96_22_Y_u6_div_90_17_n_118),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_785));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2829),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_118));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2842));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_33),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2843));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230185 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_33));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230186 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2841),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2840));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230190 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2841));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230191 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2838));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230192 (.A(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2839));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230194 (.A(u6_rem_96_22_Y_u6_div_90_17_n_198),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_778));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_198));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230204 (.A(u6_rem_96_22_Y_u6_div_90_17_n_117),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_780));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2660),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_117));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230208 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2836),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2837));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230209 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .A2(n_3647),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2831),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2836));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230211 (.A(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2834));
 NAND5xp2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230213 (.A(u6_rem_96_22_Y_u6_div_90_17_n_182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_721),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_705),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_2524),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2832));
 NOR5xp2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230214 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2758),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2755),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_703),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_688),
    .E(u6_rem_96_22_Y_u6_div_90_17_n_700),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2831));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230217 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2830),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_777));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230218 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2624),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_762),
    .B(n_13867),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2830));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230219 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_704),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_698),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2829));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230239 (.A(u6_rem_96_22_Y_u6_div_90_17_n_774),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_773));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230248 (.A(u6_rem_96_22_Y_u6_div_90_17_n_772),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_774));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_196),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_772));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230257 (.A(u6_rem_96_22_Y_u6_div_90_17_n_116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_196));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230268 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_116));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230279 (.A(u6_rem_96_22_Y_u6_div_90_17_n_775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_115));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230284 (.A(u6_rem_96_22_Y_u6_div_90_17_n_114),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_775));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230285 (.A(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_114));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230298 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_113));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_245),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_13));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_195),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_245));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_776),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_195));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_776));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230319 (.A(u6_rem_96_22_Y_u6_div_90_17_n_771),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_32));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230322 (.A(u6_rem_96_22_Y_u6_div_90_17_n_762),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_771));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_194),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_766));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230347 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_194));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_193),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_765));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230354 (.A(u6_rem_96_22_Y_u6_div_90_17_n_111),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_193));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_110),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_111));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_109),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_110));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230378 (.A(u6_rem_96_22_Y_u6_div_90_17_n_763),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_109));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230381 (.A(u6_rem_96_22_Y_u6_div_90_17_n_192),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_763));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230390 (.A(u6_rem_96_22_Y_u6_div_90_17_n_191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_192));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_191));
 XNOR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230399 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2821),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_770));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230400 (.A(u6_rem_96_22_Y_u6_div_90_17_n_702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2825),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2828));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230401 (.A(n_14269),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_704),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2827));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .B(n_14291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2826));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230405 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2724),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2823));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230406 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2723),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2822));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230407 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_688),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2552),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2821));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_704),
    .B(n_14269),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2820));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230409 (.A(u6_rem_96_22_Y_u6_div_90_17_n_182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_721),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2825));
 AOI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230410 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2772),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_762));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230423 (.A(u6_rem_96_22_Y_u6_div_90_17_n_754),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2818));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_754));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230431 (.A(u6_rem_96_22_Y_u6_div_90_17_n_190),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_753));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230433 (.A(u6_rem_96_22_Y_u6_div_90_17_n_755),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_190));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230438 (.A(u6_rem_96_22_Y_u6_div_90_17_n_756),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_755));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230445 (.A(u6_rem_96_22_Y_u6_div_90_17_n_189),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_756));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230448 (.A(u6_rem_96_22_Y_u6_div_90_17_n_752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_189));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_108),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_752));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230466 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2816),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_108));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_187),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2816));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_186),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_187));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_186));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230483 (.A(u6_rem_96_22_Y_u6_div_90_17_n_759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_107));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_759));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230489 (.A(n_14291),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_105));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2813));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_746));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230520 (.A(u6_rem_96_22_Y_u6_div_90_17_n_745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_30));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_104),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_745));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230524 (.A(u6_rem_96_22_Y_u6_div_90_17_n_185),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_104));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_185));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_184));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_183),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_40));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_183));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230572 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_743));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230584 (.A(u6_rem_96_22_Y_u6_div_90_17_n_749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_31));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230586 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2808));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2725),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2807));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2722),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2806));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230589 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2805));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230590 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2720),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2804));
 XOR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2753),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2672),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_749));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230593 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2749),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2803));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230594 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2577),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2802));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230595 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2801));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230596 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2573),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2800));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2578),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2752),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2799));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230603 (.A(u6_rem_96_22_Y_u6_div_90_17_n_182),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2796));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230608 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2795),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2794));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2563),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2750),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2793));
 O2A1O1Ixp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230610 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2572),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2652),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2716),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_739),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2792));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230611 (.A(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2798));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230613 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2539),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_182));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2795));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2791),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2790));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230616 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2789),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2788));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2782),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2783));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230622 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2781),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2780));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2778),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2779));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230625 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2775),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2776));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2771));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230629 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2769),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2768));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230630 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2766));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230631 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2765),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2764));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2762),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2763));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230633 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2760),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2761));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230637 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2758),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_739));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230640 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2757));
 NOR4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230641 (.A(u6_rem_96_22_Y_u6_div_90_17_n_693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_257),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_689),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2756));
 NAND4xp25_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230642 (.A(u6_rem_96_22_Y_u6_div_90_17_n_692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_697),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2534),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2755));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230643 (.A(u6_rem_96_22_Y_u6_div_90_17_n_707),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2754));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230644 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_700),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2545),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2753));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230645 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2791));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230646 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2693),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2789));
 MAJIxp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230647 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_740));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230648 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2692),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_716),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2787));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230649 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2786));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230650 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2785));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230651 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2784));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230652 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2782));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230653 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2781));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230654 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2778));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230655 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2708),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2777));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230656 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2775));
 OAI211xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230657 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2622),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_718),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_699),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2772));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230658 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2770));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230659 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2769));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230660 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2703),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2767));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230661 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2702),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2765));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230662 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2704),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2762));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230663 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2705),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2760));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230664 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2759));
 NAND4xp25_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230665 (.A(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_710),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_694),
    .D(u6_rem_96_22_Y_u6_div_90_17_n_695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2758));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230666 (.A(u6_rem_96_22_Y_u6_div_90_17_n_696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_738));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230667 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2751),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2752));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230668 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2748),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2749));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230669 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2746),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2747));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230670 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2745),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2744));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230673 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_730));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230682 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2742),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_733));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230683 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2742));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230689 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2741),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_732));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230690 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2741));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2740),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_734));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2740));
 INVx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230703 (.A(u6_rem_96_22_Y_u6_div_90_17_n_255),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_731));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_255));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_10));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230725 (.A(u6_rem_96_22_Y_u6_div_90_17_n_737),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_181));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_736),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_737));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230734 (.A(u6_rem_96_22_Y_u6_div_90_17_n_103),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_736));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230742 (.A(u6_rem_96_22_Y_u6_div_90_17_n_406),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_725));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_406));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230759 (.A(u6_rem_96_22_Y_u6_div_90_17_n_102),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_723));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_101),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_102));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230772 (.A(u6_rem_96_22_Y_u6_div_90_17_n_726),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_101));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_727),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_726));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230783 (.A(u6_rem_96_22_Y_u6_div_90_17_n_228),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_727));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230786 (.A(u6_rem_96_22_Y_u6_div_90_17_n_728),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_228));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230791 (.A(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_728));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_729),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2737));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230794 (.A(u6_rem_96_22_Y_u6_div_90_17_n_100),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_729));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230804 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2609),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2736));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2673),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_708),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2735));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230806 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2607),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2568),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2734));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230807 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2608),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2733));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230808 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2732));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230809 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2613),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2731));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230810 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2611),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2730));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2610),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2729));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2728));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230813 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2579),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2727));
 OAI211xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230814 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2649),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_719),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2541),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2726));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230815 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2454),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_716),
    .B2(n_3631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2751));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230816 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2508),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_716),
    .B2(n_3635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2725));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230817 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2459),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .B1(n_3627),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_715),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2724));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230818 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2458),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_716),
    .B2(n_3633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2723));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230819 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2509),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B2(n_3637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2722));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230820 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2457),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B2(n_3643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2721));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230821 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_716),
    .A2(n_3629),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2750));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230822 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2507),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B2(n_3641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2720));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230823 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2506),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B2(n_3639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2748));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230824 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B2(n_3839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2719));
 MAJIxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2574),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2746));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230826 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2745));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230827 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2657),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_103));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2540),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_100));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230829 (.A(u6_rem_96_22_Y_u6_div_90_17_n_717),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2718));
 A2O1A1Ixp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230830 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2511),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_708),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2717));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230831 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2572),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2716));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230832 (.A(u6_rem_96_22_Y_u6_div_90_17_n_722),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2715));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230834 (.A(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_710),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_722));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230836 (.A(u6_rem_96_22_Y_u6_div_90_17_n_721),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2714));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_721));
 NOR3xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230840 (.A(u6_rem_96_22_Y_u6_div_90_17_n_692),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2649),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_2543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2713));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230841 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2712));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2711));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230843 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2710));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2628),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2709));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230845 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2692),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2693));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230846 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2691));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230847 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2687));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230848 (.A(u6_rem_96_22_Y_u6_div_90_17_n_720),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2686));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230850 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2684),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2685));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230851 (.A(u6_rem_96_22_Y_u6_div_90_17_n_701),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2683));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230852 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2547),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2682));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2681));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230854 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2546),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2680));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230855 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2536),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2679));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2678));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230858 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2676));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230859 (.A1(n_3647),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2675));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230860 (.A(n_3641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2708));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230861 (.A(n_3641),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2707));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230862 (.A(n_3643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2706));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230863 (.A(n_3637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2705));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230864 (.A(n_3627),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2704));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230865 (.A(n_3631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2703));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230866 (.A(n_3639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2702));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230867 (.A(n_3637),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2701));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230868 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2567),
    .B(n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2700));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230869 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2564),
    .B(n_3629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2699));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230870 (.A(n_3633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2698));
 OAI21xp33_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230871 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2674));
 OAI22xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230872 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2511),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2673));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230873 (.A(n_3639),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2697));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230874 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2564),
    .B(n_3629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2696));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230875 (.A(n_3643),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2695));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230876 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .B2(u5_mul_69_18_n_89),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2672));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230877 (.A(n_3633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2694));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230878 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2544),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2671));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230879 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2692));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230880 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2690));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230881 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2551),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_688),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2670));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230882 (.A(u6_rem_96_22_Y_u6_div_90_17_n_711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2669));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230883 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2668));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230884 (.A(n_3631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2577),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2689));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230885 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2605),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2667));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230886 (.A(u6_rem_96_22_Y_u6_div_90_17_n_694),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2548),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2666));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230887 (.A(u6_rem_96_22_Y_u6_div_90_17_n_696),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2549),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2665));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230888 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .A2(n_14150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_690),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2664));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230889 (.A(u6_rem_96_22_Y_u6_div_90_17_n_691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2556),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2663));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2554),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2662));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230891 (.A(u6_rem_96_22_Y_u6_div_90_17_n_697),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2661));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230892 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2550),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_693),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2660));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230893 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2522),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_705),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2659));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230894 (.A(u6_rem_96_22_Y_u6_div_90_17_n_698),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2658));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230895 (.A(u6_rem_96_22_Y_u6_div_90_17_n_700),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2657));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230896 (.A(u6_rem_96_22_Y_u6_div_90_17_n_691),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2688));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230897 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2537),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_720));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_710),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_709),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2684));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230899 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2656));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230900 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2650),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2651));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230902 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2648));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230904 (.A(u6_rem_96_22_Y_u6_div_90_17_n_718),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2646));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230917 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_715));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230918 (.A(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2645));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230922 (.A(u6_rem_96_22_Y_u6_div_90_17_n_714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_716));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230924 (.A(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_714));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230936 (.A(u6_rem_96_22_Y_u6_div_90_17_n_713),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_717));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230939 (.A1(n_3634),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2565),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2655));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230940 (.A1(n_3630),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2643));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230941 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2457),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2642));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230942 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2459),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2641));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230943 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2508),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2640));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230944 (.A1(n_3642),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2570),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2639));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230945 (.A1(n_3629),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2638));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230946 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2511),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2637));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230947 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2597),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2636));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230949 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2509),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2634));
 AOI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230950 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2467),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_706),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2633));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230951 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .A2(n_3633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2632));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230952 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .A2(n_3631),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2590),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2631));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230953 (.A1(n_3636),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2575),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2630));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230954 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2629));
 NAND3xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230955 (.A(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .C(u5_mul_69_18_n_146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2628));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230956 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2627));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230957 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2626));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230958 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(n_14146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2625));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230959 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .B(n_14134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2624));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230960 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2623));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230961 (.A1(n_14128),
    .A2(n_14178),
    .B(n_14126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2622));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230962 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2460),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2654));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230963 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2621));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230964 (.A1(n_3628),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2653));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230965 (.A(u6_rem_96_22_Y_u6_div_90_17_n_702),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2527),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2620));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230966 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2483),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2619));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230967 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .A2(n_3639),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2652));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230968 (.A1(n_3626),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2650));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230969 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2618));
 AOI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230970 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2649));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230971 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_719));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230972 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2617));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230973 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .A2(n_3643),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2424),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2616));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230974 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .A2(n_14146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2615));
 AOI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230975 (.A1(n_14164),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2584),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2614));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230976 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2509),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .B2(n_3637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2613));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230977 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2507),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .B2(n_3641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2612));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230978 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_585),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .B2(n_3839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2611));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230979 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_44),
    .A2(n_3635),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2610));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230980 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2459),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .B2(n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2609));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230981 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .A2(n_3629),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2608));
 OAI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230982 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2458),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .B2(n_3633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2607));
 AOI22xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230983 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .A2(n_3631),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_496),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_2454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2606));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230984 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2463),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2647));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g230985 (.A1(n_14178),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(n_14124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_718));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g230986 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2528),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_713));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230988 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2605));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230990 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2600));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230994 (.A(u6_rem_96_22_Y_u6_div_90_17_n_710),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_711));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g230999 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2597));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231000 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2594),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2595));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231001 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2593),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2592));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231002 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2588));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231003 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2586),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2587));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231004 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2585),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2584));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2582));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231009 (.A(u6_rem_96_22_Y_u6_div_90_17_n_707),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_708));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231011 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2580),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2579));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231012 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2578),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2577));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231013 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2576),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2575));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231015 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2574),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_706));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231016 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2572));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231017 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2570));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231018 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2568));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231019 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2566));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231020 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2564),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2563));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231021 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2562));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231022 (.A(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2561));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231025 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .B(n_3646),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2559));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231026 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2604));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231027 (.A(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2603));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231028 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_230),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2558));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231029 (.A(n_14164),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2602));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231030 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2557));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_712));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231032 (.A(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .B(n_3643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2601));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231035 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_709));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .B(n_3839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2596));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231038 (.A(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2506),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2594));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231039 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2593));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231040 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2591));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231041 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2590));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .B(n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2589));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231043 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2586));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231044 (.A(u6_rem_96_22_Y_u6_div_90_17_n_584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2585));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231045 (.A(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2510),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2583));
 NAND2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231046 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(n_14270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_707));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231047 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2464),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2580));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231048 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2578));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231049 (.A(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2521),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2576));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231050 (.A(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .B(n_3838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2574));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231051 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2460),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2573));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2571));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231053 (.A(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2463),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2569));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2567));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231055 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .B(n_3634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2565));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231056 (.A(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2564));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231059 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2553),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2554));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231060 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2552));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231061 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2547),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2548));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231063 (.A(u6_rem_96_22_Y_u6_div_90_17_n_703),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_704));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_701),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_702));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231071 (.A(u6_rem_96_22_Y_u6_div_90_17_n_699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2545));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231074 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2544));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2541),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2542));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231079 (.A(u6_rem_96_22_Y_u6_div_90_17_n_257),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_697));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231080 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2539),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2538));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231084 (.A(u6_rem_96_22_Y_u6_div_90_17_n_695),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_696));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231085 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2537),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2536));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231086 (.A(u6_rem_96_22_Y_u6_div_90_17_n_694),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2535));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231093 (.A(u6_rem_96_22_Y_u6_div_90_17_n_691),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2534));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231102 (.A(u6_rem_96_22_Y_u6_div_90_17_n_689),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_690));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231108 (.A(u6_rem_96_22_Y_u6_div_90_17_n_687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_688));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231109 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2533),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2532));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231113 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2530),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_685));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2530));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231125 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_684));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231129 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2529));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2531),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_686));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231135 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2528));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231136 (.A(n_14130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2527));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231137 (.A(n_14128),
    .B(n_14126),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2526));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231138 (.A(n_14150),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2525));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231139 (.A(n_14134),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_705));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231140 (.A(n_14146),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2556));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231141 (.A(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2555));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231142 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_648),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2553));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2524));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231144 (.A(n_14130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_492),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2551));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231145 (.A(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2523));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2550));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231147 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2549));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2522));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231149 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2547));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231150 (.A(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_703));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231151 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2442),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2546));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231152 (.A(n_14132),
    .B(n_14130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_701));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231153 (.A(u5_mul_69_18_n_89),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_700));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231154 (.A(n_14126),
    .B(n_14178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_699));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231155 (.A(u6_rem_96_22_Y_u6_div_90_17_n_523),
    .B(n_14134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_698));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231156 (.A(u6_rem_96_22_Y_u6_div_90_17_n_20),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2543));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231157 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2541));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231158 (.A(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_588),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2540));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231160 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2539));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231161 (.A(u5_mul_69_18_n_130),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_695));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2537));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231163 (.A(u6_rem_96_22_Y_u6_div_90_17_n_668),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_694));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231164 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2477),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_693));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231165 (.A(n_14136),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_692));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231166 (.A(u6_rem_96_22_Y_u6_div_90_17_n_655),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_691));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231167 (.A(u6_rem_96_22_Y_u6_div_90_17_n_661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_689));
 NOR2xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231168 (.A(n_14130),
    .B(n_14128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_687));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231169 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2533));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231170 (.A(u6_rem_96_22_Y_u6_div_90_17_n_378),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2531));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231171 (.A(n_3636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2521));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231172 (.A(n_3642),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2520));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231174 (.A(n_3626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2518));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231175 (.A(n_3645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2517));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231176 (.A(u6_rem_96_22_Y_u6_div_90_17_n_683),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2511));
 BUFx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231183 (.A(n_3645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_683));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231184 (.A(n_3629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2510));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231185 (.A(n_3637),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2509));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231186 (.A(n_3635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2508));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231187 (.A(n_3641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2507));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231188 (.A(n_3639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2506));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231202 (.A(u6_rem_96_22_Y_u6_div_90_17_n_675),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_676));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231209 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_675));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231226 (.A(u6_rem_96_22_Y_u6_div_90_17_n_678),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_677));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231228 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_678));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231232 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_679));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231234 (.A(u6_rem_96_22_Y_u6_div_90_17_n_180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_7));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_680),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_180));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231252 (.A(u6_rem_96_22_Y_u6_div_90_17_n_179),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_680));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231259 (.A(u6_rem_96_22_Y_u6_div_90_17_n_681),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_179));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231262 (.A(u5_mul_69_18_n_143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_681));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231293 (.A(u6_rem_96_22_Y_u6_div_90_17_n_669),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_379));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231301 (.A(u6_rem_96_22_Y_u6_div_90_17_n_670),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_669));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231307 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_670));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_671));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231318 (.A(u6_rem_96_22_Y_u6_div_90_17_n_673),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_178));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231325 (.A(u6_rem_96_22_Y_u6_div_90_17_n_99),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_673));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_99));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_674),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_668));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231371 (.A(u6_rem_96_22_Y_u6_div_90_17_n_663),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_664));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231372 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_663));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231393 (.A(u6_rem_96_22_Y_u6_div_90_17_n_404),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_665));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231395 (.A(u6_rem_96_22_Y_u6_div_90_17_n_662),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_404));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231403 (.A(u6_rem_96_22_Y_u6_div_90_17_n_98),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_662));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231411 (.A(u6_rem_96_22_Y_u6_div_90_17_n_29),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_98));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231430 (.A(u6_rem_96_22_Y_u6_div_90_17_n_393),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_29));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231433 (.A(n_14152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_393));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231455 (.A(u6_rem_96_22_Y_u6_div_90_17_n_96),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_656));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_657),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_96));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_658),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_657));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_658));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231477 (.A(u6_rem_96_22_Y_u6_div_90_17_n_244),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_229));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_659),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_244));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_95),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_659));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_95));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_227),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_660));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231516 (.A(n_14150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_227));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231529 (.A(n_14150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_661));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2500));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_651),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_650));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_651));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231577 (.A(u6_rem_96_22_Y_u6_div_90_17_n_254),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_652));
 BUFx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_254));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_653),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_654));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231588 (.A(u6_rem_96_22_Y_u6_div_90_17_n_392),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_653));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231598 (.A(u6_rem_96_22_Y_u6_div_90_17_n_94),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_392));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231609 (.A(u6_rem_96_22_Y_u6_div_90_17_n_93),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_94));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231614 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_93));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231617 (.A(n_14146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2501));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231630 (.A(n_14146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_655));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231649 (.A(u6_rem_96_22_Y_u6_div_90_17_n_391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_644));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231657 (.A(u6_rem_96_22_Y_u6_div_90_17_n_645),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_391));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_645));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_647),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_92));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_647));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231696 (.A(u6_rem_96_22_Y_u6_div_90_17_n_172),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_226));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231702 (.A(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_172));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231726 (.A(u6_rem_96_22_Y_u6_div_90_17_n_91),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_648));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231729 (.A(u6_rem_96_22_Y_u6_div_90_17_n_643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_91));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231754 (.A(u6_rem_96_22_Y_u6_div_90_17_n_634),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_243));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231767 (.A(u6_rem_96_22_Y_u6_div_90_17_n_635),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_634));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231768 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_635));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231775 (.A(u6_rem_96_22_Y_u6_div_90_17_n_242),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_90));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231787 (.A(u6_rem_96_22_Y_u6_div_90_17_n_636),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_242));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231788 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_636));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231801 (.A(u6_rem_96_22_Y_u6_div_90_17_n_27),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_390));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g231812 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_27));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231820 (.A(u6_rem_96_22_Y_u6_div_90_17_n_638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_637));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231825 (.A(u6_rem_96_22_Y_u6_div_90_17_n_639),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_638));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231828 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_639));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231839 (.A(u6_rem_96_22_Y_u6_div_90_17_n_640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_28));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231850 (.A(n_14142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_640));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_631));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231890 (.A(u6_rem_96_22_Y_u6_div_90_17_n_623),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_389));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231898 (.A(u6_rem_96_22_Y_u6_div_90_17_n_624),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_623));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231906 (.A(u6_rem_96_22_Y_u6_div_90_17_n_625),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_624));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231928 (.A(u6_rem_96_22_Y_u6_div_90_17_n_626),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_625));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231937 (.A(u6_rem_96_22_Y_u6_div_90_17_n_627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_626));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231946 (.A(u6_rem_96_22_Y_u6_div_90_17_n_88),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_627));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231949 (.A(u6_rem_96_22_Y_u6_div_90_17_n_87),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_88));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231951 (.A(u6_rem_96_22_Y_u6_div_90_17_n_628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_87));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_26));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231961 (.A(u6_rem_96_22_Y_u6_div_90_17_n_629),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_628));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231963 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2494),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_629));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_171),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2494));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231969 (.A(u6_rem_96_22_Y_u6_div_90_17_n_630),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_171));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231971 (.A(u6_rem_96_22_Y_u6_div_90_17_n_622),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_630));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231980 (.A(u6_rem_96_22_Y_u6_div_90_17_n_170),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_622));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231984 (.A(u6_rem_96_22_Y_u6_div_90_17_n_631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_170));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g231989 (.A(u6_rem_96_22_Y_u6_div_90_17_n_86),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_632));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231991 (.A(u6_rem_96_22_Y_u6_div_90_17_n_86),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2488));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231997 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_86));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g231998 (.A(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2487));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232005 (.A(u6_rem_96_22_Y_u6_div_90_17_n_169),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2483));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232010 (.A(n_14178),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_169));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232031 (.A(u6_rem_96_22_Y_u6_div_90_17_n_615),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2480));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232042 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2480),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_614));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_615));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232067 (.A(u6_rem_96_22_Y_u6_div_90_17_n_85),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_403));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_377),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_85));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232087 (.A(u6_rem_96_22_Y_u6_div_90_17_n_84),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_377));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232096 (.A(u6_rem_96_22_Y_u6_div_90_17_n_232),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_84));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232100 (.A(u6_rem_96_22_Y_u6_div_90_17_n_82),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_232));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232112 (.A(u6_rem_96_22_Y_u6_div_90_17_n_80),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_82));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232123 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2481),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_80));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232124 (.A(u6_rem_96_22_Y_u6_div_90_17_n_619),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2481));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232127 (.A(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_619));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232130 (.A(u6_rem_96_22_Y_u6_div_90_17_n_618),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2478));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232131 (.A(u6_rem_96_22_Y_u6_div_90_17_n_168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_618));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232140 (.A(u6_rem_96_22_Y_u6_div_90_17_n_621),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_168));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232143 (.A(u6_rem_96_22_Y_u6_div_90_17_n_620),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_621));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232160 (.A(n_14134),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_620));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232161 (.A(n_14136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2477));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232177 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2474));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_607),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_79));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232197 (.A(u6_rem_96_22_Y_u6_div_90_17_n_77),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_607));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232201 (.A(u6_rem_96_22_Y_u6_div_90_17_n_78),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_77));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232206 (.A(u6_rem_96_22_Y_u6_div_90_17_n_608),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_78));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232212 (.A(u6_rem_96_22_Y_u6_div_90_17_n_166),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_608));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232219 (.A(u6_rem_96_22_Y_u6_div_90_17_n_76),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_166));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_388),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_76));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_609),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_388));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232243 (.A(u6_rem_96_22_Y_u6_div_90_17_n_610),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_609));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232244 (.A(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_610));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232246 (.A(u6_rem_96_22_Y_u6_div_90_17_n_165),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2473));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232251 (.A(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_165));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232263 (.A(u6_rem_96_22_Y_u6_div_90_17_n_164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_167));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232265 (.A(u6_rem_96_22_Y_u6_div_90_17_n_75),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_164));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232278 (.A(u6_rem_96_22_Y_u6_div_90_17_n_606),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_75));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232280 (.A(u6_rem_96_22_Y_u6_div_90_17_n_613),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_606));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232293 (.A(n_14136),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_613));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232320 (.A(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_25));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232326 (.A(u6_rem_96_22_Y_u6_div_90_17_n_598),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_597));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232327 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_598));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232349 (.A(u6_rem_96_22_Y_u6_div_90_17_n_402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_599));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232351 (.A(u6_rem_96_22_Y_u6_div_90_17_n_73),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_402));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232357 (.A(u6_rem_96_22_Y_u6_div_90_17_n_74),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_73));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232367 (.A(u6_rem_96_22_Y_u6_div_90_17_n_600),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_74));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232368 (.A(u6_rem_96_22_Y_u6_div_90_17_n_72),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_600));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232387 (.A(u6_rem_96_22_Y_u6_div_90_17_n_601),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_72));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232388 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_601));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232402 (.A(u6_rem_96_22_Y_u6_div_90_17_n_162),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_596));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232408 (.A(u6_rem_96_22_Y_u6_div_90_17_n_602),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_162));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232410 (.A(u6_rem_96_22_Y_u6_div_90_17_n_604),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_602));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232415 (.A(u6_rem_96_22_Y_u6_div_90_17_n_603),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_604));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232422 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_603));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232424 (.A(n_14130),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_6));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232441 (.A(u6_rem_96_22_Y_u6_div_90_17_n_387),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2469));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_231));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2469),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_5));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_591),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_387));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_386),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_591));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_592),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_386));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_589),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_592));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232508 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_589));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_70),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_588));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232525 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2467),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2468));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232526 (.A(n_3838),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2467));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_587),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2466));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232529 (.A(n_14270),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_587));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232531 (.A(n_3640),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2464));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232532 (.A(n_3632),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2463));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232534 (.A(n_3628),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2461));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232535 (.A(n_3638),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2460));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232536 (.A(n_3627),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2459));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232537 (.A(n_3633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2458));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232538 (.A(n_3643),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2457));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232545 (.A(n_3839),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_585));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232548 (.A(n_3631),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2454));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_579));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232574 (.A(u6_rem_96_22_Y_u6_div_90_17_n_401),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_580));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_581),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_401));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_583),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_581));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_582),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_583));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232609 (.A(n_14164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_582));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232617 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2449),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2450));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232621 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2449));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232623 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2448),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_578));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232626 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2448));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232628 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2447),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_577));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2447));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232638 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_576));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232640 (.A(fractb_mul[23]),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2445));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232674 (.A(u6_rem_96_22_Y_u6_div_90_17_n_571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_570));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232675 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_571));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232685 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2443));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232686 (.A(u6_rem_96_22_Y_u6_div_90_17_n_241),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_12));
 HB1xp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232687 (.A(u6_rem_96_22_Y_u6_div_90_17_n_572),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_241));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232692 (.A(u6_rem_96_22_Y_u6_div_90_17_n_253),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_572));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232697 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_253));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232714 (.A(u6_rem_96_22_Y_u6_div_90_17_n_573),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_230));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232717 (.A(n_14160),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_573));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232737 (.A(u6_rem_96_22_Y_u6_div_90_17_n_567),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_160));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232741 (.A(u6_rem_96_22_Y_u6_div_90_17_n_566),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_567));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232749 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_566));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232760 (.A(u6_rem_96_22_Y_u6_div_90_17_n_400),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_565));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232763 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_400));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_569),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_564));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_252),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_569));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232784 (.A(u6_rem_96_22_Y_u6_div_90_17_n_563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2442));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232792 (.A(u6_rem_96_22_Y_u6_div_90_17_n_563),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_252));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232797 (.A(n_14156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_563));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232819 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_556));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232830 (.A(u6_rem_96_22_Y_u6_div_90_17_n_557),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2440));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232838 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_557));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232842 (.A(u6_rem_96_22_Y_u6_div_90_17_n_159),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2439));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232844 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_159));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232849 (.A(u6_rem_96_22_Y_u6_div_90_17_n_158),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_559));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232853 (.A(u6_rem_96_22_Y_u6_div_90_17_n_560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_158));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232856 (.A(u6_rem_96_22_Y_u6_div_90_17_n_560),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2438));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232857 (.A(u6_rem_96_22_Y_u6_div_90_17_n_157),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_560));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232859 (.A(u6_rem_96_22_Y_u6_div_90_17_n_251),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_157));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232863 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_251));
 INVxp67_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232870 (.A(u6_rem_96_22_Y_u6_div_90_17_n_561),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_24));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232884 (.A(n_14154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_561));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232912 (.A(u6_rem_96_22_Y_u6_div_90_17_n_550),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_225));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232929 (.A(u6_rem_96_22_Y_u6_div_90_17_n_250),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_550));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232932 (.A(u6_rem_96_22_Y_u6_div_90_17_n_551),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_250));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g232940 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_551));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232960 (.A(u6_rem_96_22_Y_u6_div_90_17_n_69),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_68));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g232962 (.A(u6_rem_96_22_Y_u6_div_90_17_n_23),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_69));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232978 (.A(u6_rem_96_22_Y_u6_div_90_17_n_555),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_23));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g232980 (.A(n_14148),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_555));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233014 (.A(u6_rem_96_22_Y_u6_div_90_17_n_67),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_21));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_540),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_67));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233037 (.A(u6_rem_96_22_Y_u6_div_90_17_n_543),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_540));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233052 (.A(u6_rem_96_22_Y_u6_div_90_17_n_542),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_543));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233054 (.A(u6_rem_96_22_Y_u6_div_90_17_n_544),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_542));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_65),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_544));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233075 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_65));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233082 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_4));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233091 (.A(u6_rem_96_22_Y_u6_div_90_17_n_22),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_546));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233092 (.A(u6_rem_96_22_Y_u6_div_90_17_n_156),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_22));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233115 (.A(u6_rem_96_22_Y_u6_div_90_17_n_538),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_156));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233117 (.A(n_14140),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_538));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233146 (.A(u6_rem_96_22_Y_u6_div_90_17_n_62),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_526));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233148 (.A(u6_rem_96_22_Y_u6_div_90_17_n_240),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_62));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233162 (.A(u6_rem_96_22_Y_u6_div_90_17_n_61),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_240));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233165 (.A(u6_rem_96_22_Y_u6_div_90_17_n_528),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_61));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233168 (.A(u6_rem_96_22_Y_u6_div_90_17_n_529),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_528));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233169 (.A(u6_rem_96_22_Y_u6_div_90_17_n_60),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_529));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233178 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_60));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233189 (.A(u6_rem_96_22_Y_u6_div_90_17_n_532),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_531));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233193 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_532));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233198 (.A(u6_rem_96_22_Y_u6_div_90_17_n_59),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_533));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233199 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_59));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233221 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_63));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233224 (.A(u6_rem_96_22_Y_u6_div_90_17_n_154),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_20));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233235 (.A(u6_rem_96_22_Y_u6_div_90_17_n_155),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_154));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233249 (.A(u6_rem_96_22_Y_u6_div_90_17_n_56),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_519));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233275 (.A(u6_rem_96_22_Y_u6_div_90_17_n_514),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_513));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233277 (.A(u6_rem_96_22_Y_u6_div_90_17_n_515),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_514));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233286 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_515));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233295 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_385));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233299 (.A(u6_rem_96_22_Y_u6_div_90_17_n_516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_18));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233303 (.A(u6_rem_96_22_Y_u6_div_90_17_n_517),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_516));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233316 (.A(u6_rem_96_22_Y_u6_div_90_17_n_19),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_517));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233323 (.A(u6_rem_96_22_Y_u6_div_90_17_n_518),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_19));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233333 (.A(u6_rem_96_22_Y_u6_div_90_17_n_152),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_518));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233340 (.A(u6_rem_96_22_Y_u6_div_90_17_n_57),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_152));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233342 (.A(u6_rem_96_22_Y_u6_div_90_17_n_58),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_57));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_58));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233355 (.A(u6_rem_96_22_Y_u6_div_90_17_n_151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_56));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233364 (.A(u6_rem_96_22_Y_u6_div_90_17_n_520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_151));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233365 (.A(u6_rem_96_22_Y_u6_div_90_17_n_55),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_520));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233379 (.A(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_55));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233391 (.A(u6_rem_96_22_Y_u6_div_90_17_n_524),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_523));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233392 (.A(n_14132),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_524));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233427 (.A(u6_rem_96_22_Y_u6_div_90_17_n_501),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_502));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233436 (.A(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_501));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233440 (.A(u6_rem_96_22_Y_u6_div_90_17_n_150),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_500));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_150));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233459 (.A(u6_rem_96_22_Y_u6_div_90_17_n_503),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_499));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_503));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_3));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_54),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_504));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_249),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_54));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233493 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_249));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_53),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_507));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_17),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_53));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_508),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_17));
 INVx1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233531 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_508));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_41));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_0),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_51));
 INVx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233554 (.A(u5_mul_69_18_n_89),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_0));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_144));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233576 (.A(u6_rem_96_22_Y_u6_div_90_17_n_493),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_494));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_49),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_493));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233581 (.A(u6_rem_96_22_Y_u6_div_90_17_n_48),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_49));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233585 (.A(u6_rem_96_22_Y_u6_div_90_17_n_47),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_48));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233592 (.A(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_47));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233597 (.A(u6_rem_96_22_Y_u6_div_90_17_n_147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2422));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233599 (.A(u6_rem_96_22_Y_u6_div_90_17_n_146),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_147));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233606 (.A(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_146));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233615 (.A(u6_rem_96_22_Y_u6_div_90_17_n_145),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_378));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233618 (.A(u6_rem_96_22_Y_u6_div_90_17_n_16),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_145));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233632 (.A(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_16));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233636 (.A(u6_rem_96_22_Y_u6_div_90_17_n_495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_496));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233639 (.A(u6_rem_96_22_Y_u6_div_90_17_n_46),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_495));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233652 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2423),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_46));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233653 (.A(u6_rem_96_22_Y_u6_div_90_17_n_44),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2423));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233655 (.A(u6_rem_96_22_Y_u6_div_90_17_n_45),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_44));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233663 (.A(u6_rem_96_22_Y_u6_div_90_17_n_497),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_45));
 HB1xp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233664 (.A(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_497));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233672 (.A(u6_rem_96_22_Y_u6_div_90_17_n_144),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2424));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233684 (.A(u6_rem_96_22_Y_u6_div_90_17_n_50),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2));
 BUFx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233687 (.A(n_14124),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_50));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233711 (.A(u6_rem_96_22_Y_u6_div_90_17_n_486),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2419));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233715 (.A(u6_rem_96_22_Y_u6_div_90_17_n_487),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_486));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233716 (.A(u6_rem_96_22_Y_u6_div_90_17_n_399),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_487));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233731 (.A(u6_rem_96_22_Y_u6_div_90_17_n_485),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_399));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233743 (.A(u6_rem_96_22_Y_u6_div_90_17_n_484),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_485));
 BUFx2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233751 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_484));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233755 (.A(u6_rem_96_22_Y_u6_div_90_17_n_398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_2418));
 HB1xp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233765 (.A(u6_rem_96_22_Y_u6_div_90_17_n_143),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_398));
 INVxp67_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_143));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233795 (.A(u6_rem_96_22_Y_u6_div_90_17_n_142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_224));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233797 (.A(u6_rem_96_22_Y_u6_div_90_17_n_490),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_142));
 INVxp67_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233805 (.A(u6_rem_96_22_Y_u6_div_90_17_n_43),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_490));
 INVxp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233811 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_43));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233818 (.A(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1));
 INVx1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g233826 (.A(u6_rem_96_22_Y_u6_div_90_17_n_42),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_492));
 INVx1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g233827 (.A(n_14128),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_42));
 INVx2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g233964 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13699),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_457));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234033 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_1465));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234069 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11941),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11974),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_445));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234121 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5670),
    .B(u6_n_105),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_439));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234207 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8495),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_430));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234348 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11396),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_465));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234356 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7920),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7909),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_422));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234389 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7293),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7340),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_443));
 INVx3_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234416 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_433));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234424 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6155),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6181),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_219));
 AND2x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234432 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5177),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5147),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_411));
 NOR2x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234440 (.A(fractb_mul[23]),
    .B(n_14164),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_710));
 OAI21xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234441 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_2540),
    .A2(n_3646),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2837),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_788));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234442 (.A(u6_rem_96_22_Y_u6_div_90_17_n_743),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_975),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_409));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234450 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13661),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13461),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_375));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234451 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13660),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13457),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_374));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234452 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13379),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2402),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_373));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234453 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13426),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2398),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_372));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234454 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13436),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13337),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_371));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234456 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12822),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_13090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_369));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234457 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13080),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12843),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_368));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234458 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13060),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12808),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_367));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234459 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_12876),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2322),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12913),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_366));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234460 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12825),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2321),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_365));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234461 (.A(u6_rem_96_22_Y_u6_div_90_17_n_13002),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12803),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_364));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234462 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12788),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_363));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234463 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12682),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12824),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_362));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234464 (.A(u6_rem_96_22_Y_u6_div_90_17_n_579),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12652),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_361));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234465 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12598),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12353),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_360));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234467 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12469),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12266),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_358));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234468 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_12218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_357));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234469 (.A(u6_rem_96_22_Y_u6_div_90_17_n_12019),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11738),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_356));
 XNOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234470 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11939),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11687),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_355));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234471 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11938),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11723),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_354));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234472 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11926),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11725),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_353));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234473 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11777),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11896),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_352));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234474 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11720),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2169),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11797),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_351));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234475 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11671),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2168),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_350));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234476 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11709),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11546),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_349));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234477 (.A(u6_rem_96_22_Y_u6_div_90_17_n_141),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11520),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_348));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234478 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11331),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11090),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_347));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234480 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11302),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_346));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234481 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11116),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_345));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234482 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11250),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11046),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_344));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234483 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11249),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11049),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_343));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234484 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11076),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2101),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11151),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_342));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234486 (.A(u6_rem_96_22_Y_u6_div_90_17_n_403),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10903),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_340));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234487 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10771),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10571),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_339));
 AND2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234488 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10595),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10770),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_338));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234489 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10597),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10764),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_337));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234490 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10699),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10526),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_336));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234491 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10695),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10522),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_335));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234492 (.A(u6_rem_96_22_Y_u6_div_90_17_n_333),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10519),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_334));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234493 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_10599),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_2042),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10633),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_333));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234494 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_10391),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_332));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234495 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10152),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9899),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_331));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234496 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10149),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9932),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_330));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234497 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10148),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9892),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_329));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234498 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10143),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9898),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_328));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234499 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10121),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9885),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_327));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234500 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10097),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9881),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_326));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234501 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10096),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9887),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_325));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234502 (.A(u6_rem_96_22_Y_u6_div_90_17_n_10035),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1986),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_324));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234503 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9811),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9794),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_323));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234504 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9585),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9339),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_322));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234505 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9584),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9338),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_321));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234506 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9553),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_9350),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_320));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234507 (.A(u6_rem_96_22_Y_u6_div_90_17_n_9031),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8767),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_319));
 AO21x1_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234508 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8808),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8958),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8844),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_318));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234509 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1837),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8810),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_317));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234510 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8461),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8200),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_316));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234511 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8446),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8180),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_315));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234512 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8427),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8197),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_314));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234513 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8414),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8221),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_313));
 AO21x1_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234514 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_8330),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_8381),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8361),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_312));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234515 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8382),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8177),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_311));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234516 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8371),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8176),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_310));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234517 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8369),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8191),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_309));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234518 (.A(u6_rem_96_22_Y_u6_div_90_17_n_8040),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_8210),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_308));
 XOR2xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234519 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7902),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7596),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_307));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234521 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7672),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7894),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_305));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234522 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7865),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7612),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_304));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234523 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7864),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7644),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_303));
 AO21x1_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234525 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_7679),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_1721),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7711),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_301));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234526 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7683),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1714),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_300));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234527 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7633),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7475),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_299));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234528 (.A(u6_rem_96_22_Y_u6_div_90_17_n_839),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7454),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_298));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234529 (.A(u6_rem_96_22_Y_u6_div_90_17_n_185),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7430),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_297));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234530 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7307),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7099),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_296));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234532 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7304),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7055),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_294));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234533 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7081),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7301),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_293));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234534 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7219),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7106),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_292));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234535 (.A(u6_rem_96_22_Y_u6_div_90_17_n_7120),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_7123),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_291));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234536 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6711),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6516),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_290));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234537 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1560),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_6415),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_289));
 NOR2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234539 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1475),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1482),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_287));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234540 (.A(u6_rem_96_22_Y_u6_div_90_17_n_184),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1471),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_286));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234541 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6128),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5963),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_285));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234542 (.A(u6_rem_96_22_Y_u6_div_90_17_n_6092),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5923),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_284));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234543 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5953),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_1446),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_283));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234544 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5642),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5413),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_282));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234546 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5576),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5394),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_281));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234548 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4931),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_5107),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_279));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234549 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5071),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4886),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_278));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234550 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5068),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4951),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_277));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234552 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5059),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4943),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_275));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234553 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4832),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4814),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_274));
 AND2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234554 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4497),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4641),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_273));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234555 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4638),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4509),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_272));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234557 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4616),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4511),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_270));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234558 (.A(u6_rem_96_22_Y_u6_div_90_17_n_1145),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4488),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_269));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234560 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4111),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4218),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_268));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234561 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4216),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4116),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_267));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234562 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4182),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4096),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_266));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234563 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3542),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3470),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_265));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234564 (.A(u6_rem_96_22_Y_u6_div_90_17_n_970),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3466),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_264));
 XNOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234565 (.A(u6_rem_96_22_Y_u6_div_90_17_n_921),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_3247),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_263));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234567 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5395),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2786),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_262));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234568 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3093),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2785),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_261));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234569 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3449),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2784),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_260));
 XNOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234570 (.A(u6_rem_96_22_Y_u6_div_90_17_n_3251),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2777),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_259));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234571 (.A(u6_rem_96_22_Y_u6_div_90_17_n_5390),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2759),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_258));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234573 (.A(n_14140),
    .B(n_14142),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_257));
 XOR2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234578 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11314),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11060),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_223));
 OR2x2_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234579 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4879),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4848),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_222));
 XOR2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234580 (.A(u6_rem_96_22_Y_u6_div_90_17_n_4612),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_4489),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_221));
 XOR2x2_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234583 (.A(u6_rem_96_22_Y_u6_div_90_17_n_2959),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_2445),
    .Y(u6_rem_96_22_Y_u6_div_90_17_n_220));
 HAxp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234587 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11879),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11680),
    .CON(UNCONNECTED),
    .SN(u6_rem_96_22_Y_u6_div_90_17_n_2185));
 INVx2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234761 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11396),
    .Y(n_854));
 NAND2xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234762 (.A(n_14014),
    .B(u6_rem_96_22_Y_u6_div_90_17_n_11368),
    .Y(n_14015));
 AND2x4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234763 (.A(n_14012),
    .B(n_854),
    .Y(n_14014));
 OAI21xp33_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234765 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11347),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11348),
    .B(n_14014),
    .Y(n_14017));
 OAI21xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234766 (.A1(n_14468),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11318),
    .B(n_14014),
    .Y(n_14018));
 INVx4_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234767 (.A(n_14014),
    .Y(n_14019));
 OAI21xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234768 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11285),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11284),
    .B(n_14014),
    .Y(n_14020));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234769 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11274),
    .B(n_14014),
    .Y(n_14021));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234770 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11343),
    .B(n_14014),
    .Y(n_14022));
 NAND2xp5_ASAP7_75t_R u6_rem_96_22_Y_u6_div_90_17_g234771 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11353),
    .B(n_14014),
    .Y(n_14023));
 AOI22xp5_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234772 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11399),
    .A2(n_14024),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11412),
    .Y(n_14025));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234773 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11402),
    .B(n_14024),
    .Y(n_14026));
 AO221x2_ASAP7_75t_SL u6_rem_96_22_Y_u6_div_90_17_g234775 (.A1(n_14024),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11389),
    .B1(u6_rem_96_22_Y_u6_div_90_17_n_423),
    .B2(u6_rem_96_22_Y_u6_div_90_17_n_11390),
    .C(u6_rem_96_22_Y_u6_div_90_17_n_11467),
    .Y(n_14028));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234776 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11201),
    .B(n_14024),
    .Y(n_14029));
 NAND2xp5_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234777 (.A(u6_rem_96_22_Y_u6_div_90_17_n_11370),
    .B(n_14024),
    .Y(n_14030));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234778 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_345),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11316),
    .B(n_14024),
    .Y(n_14031));
 OAI21xp33_ASAP7_75t_L u6_rem_96_22_Y_u6_div_90_17_g234779 (.A1(u6_rem_96_22_Y_u6_div_90_17_n_11315),
    .A2(u6_rem_96_22_Y_u6_div_90_17_n_11317),
    .B(n_14024),
    .Y(n_14032));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[0]  (.CLK(clk),
    .D(n_14056),
    .QN(remainder[0]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[10]  (.CLK(clk),
    .D(n_14066),
    .QN(remainder[10]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[11]  (.CLK(clk),
    .D(n_14067),
    .QN(remainder[11]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[12]  (.CLK(clk),
    .D(n_14068),
    .QN(remainder[12]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[13]  (.CLK(clk),
    .D(n_14069),
    .QN(remainder[13]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[14]  (.CLK(clk),
    .D(n_14070),
    .QN(remainder[14]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[15]  (.CLK(clk),
    .D(n_14071),
    .QN(remainder[15]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[16]  (.CLK(clk),
    .D(n_14072),
    .QN(remainder[16]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[17]  (.CLK(clk),
    .D(n_14073),
    .QN(remainder[17]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[18]  (.CLK(clk),
    .D(n_14074),
    .QN(remainder[18]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[19]  (.CLK(clk),
    .D(n_14075),
    .QN(remainder[19]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[1]  (.CLK(clk),
    .D(n_14057),
    .QN(remainder[1]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[20]  (.CLK(clk),
    .D(n_14076),
    .QN(remainder[20]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[21]  (.CLK(clk),
    .D(n_14077),
    .QN(remainder[21]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[22]  (.CLK(clk),
    .D(n_14078),
    .QN(remainder[22]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[23]  (.CLK(clk),
    .D(n_14079),
    .QN(remainder[23]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[2]  (.CLK(clk),
    .D(n_14058),
    .QN(remainder[2]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[3]  (.CLK(clk),
    .D(n_14059),
    .QN(remainder[3]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[4]  (.CLK(clk),
    .D(n_14060),
    .QN(remainder[4]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[5]  (.CLK(clk),
    .D(n_14061),
    .QN(remainder[5]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[6]  (.CLK(clk),
    .D(n_14062),
    .QN(remainder[6]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[7]  (.CLK(clk),
    .D(n_14063),
    .QN(remainder[7]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[8]  (.CLK(clk),
    .D(n_14064),
    .QN(remainder[8]));
 DFFHQNx1_ASAP7_75t_R \u6_rem_reg[9]  (.CLK(clk),
    .D(n_14065),
    .QN(remainder[9]));
 DFFHQNx1_ASAP7_75t_L \u6_remainder_reg[0]  (.CLK(clk),
    .D(n_14054),
    .QN(n_14055));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[10]  (.CLK(clk),
    .D(u6_n_136),
    .Q(u6_remainder[10]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[11]  (.CLK(clk),
    .D(u6_n_137),
    .Q(u6_remainder[11]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[12]  (.CLK(clk),
    .D(u6_n_138),
    .Q(u6_remainder[12]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[13]  (.CLK(clk),
    .D(u6_n_139),
    .Q(u6_remainder[13]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[14]  (.CLK(clk),
    .D(u6_n_140),
    .Q(u6_remainder[14]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[15]  (.CLK(clk),
    .D(u6_n_141),
    .Q(u6_remainder[15]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[16]  (.CLK(clk),
    .D(u6_n_142),
    .Q(u6_remainder[16]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[17]  (.CLK(clk),
    .D(u6_n_143),
    .Q(u6_remainder[17]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[18]  (.CLK(clk),
    .D(u6_n_144),
    .Q(u6_remainder[18]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[19]  (.CLK(clk),
    .D(u6_n_145),
    .Q(u6_remainder[19]));
 DFFHQx4_ASAP7_75t_SL \u6_remainder_reg[1]  (.CLK(clk),
    .D(u6_n_127),
    .Q(u6_remainder[1]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[20]  (.CLK(clk),
    .D(u6_n_146),
    .Q(u6_remainder[20]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[21]  (.CLK(clk),
    .D(u6_n_147),
    .Q(u6_remainder[21]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[22]  (.CLK(clk),
    .D(u6_n_148),
    .Q(u6_remainder[22]));
 DFFHQx4_ASAP7_75t_SL \u6_remainder_reg[23]  (.CLK(clk),
    .D(u6_n_149),
    .Q(u6_remainder[23]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[2]  (.CLK(clk),
    .D(u6_n_128),
    .Q(u6_remainder[2]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[3]  (.CLK(clk),
    .D(u6_n_129),
    .Q(u6_remainder[3]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[4]  (.CLK(clk),
    .D(u6_n_130),
    .Q(u6_remainder[4]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[5]  (.CLK(clk),
    .D(u6_n_131),
    .Q(u6_remainder[5]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[6]  (.CLK(clk),
    .D(u6_n_132),
    .Q(u6_remainder[6]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[7]  (.CLK(clk),
    .D(u6_n_133),
    .Q(u6_remainder[7]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[8]  (.CLK(clk),
    .D(u6_n_134),
    .Q(u6_remainder[8]));
 DFFHQx4_ASAP7_75t_L \u6_remainder_reg[9]  (.CLK(clk),
    .D(u6_n_135),
    .Q(u6_remainder[9]));
 DFFHQNx1_ASAP7_75t_R \underflow_fmul_r_reg[0]  (.CLK(clk),
    .D(n_2195),
    .QN(underflow_fmul_r[0]));
 DFFHQNx1_ASAP7_75t_R \underflow_fmul_r_reg[1]  (.CLK(clk),
    .D(n_2509),
    .QN(underflow_fmul_r[1]));
 DFFHQNx1_ASAP7_75t_R \underflow_fmul_r_reg[2]  (.CLK(clk),
    .D(n_2539),
    .QN(underflow_fmul_r[2]));
 DFFHQNx1_ASAP7_75t_R underflow_reg (.CLK(clk),
    .D(n_616),
    .QN(underflow));
 DFFHQNx1_ASAP7_75t_R zero_reg (.CLK(clk),
    .D(n_613),
    .QN(zero));
endmodule
