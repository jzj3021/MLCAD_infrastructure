module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire UNCONNECTED;
 wire done_3039;
 wire ld_r;
 wire n_0;
 wire n_1;
 wire n_10;
 wire n_100;
 wire n_1000;
 wire n_10003;
 wire n_10008;
 wire n_1001;
 wire n_10013;
 wire n_10018;
 wire n_1002;
 wire n_10023;
 wire n_10028;
 wire n_1003;
 wire n_10033;
 wire n_1004;
 wire n_1005;
 wire n_1006;
 wire n_1007;
 wire n_1008;
 wire n_1009;
 wire n_101;
 wire n_1010;
 wire n_1011;
 wire n_1012;
 wire n_1013;
 wire n_1014;
 wire n_1015;
 wire n_1016;
 wire n_1017;
 wire n_1018;
 wire n_1019;
 wire n_102;
 wire n_1020;
 wire n_1021;
 wire n_1022;
 wire n_1024;
 wire n_1025;
 wire n_1026;
 wire n_1027;
 wire n_1028;
 wire n_1029;
 wire n_103;
 wire n_1030;
 wire n_1031;
 wire n_1032;
 wire n_1033;
 wire n_1034;
 wire n_1035;
 wire n_1036;
 wire n_1037;
 wire n_1038;
 wire n_1039;
 wire n_104;
 wire n_1040;
 wire n_1041;
 wire n_1042;
 wire n_1043;
 wire n_1044;
 wire n_1045;
 wire n_1046;
 wire n_1047;
 wire n_1048;
 wire n_1049;
 wire n_105;
 wire n_1050;
 wire n_1051;
 wire n_1052;
 wire n_1053;
 wire n_1054;
 wire n_1055;
 wire n_1056;
 wire n_1057;
 wire n_1058;
 wire n_1059;
 wire n_106;
 wire n_1060;
 wire n_1061;
 wire n_1062;
 wire n_1063;
 wire n_1064;
 wire n_1065;
 wire n_1066;
 wire n_1067;
 wire n_1068;
 wire n_1069;
 wire n_107;
 wire n_1070;
 wire n_1071;
 wire n_1072;
 wire n_1073;
 wire n_1074;
 wire n_1075;
 wire n_1076;
 wire n_1077;
 wire n_1078;
 wire n_1079;
 wire n_108;
 wire n_1080;
 wire n_1081;
 wire n_1082;
 wire n_1083;
 wire n_1084;
 wire n_1085;
 wire n_1086;
 wire n_1087;
 wire n_1088;
 wire n_1089;
 wire n_109;
 wire n_1090;
 wire n_1091;
 wire n_1092;
 wire n_1093;
 wire n_1094;
 wire n_1095;
 wire n_1096;
 wire n_1097;
 wire n_1098;
 wire n_1099;
 wire n_11;
 wire n_110;
 wire n_1100;
 wire n_1101;
 wire n_1102;
 wire n_1103;
 wire n_1104;
 wire n_1105;
 wire n_1106;
 wire n_1107;
 wire n_1108;
 wire n_1109;
 wire n_111;
 wire n_1110;
 wire n_1111;
 wire n_1112;
 wire n_1113;
 wire n_1114;
 wire n_1115;
 wire n_1116;
 wire n_1117;
 wire n_1118;
 wire n_1119;
 wire n_112;
 wire n_1120;
 wire n_1121;
 wire n_1122;
 wire n_1123;
 wire n_1124;
 wire n_1125;
 wire n_1126;
 wire n_1127;
 wire n_1128;
 wire n_1129;
 wire n_113;
 wire n_1130;
 wire n_1131;
 wire n_1132;
 wire n_1133;
 wire n_1134;
 wire n_11346;
 wire n_1135;
 wire n_1136;
 wire n_1137;
 wire n_11371;
 wire n_1138;
 wire n_1139;
 wire n_114;
 wire n_1140;
 wire n_11401;
 wire n_1141;
 wire n_1142;
 wire n_1143;
 wire n_11435;
 wire n_1144;
 wire n_1145;
 wire n_11457;
 wire n_1146;
 wire n_1147;
 wire n_1148;
 wire n_11482;
 wire n_1149;
 wire n_1150;
 wire n_11507;
 wire n_1151;
 wire n_11516;
 wire n_11517;
 wire n_11518;
 wire n_1152;
 wire n_11520;
 wire n_11521;
 wire n_11524;
 wire n_1153;
 wire n_1154;
 wire n_1155;
 wire n_1156;
 wire n_1157;
 wire n_1158;
 wire n_1159;
 wire n_116;
 wire n_1160;
 wire n_1161;
 wire n_1162;
 wire n_1163;
 wire n_1164;
 wire n_1165;
 wire n_1166;
 wire n_1167;
 wire n_1168;
 wire n_1169;
 wire n_117;
 wire n_1170;
 wire n_1171;
 wire n_1172;
 wire n_1173;
 wire n_1174;
 wire n_1175;
 wire n_1176;
 wire n_1177;
 wire n_1178;
 wire n_1179;
 wire n_1180;
 wire n_1181;
 wire n_1182;
 wire n_1183;
 wire n_1184;
 wire n_1185;
 wire n_1186;
 wire n_1187;
 wire n_1188;
 wire n_1189;
 wire n_119;
 wire n_1190;
 wire n_1192;
 wire n_1193;
 wire n_1194;
 wire n_1195;
 wire n_1196;
 wire n_1197;
 wire n_1198;
 wire n_1199;
 wire n_12;
 wire n_120;
 wire n_1200;
 wire n_1201;
 wire n_1202;
 wire n_1203;
 wire n_1204;
 wire n_1205;
 wire n_1206;
 wire n_1207;
 wire n_1208;
 wire n_1209;
 wire n_121;
 wire n_1210;
 wire n_1211;
 wire n_1212;
 wire n_1213;
 wire n_1214;
 wire n_1215;
 wire n_1216;
 wire n_1217;
 wire n_1218;
 wire n_1219;
 wire n_122;
 wire n_1220;
 wire n_1221;
 wire n_1222;
 wire n_1223;
 wire n_1224;
 wire n_1225;
 wire n_1226;
 wire n_1227;
 wire n_1228;
 wire n_1229;
 wire n_1230;
 wire n_1231;
 wire n_1232;
 wire n_1233;
 wire n_1234;
 wire n_1235;
 wire n_1236;
 wire n_1237;
 wire n_1238;
 wire n_1239;
 wire n_1240;
 wire n_1241;
 wire n_1242;
 wire n_1243;
 wire n_1244;
 wire n_1245;
 wire n_1246;
 wire n_1247;
 wire n_1248;
 wire n_1249;
 wire n_125;
 wire n_1250;
 wire n_1251;
 wire n_1252;
 wire n_1253;
 wire n_1254;
 wire n_1255;
 wire n_1256;
 wire n_1257;
 wire n_1258;
 wire n_1259;
 wire n_126;
 wire n_1260;
 wire n_1261;
 wire n_1262;
 wire n_1263;
 wire n_1264;
 wire n_1265;
 wire n_1266;
 wire n_1267;
 wire n_1268;
 wire n_1269;
 wire n_127;
 wire n_1270;
 wire n_1271;
 wire n_1272;
 wire n_1273;
 wire n_1274;
 wire n_1275;
 wire n_1276;
 wire n_1277;
 wire n_1278;
 wire n_1279;
 wire n_128;
 wire n_1280;
 wire n_1281;
 wire n_12816;
 wire n_1282;
 wire n_1283;
 wire n_1284;
 wire n_1285;
 wire n_1286;
 wire n_1287;
 wire n_1288;
 wire n_1289;
 wire n_129;
 wire n_1290;
 wire n_1291;
 wire n_1292;
 wire n_1293;
 wire n_1294;
 wire n_1295;
 wire n_1296;
 wire n_1297;
 wire n_1298;
 wire n_1299;
 wire n_13;
 wire n_130;
 wire n_1300;
 wire n_1301;
 wire n_1302;
 wire n_1303;
 wire n_1304;
 wire n_1305;
 wire n_1306;
 wire n_1307;
 wire n_1308;
 wire n_1309;
 wire n_131;
 wire n_1310;
 wire n_1311;
 wire n_1312;
 wire n_1313;
 wire n_1314;
 wire n_1315;
 wire n_1316;
 wire n_1317;
 wire n_1318;
 wire n_1319;
 wire n_1320;
 wire n_1321;
 wire n_1322;
 wire n_1323;
 wire n_1324;
 wire n_1325;
 wire n_1326;
 wire n_1327;
 wire n_1328;
 wire n_1329;
 wire n_1330;
 wire n_1331;
 wire n_1332;
 wire n_1333;
 wire n_1334;
 wire n_1335;
 wire n_1336;
 wire n_1337;
 wire n_1338;
 wire n_1339;
 wire n_134;
 wire n_1340;
 wire n_1341;
 wire n_1342;
 wire n_1343;
 wire n_1344;
 wire n_1345;
 wire n_1346;
 wire n_1348;
 wire n_1349;
 wire n_135;
 wire n_1350;
 wire n_1351;
 wire n_1352;
 wire n_1353;
 wire n_1354;
 wire n_1355;
 wire n_1356;
 wire n_1357;
 wire n_1358;
 wire n_1359;
 wire n_136;
 wire n_1360;
 wire n_1361;
 wire n_1362;
 wire n_1363;
 wire n_1364;
 wire n_1365;
 wire n_1366;
 wire n_1367;
 wire n_1368;
 wire n_1369;
 wire n_137;
 wire n_1370;
 wire n_1371;
 wire n_1372;
 wire n_1373;
 wire n_1374;
 wire n_1375;
 wire n_1376;
 wire n_1377;
 wire n_1378;
 wire n_1379;
 wire n_138;
 wire n_1380;
 wire n_1381;
 wire n_1382;
 wire n_1383;
 wire n_1384;
 wire n_1385;
 wire n_1386;
 wire n_1387;
 wire n_1389;
 wire n_1390;
 wire n_1391;
 wire n_1392;
 wire n_1393;
 wire n_1394;
 wire n_1395;
 wire n_1396;
 wire n_1397;
 wire n_1398;
 wire n_1399;
 wire n_14;
 wire n_1400;
 wire n_1401;
 wire n_1402;
 wire n_1403;
 wire n_1404;
 wire n_1405;
 wire n_1406;
 wire n_1407;
 wire n_1408;
 wire n_1409;
 wire n_1410;
 wire n_1411;
 wire n_1412;
 wire n_1413;
 wire n_1414;
 wire n_1415;
 wire n_1416;
 wire n_1417;
 wire n_1418;
 wire n_1419;
 wire n_1420;
 wire n_1421;
 wire n_1422;
 wire n_1423;
 wire n_1424;
 wire n_1425;
 wire n_1426;
 wire n_1427;
 wire n_1429;
 wire n_143;
 wire n_1430;
 wire n_1431;
 wire n_1432;
 wire n_1433;
 wire n_1434;
 wire n_1435;
 wire n_1436;
 wire n_1437;
 wire n_1438;
 wire n_1439;
 wire n_144;
 wire n_1440;
 wire n_1441;
 wire n_1442;
 wire n_1443;
 wire n_1444;
 wire n_1445;
 wire n_1446;
 wire n_1447;
 wire n_1448;
 wire n_1449;
 wire n_145;
 wire n_1450;
 wire n_1451;
 wire n_1452;
 wire n_1453;
 wire n_1454;
 wire n_1455;
 wire n_1456;
 wire n_1457;
 wire n_1458;
 wire n_1459;
 wire n_1460;
 wire n_1461;
 wire n_1462;
 wire n_1463;
 wire n_1464;
 wire n_1465;
 wire n_1466;
 wire n_1467;
 wire n_1469;
 wire n_147;
 wire n_1470;
 wire n_1471;
 wire n_1472;
 wire n_1473;
 wire n_1474;
 wire n_1475;
 wire n_1476;
 wire n_1477;
 wire n_1478;
 wire n_1479;
 wire n_148;
 wire n_1480;
 wire n_1481;
 wire n_1482;
 wire n_1483;
 wire n_1484;
 wire n_1485;
 wire n_1486;
 wire n_1487;
 wire n_149;
 wire n_1490;
 wire n_1491;
 wire n_1492;
 wire n_1493;
 wire n_1494;
 wire n_1495;
 wire n_1496;
 wire n_1497;
 wire n_1498;
 wire n_1499;
 wire n_15;
 wire n_150;
 wire n_1500;
 wire n_1501;
 wire n_1502;
 wire n_1503;
 wire n_1504;
 wire n_1505;
 wire n_1506;
 wire n_1507;
 wire n_1509;
 wire n_151;
 wire n_1510;
 wire n_1511;
 wire n_1512;
 wire n_1513;
 wire n_1517;
 wire n_1518;
 wire n_1519;
 wire n_152;
 wire n_1522;
 wire n_1523;
 wire n_1524;
 wire n_1525;
 wire n_1526;
 wire n_1527;
 wire n_1528;
 wire n_1529;
 wire n_153;
 wire n_1530;
 wire n_1531;
 wire n_1532;
 wire n_1533;
 wire n_1534;
 wire n_1535;
 wire n_1536;
 wire n_1537;
 wire n_1538;
 wire n_154;
 wire n_1540;
 wire n_1541;
 wire n_1542;
 wire n_1543;
 wire n_1544;
 wire n_1545;
 wire n_1546;
 wire n_1547;
 wire n_1548;
 wire n_1549;
 wire n_1550;
 wire n_1551;
 wire n_1552;
 wire n_1553;
 wire n_1554;
 wire n_1555;
 wire n_1556;
 wire n_1557;
 wire n_1558;
 wire n_1559;
 wire n_156;
 wire n_1560;
 wire n_1561;
 wire n_1562;
 wire n_1565;
 wire n_1566;
 wire n_1567;
 wire n_1568;
 wire n_1569;
 wire n_157;
 wire n_1570;
 wire n_1571;
 wire n_1572;
 wire n_1573;
 wire n_1575;
 wire n_1576;
 wire n_1577;
 wire n_1578;
 wire n_158;
 wire n_1580;
 wire n_1581;
 wire n_1582;
 wire n_1583;
 wire n_1584;
 wire n_1585;
 wire n_1586;
 wire n_1587;
 wire n_1588;
 wire n_1589;
 wire n_159;
 wire n_1590;
 wire n_1591;
 wire n_1592;
 wire n_1593;
 wire n_1594;
 wire n_1595;
 wire n_1596;
 wire n_1597;
 wire n_1598;
 wire n_1599;
 wire n_16;
 wire n_1600;
 wire n_1601;
 wire n_1602;
 wire n_1603;
 wire n_1604;
 wire n_1605;
 wire n_1606;
 wire n_1607;
 wire n_1608;
 wire n_1609;
 wire n_161;
 wire n_1610;
 wire n_1611;
 wire n_1612;
 wire n_1613;
 wire n_1614;
 wire n_1615;
 wire n_1616;
 wire n_1617;
 wire n_1618;
 wire n_1619;
 wire n_1620;
 wire n_1621;
 wire n_1622;
 wire n_1623;
 wire n_1624;
 wire n_1625;
 wire n_1626;
 wire n_1627;
 wire n_1628;
 wire n_1629;
 wire n_163;
 wire n_1632;
 wire n_1633;
 wire n_1634;
 wire n_1635;
 wire n_1636;
 wire n_1637;
 wire n_1638;
 wire n_1639;
 wire n_164;
 wire n_1640;
 wire n_1641;
 wire n_1642;
 wire n_1643;
 wire n_1644;
 wire n_1645;
 wire n_1646;
 wire n_1647;
 wire n_165;
 wire n_1650;
 wire n_1651;
 wire n_1652;
 wire n_1653;
 wire n_1654;
 wire n_1655;
 wire n_1656;
 wire n_1657;
 wire n_1658;
 wire n_1659;
 wire n_166;
 wire n_1660;
 wire n_1662;
 wire n_1663;
 wire n_1664;
 wire n_1665;
 wire n_1666;
 wire n_1667;
 wire n_1668;
 wire n_1669;
 wire n_167;
 wire n_1670;
 wire n_1671;
 wire n_1672;
 wire n_1673;
 wire n_1674;
 wire n_1675;
 wire n_1676;
 wire n_1677;
 wire n_1678;
 wire n_1679;
 wire n_168;
 wire n_1680;
 wire n_1681;
 wire n_1682;
 wire n_1683;
 wire n_1686;
 wire n_1687;
 wire n_1688;
 wire n_1689;
 wire n_169;
 wire n_1690;
 wire n_1691;
 wire n_1693;
 wire n_1694;
 wire n_1695;
 wire n_1696;
 wire n_1697;
 wire n_1698;
 wire n_1699;
 wire n_17;
 wire n_1700;
 wire n_1701;
 wire n_1702;
 wire n_1703;
 wire n_1704;
 wire n_1705;
 wire n_1706;
 wire n_1707;
 wire n_1708;
 wire n_1709;
 wire n_1710;
 wire n_1711;
 wire n_1712;
 wire n_1713;
 wire n_1714;
 wire n_1715;
 wire n_1716;
 wire n_1717;
 wire n_1718;
 wire n_1719;
 wire n_172;
 wire n_1720;
 wire n_1721;
 wire n_1722;
 wire n_1723;
 wire n_1724;
 wire n_1725;
 wire n_1726;
 wire n_1727;
 wire n_1728;
 wire n_1729;
 wire n_173;
 wire n_1730;
 wire n_1731;
 wire n_1732;
 wire n_1733;
 wire n_1734;
 wire n_1735;
 wire n_1736;
 wire n_1737;
 wire n_1738;
 wire n_1739;
 wire n_174;
 wire n_1740;
 wire n_1741;
 wire n_1742;
 wire n_1743;
 wire n_1744;
 wire n_1745;
 wire n_1746;
 wire n_1747;
 wire n_1748;
 wire n_1749;
 wire n_175;
 wire n_1750;
 wire n_1751;
 wire n_1752;
 wire n_1753;
 wire n_1754;
 wire n_1755;
 wire n_1756;
 wire n_1757;
 wire n_1758;
 wire n_1759;
 wire n_176;
 wire n_1760;
 wire n_1761;
 wire n_1762;
 wire n_1763;
 wire n_1764;
 wire n_1765;
 wire n_1766;
 wire n_1767;
 wire n_1768;
 wire n_1769;
 wire n_177;
 wire n_1770;
 wire n_1771;
 wire n_1772;
 wire n_1773;
 wire n_1774;
 wire n_1775;
 wire n_1776;
 wire n_1777;
 wire n_1778;
 wire n_1779;
 wire n_178;
 wire n_1780;
 wire n_1781;
 wire n_1782;
 wire n_1783;
 wire n_1784;
 wire n_1785;
 wire n_1786;
 wire n_1787;
 wire n_1788;
 wire n_1789;
 wire n_179;
 wire n_1790;
 wire n_1791;
 wire n_1792;
 wire n_1793;
 wire n_1794;
 wire n_1795;
 wire n_1796;
 wire n_1797;
 wire n_18;
 wire n_180;
 wire n_1800;
 wire n_1801;
 wire n_1802;
 wire n_1803;
 wire n_1804;
 wire n_1805;
 wire n_1806;
 wire n_1807;
 wire n_1808;
 wire n_1809;
 wire n_181;
 wire n_1810;
 wire n_1812;
 wire n_1813;
 wire n_1814;
 wire n_1815;
 wire n_1817;
 wire n_1818;
 wire n_1819;
 wire n_182;
 wire n_1820;
 wire n_1821;
 wire n_1822;
 wire n_1823;
 wire n_1824;
 wire n_1825;
 wire n_1826;
 wire n_1827;
 wire n_1828;
 wire n_1829;
 wire n_183;
 wire n_1830;
 wire n_1831;
 wire n_1832;
 wire n_1833;
 wire n_1834;
 wire n_1835;
 wire n_1836;
 wire n_1837;
 wire n_1838;
 wire n_1839;
 wire n_184;
 wire n_1840;
 wire n_1843;
 wire n_1844;
 wire n_1845;
 wire n_1846;
 wire n_1850;
 wire n_1851;
 wire n_1852;
 wire n_1853;
 wire n_1855;
 wire n_1856;
 wire n_1857;
 wire n_1859;
 wire n_186;
 wire n_1860;
 wire n_1862;
 wire n_1865;
 wire n_1866;
 wire n_1867;
 wire n_1869;
 wire n_187;
 wire n_1870;
 wire n_1871;
 wire n_1873;
 wire n_1874;
 wire n_1876;
 wire n_1877;
 wire n_1878;
 wire n_1879;
 wire n_1880;
 wire n_1884;
 wire n_1886;
 wire n_1888;
 wire n_189;
 wire n_1890;
 wire n_1891;
 wire n_1893;
 wire n_1894;
 wire n_1895;
 wire n_1896;
 wire n_19;
 wire n_190;
 wire n_1900;
 wire n_1901;
 wire n_1902;
 wire n_1903;
 wire n_1904;
 wire n_1905;
 wire n_1908;
 wire n_1909;
 wire n_191;
 wire n_1910;
 wire n_1912;
 wire n_1913;
 wire n_1914;
 wire n_1915;
 wire n_1916;
 wire n_1917;
 wire n_1918;
 wire n_1921;
 wire n_1923;
 wire n_1924;
 wire n_1925;
 wire n_1926;
 wire n_1928;
 wire n_1929;
 wire n_193;
 wire n_1930;
 wire n_1933;
 wire n_1934;
 wire n_1935;
 wire n_1938;
 wire n_1939;
 wire n_194;
 wire n_1940;
 wire n_1941;
 wire n_1944;
 wire n_1945;
 wire n_1947;
 wire n_1948;
 wire n_1949;
 wire n_195;
 wire n_1950;
 wire n_1952;
 wire n_1953;
 wire n_1954;
 wire n_1955;
 wire n_1957;
 wire n_1958;
 wire n_1959;
 wire n_196;
 wire n_1960;
 wire n_1961;
 wire n_1964;
 wire n_1965;
 wire n_1966;
 wire n_1967;
 wire n_1968;
 wire n_1969;
 wire n_1970;
 wire n_1971;
 wire n_1972;
 wire n_1975;
 wire n_1979;
 wire n_1980;
 wire n_1981;
 wire n_1982;
 wire n_1983;
 wire n_1984;
 wire n_1985;
 wire n_1986;
 wire n_1987;
 wire n_199;
 wire n_1990;
 wire n_1992;
 wire n_1994;
 wire n_1995;
 wire n_2;
 wire n_20;
 wire n_200;
 wire n_2001;
 wire n_2003;
 wire n_2004;
 wire n_2005;
 wire n_2006;
 wire n_2007;
 wire n_2008;
 wire n_2009;
 wire n_2010;
 wire n_2011;
 wire n_2012;
 wire n_2013;
 wire n_2014;
 wire n_2015;
 wire n_2016;
 wire n_2017;
 wire n_2018;
 wire n_2019;
 wire n_202;
 wire n_2020;
 wire n_2022;
 wire n_2023;
 wire n_2024;
 wire n_2026;
 wire n_2028;
 wire n_2029;
 wire n_203;
 wire n_2031;
 wire n_2032;
 wire n_2033;
 wire n_2034;
 wire n_2035;
 wire n_2037;
 wire n_2038;
 wire n_2039;
 wire n_204;
 wire n_2040;
 wire n_2041;
 wire n_2042;
 wire n_2043;
 wire n_2044;
 wire n_2045;
 wire n_2046;
 wire n_2047;
 wire n_2048;
 wire n_2050;
 wire n_2051;
 wire n_2052;
 wire n_2053;
 wire n_2054;
 wire n_2055;
 wire n_2056;
 wire n_2057;
 wire n_2058;
 wire n_2059;
 wire n_206;
 wire n_2060;
 wire n_2061;
 wire n_2062;
 wire n_2063;
 wire n_2064;
 wire n_2065;
 wire n_2066;
 wire n_2067;
 wire n_2068;
 wire n_2069;
 wire n_207;
 wire n_2070;
 wire n_2072;
 wire n_2073;
 wire n_2074;
 wire n_2075;
 wire n_2076;
 wire n_2077;
 wire n_2078;
 wire n_2079;
 wire n_208;
 wire n_2080;
 wire n_2081;
 wire n_2082;
 wire n_2083;
 wire n_2084;
 wire n_2087;
 wire n_2088;
 wire n_2089;
 wire n_209;
 wire n_2090;
 wire n_2091;
 wire n_2092;
 wire n_2094;
 wire n_2095;
 wire n_2096;
 wire n_2097;
 wire n_2098;
 wire n_2099;
 wire n_21;
 wire n_210;
 wire n_2100;
 wire n_2101;
 wire n_2102;
 wire n_2103;
 wire n_2104;
 wire n_2105;
 wire n_2106;
 wire n_2107;
 wire n_2108;
 wire n_211;
 wire n_2110;
 wire n_2111;
 wire n_2112;
 wire n_2113;
 wire n_2114;
 wire n_2115;
 wire n_2116;
 wire n_2117;
 wire n_2118;
 wire n_2119;
 wire n_2120;
 wire n_2121;
 wire n_2122;
 wire n_2123;
 wire n_2124;
 wire n_2125;
 wire n_2126;
 wire n_2127;
 wire n_2128;
 wire n_2129;
 wire n_213;
 wire n_2130;
 wire n_2131;
 wire n_2132;
 wire n_2133;
 wire n_2134;
 wire n_2135;
 wire n_2136;
 wire n_2137;
 wire n_2138;
 wire n_2139;
 wire n_214;
 wire n_2140;
 wire n_2141;
 wire n_2142;
 wire n_2143;
 wire n_2144;
 wire n_2145;
 wire n_2146;
 wire n_2147;
 wire n_2148;
 wire n_2149;
 wire n_215;
 wire n_2150;
 wire n_2151;
 wire n_2152;
 wire n_2153;
 wire n_2154;
 wire n_2155;
 wire n_2156;
 wire n_2157;
 wire n_2158;
 wire n_2159;
 wire n_2160;
 wire n_2161;
 wire n_2162;
 wire n_2163;
 wire n_2164;
 wire n_2165;
 wire n_2166;
 wire n_2167;
 wire n_2168;
 wire n_2169;
 wire n_217;
 wire n_2170;
 wire n_2171;
 wire n_2172;
 wire n_2173;
 wire n_2174;
 wire n_2175;
 wire n_2176;
 wire n_2177;
 wire n_2178;
 wire n_2179;
 wire n_218;
 wire n_2180;
 wire n_2181;
 wire n_2182;
 wire n_2183;
 wire n_2184;
 wire n_2185;
 wire n_2186;
 wire n_2187;
 wire n_2188;
 wire n_2189;
 wire n_219;
 wire n_2190;
 wire n_2191;
 wire n_2192;
 wire n_2193;
 wire n_2194;
 wire n_2195;
 wire n_2196;
 wire n_2197;
 wire n_2198;
 wire n_2199;
 wire n_22;
 wire n_220;
 wire n_2200;
 wire n_2201;
 wire n_2202;
 wire n_2203;
 wire n_2204;
 wire n_2205;
 wire n_2206;
 wire n_2208;
 wire n_2209;
 wire n_221;
 wire n_2210;
 wire n_2211;
 wire n_2212;
 wire n_2213;
 wire n_2214;
 wire n_2215;
 wire n_2216;
 wire n_2217;
 wire n_2218;
 wire n_2219;
 wire n_222;
 wire n_2220;
 wire n_2221;
 wire n_2222;
 wire n_2223;
 wire n_2224;
 wire n_2225;
 wire n_2226;
 wire n_2227;
 wire n_2228;
 wire n_2229;
 wire n_223;
 wire n_2230;
 wire n_2231;
 wire n_2232;
 wire n_2233;
 wire n_2234;
 wire n_2235;
 wire n_2236;
 wire n_2237;
 wire n_2238;
 wire n_2239;
 wire n_224;
 wire n_2240;
 wire n_2241;
 wire n_2242;
 wire n_2243;
 wire n_2244;
 wire n_2245;
 wire n_2246;
 wire n_2247;
 wire n_2248;
 wire n_2249;
 wire n_225;
 wire n_2250;
 wire n_2251;
 wire n_2252;
 wire n_2253;
 wire n_2254;
 wire n_2255;
 wire n_2256;
 wire n_2257;
 wire n_2258;
 wire n_2259;
 wire n_226;
 wire n_2260;
 wire n_2261;
 wire n_2262;
 wire n_2263;
 wire n_2264;
 wire n_2265;
 wire n_2266;
 wire n_2267;
 wire n_2268;
 wire n_2269;
 wire n_227;
 wire n_2270;
 wire n_2271;
 wire n_2272;
 wire n_2273;
 wire n_2274;
 wire n_2275;
 wire n_2276;
 wire n_2277;
 wire n_2278;
 wire n_2279;
 wire n_228;
 wire n_2280;
 wire n_2281;
 wire n_2282;
 wire n_2283;
 wire n_2284;
 wire n_2285;
 wire n_2286;
 wire n_2287;
 wire n_2288;
 wire n_2289;
 wire n_229;
 wire n_2290;
 wire n_2291;
 wire n_2292;
 wire n_2293;
 wire n_2294;
 wire n_2295;
 wire n_2296;
 wire n_2297;
 wire n_2298;
 wire n_2299;
 wire n_23;
 wire n_230;
 wire n_2300;
 wire n_2301;
 wire n_2302;
 wire n_2303;
 wire n_2304;
 wire n_2305;
 wire n_2306;
 wire n_2307;
 wire n_2308;
 wire n_2309;
 wire n_231;
 wire n_2310;
 wire n_2311;
 wire n_2312;
 wire n_2313;
 wire n_2314;
 wire n_2315;
 wire n_2316;
 wire n_2317;
 wire n_2318;
 wire n_2319;
 wire n_232;
 wire n_2320;
 wire n_2321;
 wire n_2322;
 wire n_2323;
 wire n_2324;
 wire n_2325;
 wire n_2326;
 wire n_2327;
 wire n_2328;
 wire n_2329;
 wire n_233;
 wire n_2330;
 wire n_2331;
 wire n_2332;
 wire n_2333;
 wire n_2334;
 wire n_2335;
 wire n_2336;
 wire n_2337;
 wire n_2338;
 wire n_2339;
 wire n_234;
 wire n_2340;
 wire n_2341;
 wire n_2342;
 wire n_2343;
 wire n_2344;
 wire n_2345;
 wire n_2346;
 wire n_2347;
 wire n_2348;
 wire n_2349;
 wire n_235;
 wire n_2350;
 wire n_2351;
 wire n_2352;
 wire n_2353;
 wire n_2354;
 wire n_2355;
 wire n_2356;
 wire n_2357;
 wire n_2358;
 wire n_2359;
 wire n_236;
 wire n_2360;
 wire n_2361;
 wire n_2362;
 wire n_2363;
 wire n_2364;
 wire n_2365;
 wire n_2366;
 wire n_2367;
 wire n_2368;
 wire n_2369;
 wire n_237;
 wire n_2370;
 wire n_2371;
 wire n_2372;
 wire n_2373;
 wire n_2374;
 wire n_2375;
 wire n_2376;
 wire n_2377;
 wire n_2378;
 wire n_2379;
 wire n_238;
 wire n_2380;
 wire n_2381;
 wire n_2382;
 wire n_2383;
 wire n_2384;
 wire n_2385;
 wire n_2386;
 wire n_2387;
 wire n_2388;
 wire n_2389;
 wire n_239;
 wire n_2390;
 wire n_2392;
 wire n_2393;
 wire n_2394;
 wire n_2395;
 wire n_2396;
 wire n_2397;
 wire n_2398;
 wire n_2399;
 wire n_24;
 wire n_240;
 wire n_2400;
 wire n_2401;
 wire n_2402;
 wire n_2403;
 wire n_2404;
 wire n_241;
 wire n_2410;
 wire n_2411;
 wire n_2412;
 wire n_2413;
 wire n_2414;
 wire n_2415;
 wire n_2416;
 wire n_2417;
 wire n_2418;
 wire n_2419;
 wire n_242;
 wire n_2420;
 wire n_2421;
 wire n_2422;
 wire n_2423;
 wire n_2424;
 wire n_2425;
 wire n_2427;
 wire n_2428;
 wire n_2429;
 wire n_243;
 wire n_2430;
 wire n_2431;
 wire n_2432;
 wire n_2433;
 wire n_2434;
 wire n_2435;
 wire n_2436;
 wire n_2437;
 wire n_2438;
 wire n_2439;
 wire n_2440;
 wire n_2441;
 wire n_2442;
 wire n_2443;
 wire n_2444;
 wire n_2445;
 wire n_2446;
 wire n_2447;
 wire n_2448;
 wire n_2449;
 wire n_245;
 wire n_2450;
 wire n_2451;
 wire n_2452;
 wire n_2453;
 wire n_2455;
 wire n_2456;
 wire n_2457;
 wire n_2458;
 wire n_2459;
 wire n_2460;
 wire n_2461;
 wire n_2462;
 wire n_2463;
 wire n_2464;
 wire n_2465;
 wire n_2466;
 wire n_2467;
 wire n_2468;
 wire n_2469;
 wire n_247;
 wire n_2470;
 wire n_2471;
 wire n_2472;
 wire n_2473;
 wire n_2474;
 wire n_2475;
 wire n_2476;
 wire n_2477;
 wire n_2478;
 wire n_2479;
 wire n_2480;
 wire n_2481;
 wire n_2482;
 wire n_2483;
 wire n_2484;
 wire n_2485;
 wire n_2486;
 wire n_2487;
 wire n_2488;
 wire n_2489;
 wire n_2490;
 wire n_2491;
 wire n_2492;
 wire n_2494;
 wire n_2495;
 wire n_2496;
 wire n_2497;
 wire n_2499;
 wire n_25;
 wire n_2500;
 wire n_2501;
 wire n_2502;
 wire n_2503;
 wire n_2504;
 wire n_2505;
 wire n_2506;
 wire n_2507;
 wire n_2508;
 wire n_2509;
 wire n_2510;
 wire n_2511;
 wire n_2512;
 wire n_2513;
 wire n_2514;
 wire n_2515;
 wire n_2517;
 wire n_2518;
 wire n_2519;
 wire n_252;
 wire n_2520;
 wire n_2521;
 wire n_2522;
 wire n_2523;
 wire n_2524;
 wire n_2525;
 wire n_2526;
 wire n_2527;
 wire n_2528;
 wire n_2529;
 wire n_253;
 wire n_2530;
 wire n_2531;
 wire n_2532;
 wire n_2533;
 wire n_2534;
 wire n_2535;
 wire n_2536;
 wire n_2537;
 wire n_2538;
 wire n_2539;
 wire n_254;
 wire n_2540;
 wire n_2541;
 wire n_2542;
 wire n_2543;
 wire n_2544;
 wire n_2545;
 wire n_2546;
 wire n_2547;
 wire n_2548;
 wire n_2549;
 wire n_255;
 wire n_2550;
 wire n_2551;
 wire n_2552;
 wire n_2553;
 wire n_2554;
 wire n_2555;
 wire n_2556;
 wire n_2557;
 wire n_2558;
 wire n_2559;
 wire n_256;
 wire n_2560;
 wire n_2561;
 wire n_2562;
 wire n_2563;
 wire n_2564;
 wire n_2565;
 wire n_2566;
 wire n_2567;
 wire n_2568;
 wire n_2569;
 wire n_2570;
 wire n_2571;
 wire n_2572;
 wire n_2573;
 wire n_2574;
 wire n_2575;
 wire n_2576;
 wire n_2577;
 wire n_2578;
 wire n_2579;
 wire n_258;
 wire n_2580;
 wire n_2581;
 wire n_2582;
 wire n_2583;
 wire n_2584;
 wire n_2585;
 wire n_2586;
 wire n_2587;
 wire n_2588;
 wire n_2589;
 wire n_259;
 wire n_2590;
 wire n_2591;
 wire n_2592;
 wire n_2593;
 wire n_2594;
 wire n_2595;
 wire n_2596;
 wire n_2597;
 wire n_2598;
 wire n_2599;
 wire n_26;
 wire n_260;
 wire n_2600;
 wire n_2601;
 wire n_2602;
 wire n_2603;
 wire n_2604;
 wire n_2605;
 wire n_2606;
 wire n_2607;
 wire n_2608;
 wire n_2609;
 wire n_261;
 wire n_2610;
 wire n_2611;
 wire n_2612;
 wire n_2613;
 wire n_2614;
 wire n_2615;
 wire n_2616;
 wire n_2617;
 wire n_2618;
 wire n_2619;
 wire n_2620;
 wire n_2621;
 wire n_2622;
 wire n_2623;
 wire n_2624;
 wire n_2625;
 wire n_2626;
 wire n_2627;
 wire n_2628;
 wire n_2629;
 wire n_263;
 wire n_2630;
 wire n_2631;
 wire n_2632;
 wire n_2633;
 wire n_2634;
 wire n_2635;
 wire n_2636;
 wire n_2637;
 wire n_2638;
 wire n_2639;
 wire n_264;
 wire n_2640;
 wire n_2642;
 wire n_2643;
 wire n_2644;
 wire n_2645;
 wire n_2646;
 wire n_2647;
 wire n_2648;
 wire n_2649;
 wire n_265;
 wire n_2650;
 wire n_2651;
 wire n_2652;
 wire n_2653;
 wire n_2654;
 wire n_2655;
 wire n_2656;
 wire n_2657;
 wire n_2658;
 wire n_2659;
 wire n_266;
 wire n_2660;
 wire n_2661;
 wire n_2662;
 wire n_2663;
 wire n_2664;
 wire n_2665;
 wire n_2666;
 wire n_2667;
 wire n_2668;
 wire n_267;
 wire n_2670;
 wire n_2671;
 wire n_2672;
 wire n_2673;
 wire n_2674;
 wire n_2675;
 wire n_2676;
 wire n_2677;
 wire n_2678;
 wire n_2679;
 wire n_268;
 wire n_2680;
 wire n_2681;
 wire n_2682;
 wire n_2683;
 wire n_2684;
 wire n_2685;
 wire n_2686;
 wire n_2687;
 wire n_2688;
 wire n_2689;
 wire n_269;
 wire n_2690;
 wire n_2691;
 wire n_2692;
 wire n_2693;
 wire n_2694;
 wire n_2695;
 wire n_2696;
 wire n_2697;
 wire n_2698;
 wire n_2699;
 wire n_27;
 wire n_270;
 wire n_2700;
 wire n_2701;
 wire n_2702;
 wire n_2703;
 wire n_2704;
 wire n_2705;
 wire n_2706;
 wire n_2707;
 wire n_2708;
 wire n_2709;
 wire n_271;
 wire n_2710;
 wire n_2711;
 wire n_2712;
 wire n_2713;
 wire n_2714;
 wire n_2715;
 wire n_2716;
 wire n_2717;
 wire n_2718;
 wire n_2719;
 wire n_272;
 wire n_2720;
 wire n_2721;
 wire n_2722;
 wire n_2723;
 wire n_2724;
 wire n_2725;
 wire n_2726;
 wire n_2727;
 wire n_2728;
 wire n_2729;
 wire n_2730;
 wire n_2731;
 wire n_2732;
 wire n_2733;
 wire n_2734;
 wire n_2735;
 wire n_2736;
 wire n_2737;
 wire n_2738;
 wire n_2739;
 wire n_2740;
 wire n_2741;
 wire n_2742;
 wire n_2743;
 wire n_2744;
 wire n_2745;
 wire n_2746;
 wire n_2747;
 wire n_2748;
 wire n_2749;
 wire n_2750;
 wire n_2751;
 wire n_2752;
 wire n_2753;
 wire n_2754;
 wire n_2755;
 wire n_2756;
 wire n_2757;
 wire n_2758;
 wire n_2759;
 wire n_2760;
 wire n_2761;
 wire n_2762;
 wire n_2763;
 wire n_2764;
 wire n_2765;
 wire n_2766;
 wire n_2767;
 wire n_2768;
 wire n_2769;
 wire n_2770;
 wire n_2771;
 wire n_2772;
 wire n_2773;
 wire n_2774;
 wire n_2775;
 wire n_2776;
 wire n_2777;
 wire n_2778;
 wire n_2779;
 wire n_278;
 wire n_2780;
 wire n_2781;
 wire n_2782;
 wire n_2783;
 wire n_2784;
 wire n_2785;
 wire n_2786;
 wire n_2787;
 wire n_2788;
 wire n_2789;
 wire n_279;
 wire n_2790;
 wire n_2791;
 wire n_2792;
 wire n_2793;
 wire n_2794;
 wire n_2795;
 wire n_2796;
 wire n_2797;
 wire n_2798;
 wire n_2799;
 wire n_28;
 wire n_280;
 wire n_2800;
 wire n_2801;
 wire n_2802;
 wire n_2803;
 wire n_2804;
 wire n_2805;
 wire n_2806;
 wire n_2807;
 wire n_2808;
 wire n_2809;
 wire n_281;
 wire n_2811;
 wire n_2813;
 wire n_2814;
 wire n_2815;
 wire n_2816;
 wire n_2817;
 wire n_2818;
 wire n_2819;
 wire n_282;
 wire n_2820;
 wire n_2821;
 wire n_2822;
 wire n_2823;
 wire n_2824;
 wire n_2825;
 wire n_2826;
 wire n_2827;
 wire n_2828;
 wire n_2829;
 wire n_283;
 wire n_2830;
 wire n_2831;
 wire n_2832;
 wire n_2833;
 wire n_2834;
 wire n_2835;
 wire n_2837;
 wire n_2838;
 wire n_2839;
 wire n_2840;
 wire n_2841;
 wire n_2842;
 wire n_2843;
 wire n_2844;
 wire n_2845;
 wire n_2846;
 wire n_2847;
 wire n_2848;
 wire n_2849;
 wire n_285;
 wire n_2850;
 wire n_2851;
 wire n_2852;
 wire n_2853;
 wire n_2854;
 wire n_2855;
 wire n_2856;
 wire n_2857;
 wire n_2858;
 wire n_2859;
 wire n_2860;
 wire n_2861;
 wire n_2862;
 wire n_2863;
 wire n_2864;
 wire n_2865;
 wire n_2866;
 wire n_2867;
 wire n_2868;
 wire n_2869;
 wire n_2870;
 wire n_2871;
 wire n_2872;
 wire n_2873;
 wire n_2874;
 wire n_2875;
 wire n_2876;
 wire n_2877;
 wire n_2878;
 wire n_2879;
 wire n_2880;
 wire n_2881;
 wire n_2882;
 wire n_2883;
 wire n_2884;
 wire n_2885;
 wire n_2886;
 wire n_2887;
 wire n_2888;
 wire n_2889;
 wire n_289;
 wire n_2890;
 wire n_2891;
 wire n_2892;
 wire n_2893;
 wire n_2894;
 wire n_2895;
 wire n_2896;
 wire n_2897;
 wire n_2898;
 wire n_2899;
 wire n_29;
 wire n_290;
 wire n_2900;
 wire n_2901;
 wire n_2902;
 wire n_2903;
 wire n_2904;
 wire n_2905;
 wire n_2906;
 wire n_2907;
 wire n_2908;
 wire n_2909;
 wire n_291;
 wire n_2910;
 wire n_2911;
 wire n_2912;
 wire n_2913;
 wire n_2914;
 wire n_2915;
 wire n_2916;
 wire n_2917;
 wire n_2918;
 wire n_2919;
 wire n_292;
 wire n_2920;
 wire n_2921;
 wire n_2922;
 wire n_2923;
 wire n_2924;
 wire n_2925;
 wire n_2926;
 wire n_2927;
 wire n_2928;
 wire n_2929;
 wire n_293;
 wire n_2930;
 wire n_2931;
 wire n_2932;
 wire n_2933;
 wire n_2934;
 wire n_2935;
 wire n_2936;
 wire n_2937;
 wire n_2938;
 wire n_2939;
 wire n_294;
 wire n_2940;
 wire n_2941;
 wire n_2942;
 wire n_2943;
 wire n_2944;
 wire n_2945;
 wire n_2946;
 wire n_2947;
 wire n_2948;
 wire n_2949;
 wire n_295;
 wire n_2950;
 wire n_2951;
 wire n_2952;
 wire n_2953;
 wire n_2954;
 wire n_2955;
 wire n_2956;
 wire n_2957;
 wire n_2958;
 wire n_2959;
 wire n_296;
 wire n_2960;
 wire n_2961;
 wire n_2962;
 wire n_2963;
 wire n_2964;
 wire n_2965;
 wire n_2966;
 wire n_2967;
 wire n_2968;
 wire n_2969;
 wire n_2970;
 wire n_2971;
 wire n_2972;
 wire n_2973;
 wire n_2974;
 wire n_2975;
 wire n_2976;
 wire n_2977;
 wire n_2978;
 wire n_2979;
 wire n_298;
 wire n_2980;
 wire n_2981;
 wire n_2982;
 wire n_2983;
 wire n_2984;
 wire n_2985;
 wire n_2986;
 wire n_2987;
 wire n_2988;
 wire n_2989;
 wire n_299;
 wire n_2990;
 wire n_2991;
 wire n_2992;
 wire n_2993;
 wire n_2994;
 wire n_2995;
 wire n_2996;
 wire n_2997;
 wire n_2998;
 wire n_2999;
 wire n_3;
 wire n_30;
 wire n_300;
 wire n_3000;
 wire n_3001;
 wire n_3002;
 wire n_3003;
 wire n_3004;
 wire n_3005;
 wire n_3006;
 wire n_3007;
 wire n_3008;
 wire n_3009;
 wire n_301;
 wire n_3010;
 wire n_3011;
 wire n_3012;
 wire n_3013;
 wire n_3014;
 wire n_3015;
 wire n_3016;
 wire n_3017;
 wire n_3018;
 wire n_3019;
 wire n_302;
 wire n_3020;
 wire n_3021;
 wire n_3022;
 wire n_3023;
 wire n_3024;
 wire n_3025;
 wire n_3026;
 wire n_3027;
 wire n_3028;
 wire n_3029;
 wire n_303;
 wire n_3030;
 wire n_3031;
 wire n_3032;
 wire n_3033;
 wire n_3034;
 wire n_3035;
 wire n_3036;
 wire n_3037;
 wire n_3038;
 wire n_3039;
 wire n_304;
 wire n_3040;
 wire n_3041;
 wire n_3042;
 wire n_3043;
 wire n_3044;
 wire n_3045;
 wire n_3046;
 wire n_3047;
 wire n_3048;
 wire n_3049;
 wire n_305;
 wire n_3050;
 wire n_3051;
 wire n_3052;
 wire n_3053;
 wire n_3054;
 wire n_3055;
 wire n_3056;
 wire n_3057;
 wire n_3058;
 wire n_3059;
 wire n_306;
 wire n_3060;
 wire n_3061;
 wire n_3062;
 wire n_3063;
 wire n_3064;
 wire n_3065;
 wire n_3066;
 wire n_3067;
 wire n_3068;
 wire n_3069;
 wire n_3070;
 wire n_3071;
 wire n_3072;
 wire n_3073;
 wire n_3074;
 wire n_3075;
 wire n_3076;
 wire n_3077;
 wire n_3078;
 wire n_3079;
 wire n_3080;
 wire n_3081;
 wire n_3082;
 wire n_3083;
 wire n_3084;
 wire n_3085;
 wire n_3086;
 wire n_3087;
 wire n_3088;
 wire n_3089;
 wire n_309;
 wire n_3090;
 wire n_3091;
 wire n_3092;
 wire n_3093;
 wire n_3094;
 wire n_3095;
 wire n_3096;
 wire n_3097;
 wire n_3098;
 wire n_3099;
 wire n_31;
 wire n_310;
 wire n_3100;
 wire n_3101;
 wire n_3102;
 wire n_3103;
 wire n_3104;
 wire n_3105;
 wire n_3106;
 wire n_3107;
 wire n_3108;
 wire n_3109;
 wire n_311;
 wire n_3110;
 wire n_3111;
 wire n_3112;
 wire n_3113;
 wire n_3114;
 wire n_3115;
 wire n_3116;
 wire n_3117;
 wire n_3118;
 wire n_3119;
 wire n_312;
 wire n_3120;
 wire n_3121;
 wire n_3122;
 wire n_3123;
 wire n_3124;
 wire n_3125;
 wire n_3126;
 wire n_3127;
 wire n_3128;
 wire n_3129;
 wire n_313;
 wire n_3130;
 wire n_3131;
 wire n_3132;
 wire n_3133;
 wire n_3134;
 wire n_3135;
 wire n_3136;
 wire n_3137;
 wire n_3138;
 wire n_3139;
 wire n_314;
 wire n_3140;
 wire n_3141;
 wire n_3142;
 wire n_3143;
 wire n_3144;
 wire n_3145;
 wire n_3146;
 wire n_3147;
 wire n_3148;
 wire n_3149;
 wire n_3150;
 wire n_3151;
 wire n_3152;
 wire n_3153;
 wire n_3154;
 wire n_3155;
 wire n_3156;
 wire n_3157;
 wire n_3158;
 wire n_3159;
 wire n_316;
 wire n_3160;
 wire n_3161;
 wire n_3162;
 wire n_3163;
 wire n_3164;
 wire n_3165;
 wire n_3166;
 wire n_3167;
 wire n_3168;
 wire n_3169;
 wire n_3170;
 wire n_3171;
 wire n_3172;
 wire n_3173;
 wire n_3174;
 wire n_3175;
 wire n_3176;
 wire n_3177;
 wire n_3178;
 wire n_3179;
 wire n_3180;
 wire n_3181;
 wire n_3182;
 wire n_3183;
 wire n_3184;
 wire n_3185;
 wire n_3186;
 wire n_3187;
 wire n_3188;
 wire n_3189;
 wire n_319;
 wire n_3190;
 wire n_3191;
 wire n_3192;
 wire n_3193;
 wire n_3194;
 wire n_3195;
 wire n_3196;
 wire n_3197;
 wire n_3198;
 wire n_3199;
 wire n_32;
 wire n_320;
 wire n_3200;
 wire n_3201;
 wire n_3202;
 wire n_3203;
 wire n_3204;
 wire n_3205;
 wire n_3206;
 wire n_3207;
 wire n_3208;
 wire n_3209;
 wire n_321;
 wire n_3210;
 wire n_3211;
 wire n_3212;
 wire n_3213;
 wire n_3214;
 wire n_3215;
 wire n_3216;
 wire n_3217;
 wire n_3218;
 wire n_3219;
 wire n_322;
 wire n_3220;
 wire n_3221;
 wire n_3222;
 wire n_3223;
 wire n_3224;
 wire n_3225;
 wire n_3226;
 wire n_3227;
 wire n_3228;
 wire n_3229;
 wire n_3230;
 wire n_3231;
 wire n_3232;
 wire n_3233;
 wire n_3234;
 wire n_3235;
 wire n_3236;
 wire n_3237;
 wire n_3238;
 wire n_3239;
 wire n_324;
 wire n_3240;
 wire n_3241;
 wire n_3242;
 wire n_3243;
 wire n_3244;
 wire n_3245;
 wire n_3246;
 wire n_3247;
 wire n_3248;
 wire n_3249;
 wire n_325;
 wire n_3250;
 wire n_3251;
 wire n_3252;
 wire n_3253;
 wire n_3254;
 wire n_3255;
 wire n_3256;
 wire n_3257;
 wire n_3258;
 wire n_3259;
 wire n_326;
 wire n_3260;
 wire n_3261;
 wire n_3262;
 wire n_3263;
 wire n_3265;
 wire n_3266;
 wire n_3267;
 wire n_3268;
 wire n_3269;
 wire n_3270;
 wire n_3271;
 wire n_3272;
 wire n_3273;
 wire n_3274;
 wire n_3275;
 wire n_3276;
 wire n_3277;
 wire n_3278;
 wire n_3279;
 wire n_328;
 wire n_3280;
 wire n_3281;
 wire n_3282;
 wire n_3283;
 wire n_3284;
 wire n_3285;
 wire n_3286;
 wire n_3287;
 wire n_3288;
 wire n_3289;
 wire n_3290;
 wire n_3291;
 wire n_3292;
 wire n_3293;
 wire n_3294;
 wire n_3295;
 wire n_3296;
 wire n_3297;
 wire n_3298;
 wire n_3299;
 wire n_33;
 wire n_330;
 wire n_3300;
 wire n_3301;
 wire n_3302;
 wire n_3303;
 wire n_3304;
 wire n_3305;
 wire n_3306;
 wire n_3307;
 wire n_3308;
 wire n_3309;
 wire n_331;
 wire n_3310;
 wire n_3311;
 wire n_3312;
 wire n_3313;
 wire n_3314;
 wire n_3315;
 wire n_3316;
 wire n_3317;
 wire n_3319;
 wire n_332;
 wire n_3320;
 wire n_3321;
 wire n_3322;
 wire n_3323;
 wire n_3324;
 wire n_3325;
 wire n_3326;
 wire n_3327;
 wire n_3328;
 wire n_3329;
 wire n_3330;
 wire n_3331;
 wire n_3332;
 wire n_3333;
 wire n_3334;
 wire n_3335;
 wire n_3336;
 wire n_3337;
 wire n_3338;
 wire n_334;
 wire n_3340;
 wire n_3341;
 wire n_3342;
 wire n_3343;
 wire n_3344;
 wire n_3345;
 wire n_3346;
 wire n_3347;
 wire n_3348;
 wire n_3349;
 wire n_335;
 wire n_3350;
 wire n_3351;
 wire n_3352;
 wire n_3353;
 wire n_3354;
 wire n_3355;
 wire n_3356;
 wire n_3357;
 wire n_3358;
 wire n_3359;
 wire n_336;
 wire n_3360;
 wire n_3361;
 wire n_3363;
 wire n_3364;
 wire n_3365;
 wire n_3366;
 wire n_3367;
 wire n_3368;
 wire n_3369;
 wire n_337;
 wire n_3370;
 wire n_3371;
 wire n_3372;
 wire n_3373;
 wire n_3374;
 wire n_3375;
 wire n_3376;
 wire n_3377;
 wire n_3378;
 wire n_3379;
 wire n_338;
 wire n_3380;
 wire n_3381;
 wire n_3382;
 wire n_3383;
 wire n_3384;
 wire n_3385;
 wire n_3386;
 wire n_3387;
 wire n_3388;
 wire n_3389;
 wire n_3390;
 wire n_3391;
 wire n_3392;
 wire n_3393;
 wire n_3394;
 wire n_3395;
 wire n_3396;
 wire n_3398;
 wire n_3399;
 wire n_34;
 wire n_340;
 wire n_3400;
 wire n_3401;
 wire n_3402;
 wire n_3403;
 wire n_3404;
 wire n_3405;
 wire n_3406;
 wire n_3407;
 wire n_3408;
 wire n_3409;
 wire n_341;
 wire n_3410;
 wire n_3411;
 wire n_3412;
 wire n_3413;
 wire n_3414;
 wire n_3415;
 wire n_3416;
 wire n_3417;
 wire n_3418;
 wire n_3419;
 wire n_342;
 wire n_3420;
 wire n_3421;
 wire n_3422;
 wire n_3423;
 wire n_3424;
 wire n_3425;
 wire n_3427;
 wire n_3428;
 wire n_3429;
 wire n_3430;
 wire n_3431;
 wire n_3432;
 wire n_3433;
 wire n_3434;
 wire n_3435;
 wire n_3436;
 wire n_3437;
 wire n_3438;
 wire n_3439;
 wire n_344;
 wire n_3440;
 wire n_3441;
 wire n_3442;
 wire n_3443;
 wire n_3444;
 wire n_3445;
 wire n_3446;
 wire n_3447;
 wire n_3448;
 wire n_3449;
 wire n_345;
 wire n_3450;
 wire n_3451;
 wire n_3452;
 wire n_3453;
 wire n_3454;
 wire n_3455;
 wire n_3456;
 wire n_3457;
 wire n_3458;
 wire n_3459;
 wire n_346;
 wire n_3460;
 wire n_3461;
 wire n_3462;
 wire n_3463;
 wire n_3464;
 wire n_3465;
 wire n_3466;
 wire n_3467;
 wire n_3468;
 wire n_3469;
 wire n_347;
 wire n_3470;
 wire n_3471;
 wire n_3472;
 wire n_3473;
 wire n_3474;
 wire n_3475;
 wire n_3476;
 wire n_3477;
 wire n_3478;
 wire n_3479;
 wire n_348;
 wire n_3480;
 wire n_3481;
 wire n_3482;
 wire n_3483;
 wire n_3484;
 wire n_3485;
 wire n_3486;
 wire n_3487;
 wire n_3488;
 wire n_3489;
 wire n_349;
 wire n_3490;
 wire n_3491;
 wire n_3492;
 wire n_3493;
 wire n_3494;
 wire n_3495;
 wire n_3496;
 wire n_3497;
 wire n_3498;
 wire n_3499;
 wire n_35;
 wire n_350;
 wire n_3500;
 wire n_3501;
 wire n_3502;
 wire n_3503;
 wire n_3504;
 wire n_3505;
 wire n_3506;
 wire n_3507;
 wire n_3508;
 wire n_3509;
 wire n_351;
 wire n_3510;
 wire n_3511;
 wire n_3512;
 wire n_3513;
 wire n_3514;
 wire n_3515;
 wire n_3516;
 wire n_3517;
 wire n_3518;
 wire n_3519;
 wire n_3520;
 wire n_3521;
 wire n_3522;
 wire n_3523;
 wire n_3524;
 wire n_3525;
 wire n_3526;
 wire n_3527;
 wire n_3528;
 wire n_3529;
 wire n_353;
 wire n_3530;
 wire n_3531;
 wire n_3532;
 wire n_3533;
 wire n_3534;
 wire n_3535;
 wire n_3536;
 wire n_3537;
 wire n_3538;
 wire n_3539;
 wire n_3540;
 wire n_3541;
 wire n_3542;
 wire n_3543;
 wire n_3544;
 wire n_3545;
 wire n_3546;
 wire n_3547;
 wire n_3548;
 wire n_3549;
 wire n_355;
 wire n_3550;
 wire n_3551;
 wire n_3552;
 wire n_3553;
 wire n_3554;
 wire n_3555;
 wire n_3556;
 wire n_3557;
 wire n_3558;
 wire n_3559;
 wire n_356;
 wire n_3560;
 wire n_3561;
 wire n_3562;
 wire n_3563;
 wire n_3564;
 wire n_3565;
 wire n_3566;
 wire n_3567;
 wire n_3568;
 wire n_3569;
 wire n_357;
 wire n_3570;
 wire n_3571;
 wire n_3572;
 wire n_3573;
 wire n_3574;
 wire n_3575;
 wire n_3576;
 wire n_3577;
 wire n_3578;
 wire n_3579;
 wire n_3580;
 wire n_3581;
 wire n_3582;
 wire n_3583;
 wire n_3584;
 wire n_3585;
 wire n_3586;
 wire n_3587;
 wire n_3588;
 wire n_3589;
 wire n_3590;
 wire n_3591;
 wire n_3592;
 wire n_3593;
 wire n_3594;
 wire n_3595;
 wire n_3596;
 wire n_3597;
 wire n_3598;
 wire n_3599;
 wire n_36;
 wire n_360;
 wire n_3600;
 wire n_3601;
 wire n_3602;
 wire n_3603;
 wire n_3604;
 wire n_3605;
 wire n_3606;
 wire n_3607;
 wire n_3608;
 wire n_3609;
 wire n_361;
 wire n_3610;
 wire n_3611;
 wire n_3612;
 wire n_3613;
 wire n_3614;
 wire n_3615;
 wire n_3616;
 wire n_3617;
 wire n_3618;
 wire n_3619;
 wire n_362;
 wire n_3620;
 wire n_3621;
 wire n_3622;
 wire n_3623;
 wire n_3624;
 wire n_3625;
 wire n_3626;
 wire n_3627;
 wire n_3628;
 wire n_3629;
 wire n_363;
 wire n_3630;
 wire n_3631;
 wire n_3632;
 wire n_3633;
 wire n_3634;
 wire n_3635;
 wire n_3636;
 wire n_3637;
 wire n_3638;
 wire n_3639;
 wire n_364;
 wire n_3640;
 wire n_3641;
 wire n_3642;
 wire n_3643;
 wire n_3644;
 wire n_3645;
 wire n_3646;
 wire n_3647;
 wire n_3648;
 wire n_3649;
 wire n_365;
 wire n_3650;
 wire n_3651;
 wire n_3652;
 wire n_3653;
 wire n_3654;
 wire n_3655;
 wire n_3657;
 wire n_3658;
 wire n_3659;
 wire n_3660;
 wire n_3661;
 wire n_3662;
 wire n_3663;
 wire n_3664;
 wire n_3665;
 wire n_3666;
 wire n_3667;
 wire n_3668;
 wire n_3669;
 wire n_367;
 wire n_3670;
 wire n_3671;
 wire n_3672;
 wire n_3673;
 wire n_3674;
 wire n_3675;
 wire n_3676;
 wire n_3677;
 wire n_3678;
 wire n_3679;
 wire n_368;
 wire n_3680;
 wire n_3681;
 wire n_3682;
 wire n_3683;
 wire n_3684;
 wire n_3685;
 wire n_3686;
 wire n_3687;
 wire n_3688;
 wire n_3689;
 wire n_369;
 wire n_3690;
 wire n_3691;
 wire n_3692;
 wire n_3693;
 wire n_3694;
 wire n_3695;
 wire n_3696;
 wire n_3697;
 wire n_3698;
 wire n_3699;
 wire n_37;
 wire n_370;
 wire n_3700;
 wire n_3701;
 wire n_3702;
 wire n_3703;
 wire n_3704;
 wire n_3705;
 wire n_3706;
 wire n_3707;
 wire n_3708;
 wire n_3709;
 wire n_371;
 wire n_3710;
 wire n_3711;
 wire n_3712;
 wire n_3713;
 wire n_3714;
 wire n_3715;
 wire n_3716;
 wire n_3717;
 wire n_3718;
 wire n_3719;
 wire n_3720;
 wire n_3721;
 wire n_3722;
 wire n_3723;
 wire n_3724;
 wire n_3725;
 wire n_3726;
 wire n_3727;
 wire n_3728;
 wire n_3729;
 wire n_373;
 wire n_3730;
 wire n_3731;
 wire n_3732;
 wire n_3733;
 wire n_3734;
 wire n_3735;
 wire n_3736;
 wire n_3737;
 wire n_3738;
 wire n_3739;
 wire n_3740;
 wire n_3741;
 wire n_3742;
 wire n_3743;
 wire n_3744;
 wire n_3745;
 wire n_3746;
 wire n_3747;
 wire n_3748;
 wire n_3749;
 wire n_375;
 wire n_3750;
 wire n_3751;
 wire n_3752;
 wire n_3753;
 wire n_3754;
 wire n_3755;
 wire n_3756;
 wire n_3757;
 wire n_3758;
 wire n_3759;
 wire n_376;
 wire n_3760;
 wire n_3761;
 wire n_3762;
 wire n_3763;
 wire n_3764;
 wire n_3765;
 wire n_3766;
 wire n_3767;
 wire n_3768;
 wire n_3769;
 wire n_377;
 wire n_3770;
 wire n_3771;
 wire n_3772;
 wire n_3773;
 wire n_3774;
 wire n_3775;
 wire n_3776;
 wire n_3777;
 wire n_3778;
 wire n_3779;
 wire n_378;
 wire n_3780;
 wire n_3781;
 wire n_3782;
 wire n_3783;
 wire n_3784;
 wire n_3785;
 wire n_3786;
 wire n_3787;
 wire n_3788;
 wire n_3789;
 wire n_379;
 wire n_3790;
 wire n_3791;
 wire n_3792;
 wire n_3793;
 wire n_3794;
 wire n_3795;
 wire n_3796;
 wire n_3797;
 wire n_3798;
 wire n_3799;
 wire n_380;
 wire n_3800;
 wire n_3801;
 wire n_3802;
 wire n_3803;
 wire n_3804;
 wire n_3805;
 wire n_3806;
 wire n_3807;
 wire n_3808;
 wire n_3809;
 wire n_381;
 wire n_3810;
 wire n_3811;
 wire n_3812;
 wire n_3813;
 wire n_3814;
 wire n_3815;
 wire n_3816;
 wire n_3817;
 wire n_3818;
 wire n_3819;
 wire n_3820;
 wire n_3821;
 wire n_3822;
 wire n_3823;
 wire n_3824;
 wire n_3825;
 wire n_3826;
 wire n_3827;
 wire n_3828;
 wire n_3829;
 wire n_383;
 wire n_3830;
 wire n_3831;
 wire n_3832;
 wire n_3833;
 wire n_3834;
 wire n_3835;
 wire n_3836;
 wire n_3837;
 wire n_3838;
 wire n_3839;
 wire n_384;
 wire n_3840;
 wire n_3841;
 wire n_3842;
 wire n_3843;
 wire n_3844;
 wire n_3845;
 wire n_3846;
 wire n_3847;
 wire n_3848;
 wire n_3849;
 wire n_385;
 wire n_3850;
 wire n_3851;
 wire n_3852;
 wire n_3853;
 wire n_3854;
 wire n_3855;
 wire n_3856;
 wire n_3857;
 wire n_3858;
 wire n_3859;
 wire n_386;
 wire n_3860;
 wire n_3861;
 wire n_3862;
 wire n_3863;
 wire n_3864;
 wire n_3865;
 wire n_3866;
 wire n_3867;
 wire n_3868;
 wire n_3869;
 wire n_387;
 wire n_3870;
 wire n_3871;
 wire n_3872;
 wire n_3873;
 wire n_3874;
 wire n_3875;
 wire n_3876;
 wire n_3877;
 wire n_3878;
 wire n_3879;
 wire n_388;
 wire n_3880;
 wire n_3881;
 wire n_3882;
 wire n_3883;
 wire n_3884;
 wire n_3885;
 wire n_3886;
 wire n_3887;
 wire n_3888;
 wire n_3889;
 wire n_389;
 wire n_3890;
 wire n_3891;
 wire n_3892;
 wire n_3893;
 wire n_3894;
 wire n_3895;
 wire n_3896;
 wire n_3897;
 wire n_3898;
 wire n_3899;
 wire n_39;
 wire n_390;
 wire n_3900;
 wire n_3901;
 wire n_3902;
 wire n_3903;
 wire n_3904;
 wire n_3905;
 wire n_3906;
 wire n_3907;
 wire n_3908;
 wire n_3909;
 wire n_391;
 wire n_3910;
 wire n_3911;
 wire n_3912;
 wire n_3913;
 wire n_3914;
 wire n_3915;
 wire n_3916;
 wire n_3917;
 wire n_3918;
 wire n_3919;
 wire n_392;
 wire n_3920;
 wire n_3921;
 wire n_3922;
 wire n_3923;
 wire n_3924;
 wire n_3925;
 wire n_3926;
 wire n_3927;
 wire n_3928;
 wire n_3929;
 wire n_393;
 wire n_3930;
 wire n_3931;
 wire n_3932;
 wire n_3933;
 wire n_3934;
 wire n_3935;
 wire n_3936;
 wire n_3937;
 wire n_3938;
 wire n_3939;
 wire n_394;
 wire n_3940;
 wire n_3941;
 wire n_3942;
 wire n_3943;
 wire n_3944;
 wire n_3945;
 wire n_3946;
 wire n_3947;
 wire n_3948;
 wire n_3949;
 wire n_395;
 wire n_3950;
 wire n_3951;
 wire n_3952;
 wire n_3953;
 wire n_3954;
 wire n_3955;
 wire n_3956;
 wire n_3957;
 wire n_3958;
 wire n_3959;
 wire n_396;
 wire n_3960;
 wire n_3961;
 wire n_3962;
 wire n_3963;
 wire n_3964;
 wire n_3965;
 wire n_3966;
 wire n_3967;
 wire n_3968;
 wire n_3969;
 wire n_397;
 wire n_3970;
 wire n_3971;
 wire n_3972;
 wire n_3973;
 wire n_3974;
 wire n_3975;
 wire n_3976;
 wire n_3977;
 wire n_3978;
 wire n_3979;
 wire n_398;
 wire n_3980;
 wire n_3981;
 wire n_3982;
 wire n_3983;
 wire n_3984;
 wire n_3985;
 wire n_3986;
 wire n_3987;
 wire n_3988;
 wire n_3989;
 wire n_399;
 wire n_3990;
 wire n_3991;
 wire n_3992;
 wire n_3993;
 wire n_3994;
 wire n_3995;
 wire n_3996;
 wire n_3997;
 wire n_3998;
 wire n_3999;
 wire n_4;
 wire n_40;
 wire n_400;
 wire n_4000;
 wire n_4001;
 wire n_4002;
 wire n_4003;
 wire n_4004;
 wire n_4005;
 wire n_4006;
 wire n_4007;
 wire n_4008;
 wire n_4009;
 wire n_401;
 wire n_4010;
 wire n_4011;
 wire n_4012;
 wire n_4013;
 wire n_4014;
 wire n_4015;
 wire n_4016;
 wire n_4017;
 wire n_4018;
 wire n_4019;
 wire n_402;
 wire n_4020;
 wire n_4021;
 wire n_4022;
 wire n_4023;
 wire n_4024;
 wire n_4025;
 wire n_4026;
 wire n_4027;
 wire n_4028;
 wire n_4029;
 wire n_403;
 wire n_4030;
 wire n_4031;
 wire n_4032;
 wire n_4033;
 wire n_4034;
 wire n_4035;
 wire n_4036;
 wire n_4037;
 wire n_4038;
 wire n_4039;
 wire n_404;
 wire n_4040;
 wire n_4041;
 wire n_4042;
 wire n_4043;
 wire n_4044;
 wire n_4045;
 wire n_4046;
 wire n_4047;
 wire n_4048;
 wire n_4049;
 wire n_405;
 wire n_4050;
 wire n_4051;
 wire n_4052;
 wire n_4053;
 wire n_4054;
 wire n_4055;
 wire n_4056;
 wire n_4057;
 wire n_4058;
 wire n_4059;
 wire n_406;
 wire n_4060;
 wire n_4061;
 wire n_4062;
 wire n_4063;
 wire n_4064;
 wire n_4065;
 wire n_4066;
 wire n_4067;
 wire n_4068;
 wire n_4069;
 wire n_407;
 wire n_4070;
 wire n_4071;
 wire n_4072;
 wire n_4073;
 wire n_4074;
 wire n_4075;
 wire n_4076;
 wire n_4077;
 wire n_4078;
 wire n_4079;
 wire n_408;
 wire n_4080;
 wire n_4081;
 wire n_4082;
 wire n_4083;
 wire n_4084;
 wire n_4085;
 wire n_4086;
 wire n_4087;
 wire n_4088;
 wire n_4089;
 wire n_409;
 wire n_4090;
 wire n_4091;
 wire n_4092;
 wire n_4093;
 wire n_4094;
 wire n_4095;
 wire n_4096;
 wire n_4097;
 wire n_4098;
 wire n_4099;
 wire n_41;
 wire n_410;
 wire n_4100;
 wire n_4101;
 wire n_4102;
 wire n_4103;
 wire n_4104;
 wire n_4105;
 wire n_4106;
 wire n_4107;
 wire n_4108;
 wire n_4109;
 wire n_411;
 wire n_4110;
 wire n_4111;
 wire n_4112;
 wire n_4113;
 wire n_4114;
 wire n_4115;
 wire n_4116;
 wire n_4117;
 wire n_4118;
 wire n_4119;
 wire n_412;
 wire n_4120;
 wire n_4121;
 wire n_4122;
 wire n_4123;
 wire n_4124;
 wire n_4125;
 wire n_4126;
 wire n_4127;
 wire n_4128;
 wire n_4129;
 wire n_413;
 wire n_4130;
 wire n_4131;
 wire n_4132;
 wire n_4133;
 wire n_4134;
 wire n_4135;
 wire n_4136;
 wire n_4137;
 wire n_4138;
 wire n_4139;
 wire n_414;
 wire n_4140;
 wire n_4141;
 wire n_4142;
 wire n_4143;
 wire n_4144;
 wire n_4145;
 wire n_4146;
 wire n_4147;
 wire n_4148;
 wire n_4149;
 wire n_415;
 wire n_4150;
 wire n_4151;
 wire n_4152;
 wire n_4153;
 wire n_4154;
 wire n_4155;
 wire n_4156;
 wire n_4157;
 wire n_4158;
 wire n_4159;
 wire n_416;
 wire n_4160;
 wire n_4161;
 wire n_4162;
 wire n_4163;
 wire n_4164;
 wire n_4165;
 wire n_4166;
 wire n_4167;
 wire n_4168;
 wire n_4169;
 wire n_417;
 wire n_4170;
 wire n_4171;
 wire n_4172;
 wire n_4173;
 wire n_4174;
 wire n_4175;
 wire n_4176;
 wire n_4177;
 wire n_4178;
 wire n_4179;
 wire n_418;
 wire n_4180;
 wire n_4181;
 wire n_4182;
 wire n_4183;
 wire n_4184;
 wire n_4185;
 wire n_4186;
 wire n_4187;
 wire n_4188;
 wire n_4189;
 wire n_419;
 wire n_4190;
 wire n_4191;
 wire n_4192;
 wire n_4193;
 wire n_4194;
 wire n_4195;
 wire n_4196;
 wire n_4197;
 wire n_4198;
 wire n_4199;
 wire n_42;
 wire n_420;
 wire n_4200;
 wire n_4201;
 wire n_4202;
 wire n_4203;
 wire n_4204;
 wire n_4205;
 wire n_4206;
 wire n_4207;
 wire n_4208;
 wire n_4209;
 wire n_421;
 wire n_4210;
 wire n_4211;
 wire n_4212;
 wire n_4213;
 wire n_4214;
 wire n_4215;
 wire n_4216;
 wire n_4217;
 wire n_4218;
 wire n_4219;
 wire n_422;
 wire n_4220;
 wire n_4221;
 wire n_4222;
 wire n_4223;
 wire n_4224;
 wire n_4225;
 wire n_4226;
 wire n_4227;
 wire n_4228;
 wire n_4229;
 wire n_423;
 wire n_4230;
 wire n_4231;
 wire n_4232;
 wire n_4233;
 wire n_4234;
 wire n_4235;
 wire n_4236;
 wire n_4237;
 wire n_4238;
 wire n_4239;
 wire n_424;
 wire n_4240;
 wire n_4241;
 wire n_4242;
 wire n_4243;
 wire n_4244;
 wire n_4245;
 wire n_4246;
 wire n_4247;
 wire n_4248;
 wire n_4249;
 wire n_425;
 wire n_4250;
 wire n_4251;
 wire n_4252;
 wire n_4253;
 wire n_4254;
 wire n_4255;
 wire n_4256;
 wire n_4257;
 wire n_4258;
 wire n_4259;
 wire n_426;
 wire n_4260;
 wire n_4261;
 wire n_4262;
 wire n_4263;
 wire n_4264;
 wire n_4265;
 wire n_4266;
 wire n_4267;
 wire n_4268;
 wire n_4269;
 wire n_427;
 wire n_4270;
 wire n_4271;
 wire n_4272;
 wire n_4273;
 wire n_4274;
 wire n_4275;
 wire n_4276;
 wire n_4277;
 wire n_4278;
 wire n_4279;
 wire n_428;
 wire n_4280;
 wire n_4281;
 wire n_4282;
 wire n_4283;
 wire n_4284;
 wire n_4285;
 wire n_4286;
 wire n_4287;
 wire n_4288;
 wire n_4289;
 wire n_429;
 wire n_4290;
 wire n_4291;
 wire n_4292;
 wire n_4293;
 wire n_4294;
 wire n_4295;
 wire n_4296;
 wire n_4297;
 wire n_4298;
 wire n_4299;
 wire n_43;
 wire n_430;
 wire n_4300;
 wire n_4301;
 wire n_4302;
 wire n_4303;
 wire n_4304;
 wire n_4305;
 wire n_4306;
 wire n_4307;
 wire n_4308;
 wire n_4309;
 wire n_431;
 wire n_4310;
 wire n_4311;
 wire n_4312;
 wire n_4313;
 wire n_4314;
 wire n_4315;
 wire n_4316;
 wire n_4317;
 wire n_4318;
 wire n_4319;
 wire n_432;
 wire n_4320;
 wire n_4321;
 wire n_4322;
 wire n_4323;
 wire n_4324;
 wire n_4325;
 wire n_4326;
 wire n_4327;
 wire n_4328;
 wire n_4329;
 wire n_433;
 wire n_4330;
 wire n_4331;
 wire n_4332;
 wire n_4333;
 wire n_4334;
 wire n_4335;
 wire n_4336;
 wire n_4337;
 wire n_4338;
 wire n_4339;
 wire n_434;
 wire n_4340;
 wire n_4341;
 wire n_4342;
 wire n_4343;
 wire n_4344;
 wire n_4345;
 wire n_4346;
 wire n_4347;
 wire n_4348;
 wire n_4349;
 wire n_435;
 wire n_4350;
 wire n_4351;
 wire n_4352;
 wire n_4353;
 wire n_4354;
 wire n_4355;
 wire n_4356;
 wire n_4357;
 wire n_4358;
 wire n_4359;
 wire n_436;
 wire n_4360;
 wire n_4361;
 wire n_4362;
 wire n_4363;
 wire n_4364;
 wire n_4365;
 wire n_4366;
 wire n_4367;
 wire n_4368;
 wire n_4369;
 wire n_437;
 wire n_4370;
 wire n_4371;
 wire n_4372;
 wire n_4373;
 wire n_4374;
 wire n_4375;
 wire n_4376;
 wire n_4377;
 wire n_4378;
 wire n_4379;
 wire n_438;
 wire n_4380;
 wire n_4381;
 wire n_4382;
 wire n_4383;
 wire n_4384;
 wire n_4385;
 wire n_4386;
 wire n_4387;
 wire n_4388;
 wire n_4389;
 wire n_439;
 wire n_4390;
 wire n_4391;
 wire n_4392;
 wire n_4393;
 wire n_4394;
 wire n_4395;
 wire n_4396;
 wire n_4397;
 wire n_4398;
 wire n_4399;
 wire n_44;
 wire n_440;
 wire n_4400;
 wire n_4401;
 wire n_4402;
 wire n_4403;
 wire n_4404;
 wire n_4405;
 wire n_4406;
 wire n_4407;
 wire n_4408;
 wire n_4409;
 wire n_441;
 wire n_4410;
 wire n_4411;
 wire n_4412;
 wire n_4413;
 wire n_4414;
 wire n_4415;
 wire n_4416;
 wire n_4417;
 wire n_4418;
 wire n_4419;
 wire n_442;
 wire n_4420;
 wire n_4421;
 wire n_4422;
 wire n_4423;
 wire n_4424;
 wire n_4425;
 wire n_4427;
 wire n_4428;
 wire n_4429;
 wire n_443;
 wire n_4430;
 wire n_4431;
 wire n_4432;
 wire n_4433;
 wire n_4434;
 wire n_4435;
 wire n_4436;
 wire n_4437;
 wire n_4438;
 wire n_4439;
 wire n_444;
 wire n_4440;
 wire n_4441;
 wire n_4442;
 wire n_4443;
 wire n_4444;
 wire n_4445;
 wire n_4446;
 wire n_4447;
 wire n_4448;
 wire n_4449;
 wire n_445;
 wire n_4450;
 wire n_4451;
 wire n_4452;
 wire n_4453;
 wire n_4454;
 wire n_4455;
 wire n_4456;
 wire n_4457;
 wire n_4458;
 wire n_4459;
 wire n_446;
 wire n_4460;
 wire n_4461;
 wire n_4462;
 wire n_4463;
 wire n_4464;
 wire n_4465;
 wire n_4466;
 wire n_4467;
 wire n_4468;
 wire n_4469;
 wire n_447;
 wire n_4470;
 wire n_4471;
 wire n_4473;
 wire n_4474;
 wire n_4475;
 wire n_4476;
 wire n_4477;
 wire n_4478;
 wire n_4479;
 wire n_448;
 wire n_4480;
 wire n_4481;
 wire n_4482;
 wire n_4483;
 wire n_4484;
 wire n_4485;
 wire n_4486;
 wire n_4487;
 wire n_4488;
 wire n_4489;
 wire n_449;
 wire n_4490;
 wire n_4491;
 wire n_4492;
 wire n_4493;
 wire n_4494;
 wire n_4495;
 wire n_4496;
 wire n_4497;
 wire n_4498;
 wire n_4499;
 wire n_45;
 wire n_450;
 wire n_4500;
 wire n_4501;
 wire n_4502;
 wire n_4503;
 wire n_4504;
 wire n_4505;
 wire n_4506;
 wire n_4507;
 wire n_4508;
 wire n_4509;
 wire n_451;
 wire n_4510;
 wire n_4511;
 wire n_4512;
 wire n_4513;
 wire n_4514;
 wire n_4515;
 wire n_4516;
 wire n_4517;
 wire n_4518;
 wire n_4519;
 wire n_452;
 wire n_4520;
 wire n_4521;
 wire n_4522;
 wire n_4523;
 wire n_4524;
 wire n_4525;
 wire n_4526;
 wire n_4527;
 wire n_4528;
 wire n_4529;
 wire n_453;
 wire n_4530;
 wire n_4531;
 wire n_4532;
 wire n_4533;
 wire n_4534;
 wire n_4535;
 wire n_4536;
 wire n_4537;
 wire n_4538;
 wire n_4539;
 wire n_454;
 wire n_4540;
 wire n_4541;
 wire n_4542;
 wire n_4543;
 wire n_4544;
 wire n_4545;
 wire n_4546;
 wire n_4547;
 wire n_4548;
 wire n_4549;
 wire n_455;
 wire n_4550;
 wire n_4551;
 wire n_4552;
 wire n_4553;
 wire n_4554;
 wire n_4555;
 wire n_4556;
 wire n_4557;
 wire n_4558;
 wire n_4559;
 wire n_456;
 wire n_4560;
 wire n_4561;
 wire n_4562;
 wire n_4563;
 wire n_4564;
 wire n_4565;
 wire n_4566;
 wire n_4567;
 wire n_4568;
 wire n_4569;
 wire n_457;
 wire n_4570;
 wire n_4571;
 wire n_4572;
 wire n_4573;
 wire n_4574;
 wire n_4575;
 wire n_4576;
 wire n_4577;
 wire n_4578;
 wire n_4579;
 wire n_458;
 wire n_4580;
 wire n_4581;
 wire n_4582;
 wire n_4583;
 wire n_4584;
 wire n_4585;
 wire n_4586;
 wire n_4587;
 wire n_4588;
 wire n_4589;
 wire n_459;
 wire n_4590;
 wire n_4591;
 wire n_4592;
 wire n_4593;
 wire n_4594;
 wire n_4595;
 wire n_4596;
 wire n_4597;
 wire n_4598;
 wire n_4599;
 wire n_46;
 wire n_460;
 wire n_4600;
 wire n_4601;
 wire n_4602;
 wire n_4603;
 wire n_4604;
 wire n_4605;
 wire n_4606;
 wire n_4607;
 wire n_4608;
 wire n_4609;
 wire n_461;
 wire n_4610;
 wire n_4611;
 wire n_4612;
 wire n_4613;
 wire n_4614;
 wire n_4615;
 wire n_4616;
 wire n_4617;
 wire n_4618;
 wire n_4619;
 wire n_462;
 wire n_4620;
 wire n_4621;
 wire n_4622;
 wire n_4623;
 wire n_4624;
 wire n_4625;
 wire n_4626;
 wire n_4627;
 wire n_4628;
 wire n_4629;
 wire n_463;
 wire n_4630;
 wire n_4631;
 wire n_4632;
 wire n_4633;
 wire n_4634;
 wire n_4635;
 wire n_4636;
 wire n_4637;
 wire n_4638;
 wire n_4639;
 wire n_464;
 wire n_4640;
 wire n_4641;
 wire n_4642;
 wire n_4643;
 wire n_4644;
 wire n_4645;
 wire n_4646;
 wire n_4647;
 wire n_4648;
 wire n_4649;
 wire n_465;
 wire n_4650;
 wire n_4651;
 wire n_4652;
 wire n_4653;
 wire n_4654;
 wire n_4655;
 wire n_4656;
 wire n_4657;
 wire n_4658;
 wire n_4659;
 wire n_466;
 wire n_4660;
 wire n_4661;
 wire n_4662;
 wire n_4663;
 wire n_4664;
 wire n_4665;
 wire n_4666;
 wire n_4667;
 wire n_4668;
 wire n_4669;
 wire n_467;
 wire n_4670;
 wire n_4671;
 wire n_4672;
 wire n_4673;
 wire n_4674;
 wire n_4675;
 wire n_4676;
 wire n_4677;
 wire n_4678;
 wire n_4679;
 wire n_468;
 wire n_4680;
 wire n_4681;
 wire n_4682;
 wire n_4683;
 wire n_4684;
 wire n_4685;
 wire n_4686;
 wire n_4687;
 wire n_4688;
 wire n_4689;
 wire n_469;
 wire n_4690;
 wire n_4691;
 wire n_4692;
 wire n_4693;
 wire n_4694;
 wire n_4695;
 wire n_4696;
 wire n_4697;
 wire n_4698;
 wire n_4699;
 wire n_47;
 wire n_470;
 wire n_4700;
 wire n_4701;
 wire n_4702;
 wire n_4703;
 wire n_4704;
 wire n_4705;
 wire n_4706;
 wire n_4707;
 wire n_4708;
 wire n_4709;
 wire n_471;
 wire n_4710;
 wire n_4711;
 wire n_4712;
 wire n_4713;
 wire n_4714;
 wire n_4715;
 wire n_4716;
 wire n_4717;
 wire n_4718;
 wire n_4719;
 wire n_472;
 wire n_4720;
 wire n_4721;
 wire n_4722;
 wire n_4723;
 wire n_4724;
 wire n_4725;
 wire n_4726;
 wire n_4727;
 wire n_4728;
 wire n_4729;
 wire n_473;
 wire n_4730;
 wire n_4731;
 wire n_4732;
 wire n_4733;
 wire n_4734;
 wire n_4735;
 wire n_4736;
 wire n_4737;
 wire n_4738;
 wire n_4739;
 wire n_474;
 wire n_4740;
 wire n_4741;
 wire n_4742;
 wire n_4743;
 wire n_4744;
 wire n_4745;
 wire n_4746;
 wire n_4747;
 wire n_4748;
 wire n_4749;
 wire n_475;
 wire n_4750;
 wire n_4751;
 wire n_4752;
 wire n_4753;
 wire n_4754;
 wire n_4755;
 wire n_4756;
 wire n_4757;
 wire n_4758;
 wire n_4759;
 wire n_476;
 wire n_4760;
 wire n_4761;
 wire n_4762;
 wire n_4763;
 wire n_4764;
 wire n_4765;
 wire n_4766;
 wire n_4767;
 wire n_4768;
 wire n_4769;
 wire n_477;
 wire n_4770;
 wire n_4771;
 wire n_4772;
 wire n_4773;
 wire n_4774;
 wire n_4775;
 wire n_4776;
 wire n_4777;
 wire n_4778;
 wire n_4779;
 wire n_478;
 wire n_4780;
 wire n_4781;
 wire n_4782;
 wire n_4783;
 wire n_4784;
 wire n_4785;
 wire n_4786;
 wire n_4787;
 wire n_4788;
 wire n_4789;
 wire n_479;
 wire n_4790;
 wire n_4791;
 wire n_4792;
 wire n_4793;
 wire n_4794;
 wire n_4795;
 wire n_4796;
 wire n_4797;
 wire n_4798;
 wire n_4799;
 wire n_48;
 wire n_480;
 wire n_4800;
 wire n_4801;
 wire n_4802;
 wire n_4803;
 wire n_4804;
 wire n_4805;
 wire n_4806;
 wire n_4807;
 wire n_4808;
 wire n_4809;
 wire n_481;
 wire n_4810;
 wire n_4811;
 wire n_4812;
 wire n_4813;
 wire n_4814;
 wire n_4815;
 wire n_4816;
 wire n_4817;
 wire n_4818;
 wire n_4819;
 wire n_482;
 wire n_4820;
 wire n_4821;
 wire n_4822;
 wire n_4823;
 wire n_4824;
 wire n_4825;
 wire n_4826;
 wire n_4827;
 wire n_4828;
 wire n_4829;
 wire n_483;
 wire n_4830;
 wire n_4831;
 wire n_4832;
 wire n_4833;
 wire n_4834;
 wire n_4835;
 wire n_4836;
 wire n_4837;
 wire n_4838;
 wire n_4839;
 wire n_484;
 wire n_4840;
 wire n_4841;
 wire n_4842;
 wire n_4843;
 wire n_4844;
 wire n_4845;
 wire n_4846;
 wire n_4847;
 wire n_4848;
 wire n_4849;
 wire n_485;
 wire n_4850;
 wire n_4851;
 wire n_4852;
 wire n_4853;
 wire n_4854;
 wire n_4855;
 wire n_4856;
 wire n_4857;
 wire n_4858;
 wire n_4859;
 wire n_486;
 wire n_4860;
 wire n_4861;
 wire n_4862;
 wire n_4863;
 wire n_4864;
 wire n_4865;
 wire n_4866;
 wire n_4867;
 wire n_4868;
 wire n_4869;
 wire n_487;
 wire n_4870;
 wire n_4871;
 wire n_4872;
 wire n_4873;
 wire n_4874;
 wire n_4875;
 wire n_4876;
 wire n_4877;
 wire n_4878;
 wire n_4879;
 wire n_488;
 wire n_4880;
 wire n_4881;
 wire n_4882;
 wire n_4883;
 wire n_4884;
 wire n_4885;
 wire n_4886;
 wire n_4887;
 wire n_4888;
 wire n_4889;
 wire n_489;
 wire n_4890;
 wire n_4891;
 wire n_4892;
 wire n_4893;
 wire n_4894;
 wire n_4895;
 wire n_4896;
 wire n_4897;
 wire n_4898;
 wire n_4899;
 wire n_49;
 wire n_490;
 wire n_4900;
 wire n_4901;
 wire n_4902;
 wire n_4903;
 wire n_4904;
 wire n_4905;
 wire n_4906;
 wire n_4907;
 wire n_4908;
 wire n_4909;
 wire n_491;
 wire n_4910;
 wire n_4911;
 wire n_4912;
 wire n_4913;
 wire n_4914;
 wire n_4915;
 wire n_4916;
 wire n_4917;
 wire n_4918;
 wire n_4919;
 wire n_492;
 wire n_4920;
 wire n_4921;
 wire n_4922;
 wire n_4923;
 wire n_4924;
 wire n_4925;
 wire n_4926;
 wire n_4927;
 wire n_4928;
 wire n_4929;
 wire n_493;
 wire n_4930;
 wire n_4931;
 wire n_4932;
 wire n_4933;
 wire n_4934;
 wire n_4935;
 wire n_4936;
 wire n_4937;
 wire n_4938;
 wire n_4939;
 wire n_494;
 wire n_4940;
 wire n_4941;
 wire n_4942;
 wire n_4943;
 wire n_4944;
 wire n_4945;
 wire n_4946;
 wire n_4947;
 wire n_4948;
 wire n_4949;
 wire n_495;
 wire n_4950;
 wire n_4951;
 wire n_4952;
 wire n_4953;
 wire n_4954;
 wire n_4955;
 wire n_4956;
 wire n_4957;
 wire n_4958;
 wire n_4959;
 wire n_496;
 wire n_4960;
 wire n_4961;
 wire n_4962;
 wire n_4963;
 wire n_4964;
 wire n_4965;
 wire n_4966;
 wire n_4967;
 wire n_4968;
 wire n_4969;
 wire n_497;
 wire n_4970;
 wire n_4971;
 wire n_4972;
 wire n_4973;
 wire n_4974;
 wire n_4975;
 wire n_4976;
 wire n_4977;
 wire n_4978;
 wire n_4979;
 wire n_498;
 wire n_4980;
 wire n_4981;
 wire n_4982;
 wire n_4983;
 wire n_4984;
 wire n_4985;
 wire n_4986;
 wire n_4987;
 wire n_4988;
 wire n_4989;
 wire n_499;
 wire n_4990;
 wire n_4991;
 wire n_4992;
 wire n_4993;
 wire n_4994;
 wire n_4995;
 wire n_4996;
 wire n_4997;
 wire n_4998;
 wire n_4999;
 wire n_5;
 wire n_50;
 wire n_500;
 wire n_5000;
 wire n_5001;
 wire n_5002;
 wire n_5003;
 wire n_5004;
 wire n_5005;
 wire n_5006;
 wire n_5007;
 wire n_5008;
 wire n_5009;
 wire n_501;
 wire n_5010;
 wire n_5011;
 wire n_5012;
 wire n_5013;
 wire n_5014;
 wire n_5015;
 wire n_5016;
 wire n_5017;
 wire n_5018;
 wire n_5019;
 wire n_502;
 wire n_5020;
 wire n_5021;
 wire n_5022;
 wire n_5023;
 wire n_5024;
 wire n_5025;
 wire n_5026;
 wire n_5027;
 wire n_5028;
 wire n_5029;
 wire n_503;
 wire n_5030;
 wire n_5031;
 wire n_5032;
 wire n_5033;
 wire n_5034;
 wire n_5035;
 wire n_5036;
 wire n_5037;
 wire n_5038;
 wire n_5039;
 wire n_504;
 wire n_5040;
 wire n_5041;
 wire n_5042;
 wire n_5043;
 wire n_5044;
 wire n_5045;
 wire n_5046;
 wire n_5047;
 wire n_5048;
 wire n_5049;
 wire n_505;
 wire n_5050;
 wire n_5051;
 wire n_5052;
 wire n_5053;
 wire n_5054;
 wire n_5055;
 wire n_5056;
 wire n_5057;
 wire n_5058;
 wire n_5059;
 wire n_506;
 wire n_5060;
 wire n_5061;
 wire n_5062;
 wire n_5063;
 wire n_5064;
 wire n_5065;
 wire n_5066;
 wire n_5067;
 wire n_5068;
 wire n_5069;
 wire n_507;
 wire n_5070;
 wire n_5071;
 wire n_5072;
 wire n_5073;
 wire n_5074;
 wire n_5075;
 wire n_5076;
 wire n_5077;
 wire n_5078;
 wire n_5079;
 wire n_508;
 wire n_5080;
 wire n_5081;
 wire n_5082;
 wire n_5083;
 wire n_5084;
 wire n_5085;
 wire n_5086;
 wire n_5087;
 wire n_5088;
 wire n_5089;
 wire n_509;
 wire n_5090;
 wire n_5091;
 wire n_5092;
 wire n_5093;
 wire n_5094;
 wire n_5095;
 wire n_5096;
 wire n_5097;
 wire n_5098;
 wire n_5099;
 wire n_51;
 wire n_510;
 wire n_5100;
 wire n_5101;
 wire n_5102;
 wire n_5103;
 wire n_5104;
 wire n_5105;
 wire n_5106;
 wire n_5107;
 wire n_5108;
 wire n_5109;
 wire n_511;
 wire n_5110;
 wire n_5111;
 wire n_5112;
 wire n_5113;
 wire n_5114;
 wire n_5115;
 wire n_5116;
 wire n_5117;
 wire n_5118;
 wire n_5119;
 wire n_512;
 wire n_5120;
 wire n_5121;
 wire n_5122;
 wire n_5123;
 wire n_5124;
 wire n_5125;
 wire n_5126;
 wire n_5127;
 wire n_5128;
 wire n_5129;
 wire n_513;
 wire n_5130;
 wire n_5131;
 wire n_5132;
 wire n_5133;
 wire n_5134;
 wire n_5135;
 wire n_5136;
 wire n_5137;
 wire n_5138;
 wire n_5139;
 wire n_514;
 wire n_5140;
 wire n_5141;
 wire n_5142;
 wire n_5143;
 wire n_5144;
 wire n_5145;
 wire n_5146;
 wire n_5147;
 wire n_5148;
 wire n_5149;
 wire n_515;
 wire n_5150;
 wire n_5151;
 wire n_5152;
 wire n_5153;
 wire n_5154;
 wire n_5155;
 wire n_5156;
 wire n_5157;
 wire n_5158;
 wire n_5159;
 wire n_516;
 wire n_5160;
 wire n_5161;
 wire n_5162;
 wire n_5163;
 wire n_5164;
 wire n_5165;
 wire n_5166;
 wire n_5167;
 wire n_5168;
 wire n_5169;
 wire n_517;
 wire n_5170;
 wire n_5171;
 wire n_5172;
 wire n_5173;
 wire n_5174;
 wire n_5175;
 wire n_5176;
 wire n_5177;
 wire n_5178;
 wire n_5179;
 wire n_518;
 wire n_5180;
 wire n_5181;
 wire n_5182;
 wire n_5183;
 wire n_5184;
 wire n_5185;
 wire n_5186;
 wire n_5187;
 wire n_5188;
 wire n_5189;
 wire n_519;
 wire n_5190;
 wire n_5191;
 wire n_5192;
 wire n_5193;
 wire n_5194;
 wire n_5195;
 wire n_5196;
 wire n_5197;
 wire n_5198;
 wire n_5199;
 wire n_52;
 wire n_520;
 wire n_5200;
 wire n_5201;
 wire n_5202;
 wire n_5203;
 wire n_5204;
 wire n_5205;
 wire n_5206;
 wire n_5207;
 wire n_5208;
 wire n_5209;
 wire n_521;
 wire n_5210;
 wire n_5211;
 wire n_5212;
 wire n_5213;
 wire n_5214;
 wire n_5215;
 wire n_5216;
 wire n_5217;
 wire n_5218;
 wire n_5219;
 wire n_522;
 wire n_5220;
 wire n_5221;
 wire n_5222;
 wire n_5223;
 wire n_5224;
 wire n_5225;
 wire n_5226;
 wire n_5227;
 wire n_5228;
 wire n_5229;
 wire n_523;
 wire n_5230;
 wire n_5231;
 wire n_5232;
 wire n_5233;
 wire n_5234;
 wire n_5235;
 wire n_5236;
 wire n_5237;
 wire n_5238;
 wire n_5239;
 wire n_524;
 wire n_5240;
 wire n_5241;
 wire n_5242;
 wire n_5243;
 wire n_5244;
 wire n_5245;
 wire n_5246;
 wire n_5247;
 wire n_5248;
 wire n_5249;
 wire n_525;
 wire n_5250;
 wire n_5251;
 wire n_5252;
 wire n_5253;
 wire n_5254;
 wire n_5255;
 wire n_5256;
 wire n_5257;
 wire n_5258;
 wire n_5259;
 wire n_526;
 wire n_5260;
 wire n_5261;
 wire n_5262;
 wire n_5263;
 wire n_5264;
 wire n_5265;
 wire n_5266;
 wire n_5267;
 wire n_5268;
 wire n_5269;
 wire n_527;
 wire n_5270;
 wire n_5271;
 wire n_5272;
 wire n_5273;
 wire n_5274;
 wire n_5275;
 wire n_5276;
 wire n_5277;
 wire n_5278;
 wire n_5279;
 wire n_528;
 wire n_5280;
 wire n_5281;
 wire n_5282;
 wire n_5283;
 wire n_5284;
 wire n_5285;
 wire n_5286;
 wire n_5287;
 wire n_5288;
 wire n_5289;
 wire n_529;
 wire n_5290;
 wire n_5291;
 wire n_5292;
 wire n_5293;
 wire n_5294;
 wire n_5295;
 wire n_5296;
 wire n_5297;
 wire n_5298;
 wire n_5299;
 wire n_53;
 wire n_530;
 wire n_5300;
 wire n_5301;
 wire n_5302;
 wire n_5303;
 wire n_5304;
 wire n_5305;
 wire n_5306;
 wire n_5307;
 wire n_5308;
 wire n_5309;
 wire n_531;
 wire n_5310;
 wire n_5311;
 wire n_5312;
 wire n_5313;
 wire n_5314;
 wire n_5315;
 wire n_5316;
 wire n_5317;
 wire n_5318;
 wire n_5319;
 wire n_532;
 wire n_5320;
 wire n_5321;
 wire n_5322;
 wire n_5323;
 wire n_5324;
 wire n_5325;
 wire n_5326;
 wire n_5327;
 wire n_5328;
 wire n_5329;
 wire n_533;
 wire n_5330;
 wire n_5331;
 wire n_5332;
 wire n_5333;
 wire n_5334;
 wire n_5335;
 wire n_5336;
 wire n_5337;
 wire n_5338;
 wire n_5339;
 wire n_534;
 wire n_5340;
 wire n_5341;
 wire n_5342;
 wire n_5343;
 wire n_5344;
 wire n_5345;
 wire n_5346;
 wire n_5347;
 wire n_5348;
 wire n_5349;
 wire n_535;
 wire n_5350;
 wire n_5351;
 wire n_5352;
 wire n_5353;
 wire n_5354;
 wire n_5355;
 wire n_5356;
 wire n_5357;
 wire n_5358;
 wire n_5359;
 wire n_536;
 wire n_5360;
 wire n_5361;
 wire n_5362;
 wire n_5363;
 wire n_5364;
 wire n_5365;
 wire n_5366;
 wire n_5367;
 wire n_5368;
 wire n_5369;
 wire n_537;
 wire n_5370;
 wire n_5371;
 wire n_5372;
 wire n_5373;
 wire n_5374;
 wire n_5375;
 wire n_5376;
 wire n_5377;
 wire n_5378;
 wire n_5379;
 wire n_538;
 wire n_5380;
 wire n_5381;
 wire n_5382;
 wire n_5383;
 wire n_5384;
 wire n_5385;
 wire n_5386;
 wire n_5387;
 wire n_5388;
 wire n_5389;
 wire n_539;
 wire n_5390;
 wire n_5391;
 wire n_5392;
 wire n_5393;
 wire n_5394;
 wire n_5395;
 wire n_5396;
 wire n_5397;
 wire n_5398;
 wire n_5399;
 wire n_54;
 wire n_540;
 wire n_5400;
 wire n_5401;
 wire n_5402;
 wire n_5403;
 wire n_5404;
 wire n_5405;
 wire n_5406;
 wire n_5407;
 wire n_5408;
 wire n_5409;
 wire n_541;
 wire n_5410;
 wire n_5411;
 wire n_5412;
 wire n_5413;
 wire n_5414;
 wire n_5415;
 wire n_5416;
 wire n_5417;
 wire n_5418;
 wire n_5419;
 wire n_542;
 wire n_5420;
 wire n_5421;
 wire n_5422;
 wire n_5423;
 wire n_5424;
 wire n_5425;
 wire n_5426;
 wire n_5427;
 wire n_5428;
 wire n_5429;
 wire n_543;
 wire n_5430;
 wire n_5431;
 wire n_5432;
 wire n_5433;
 wire n_5434;
 wire n_5435;
 wire n_5436;
 wire n_5437;
 wire n_5438;
 wire n_5439;
 wire n_544;
 wire n_5440;
 wire n_5441;
 wire n_5442;
 wire n_5443;
 wire n_5444;
 wire n_5445;
 wire n_5446;
 wire n_5447;
 wire n_5448;
 wire n_5449;
 wire n_545;
 wire n_5450;
 wire n_5451;
 wire n_5452;
 wire n_5453;
 wire n_5454;
 wire n_5455;
 wire n_5456;
 wire n_5457;
 wire n_5458;
 wire n_5459;
 wire n_546;
 wire n_5460;
 wire n_5461;
 wire n_5462;
 wire n_5463;
 wire n_5464;
 wire n_5465;
 wire n_5466;
 wire n_5467;
 wire n_5468;
 wire n_5469;
 wire n_547;
 wire n_5470;
 wire n_5471;
 wire n_5472;
 wire n_5473;
 wire n_5474;
 wire n_5475;
 wire n_5476;
 wire n_5477;
 wire n_5478;
 wire n_5479;
 wire n_548;
 wire n_5480;
 wire n_5481;
 wire n_5482;
 wire n_5483;
 wire n_5484;
 wire n_5485;
 wire n_5486;
 wire n_5487;
 wire n_5488;
 wire n_5489;
 wire n_549;
 wire n_5490;
 wire n_5491;
 wire n_5492;
 wire n_5493;
 wire n_5494;
 wire n_5495;
 wire n_5496;
 wire n_5497;
 wire n_5498;
 wire n_5499;
 wire n_55;
 wire n_550;
 wire n_5500;
 wire n_5501;
 wire n_5502;
 wire n_5503;
 wire n_5504;
 wire n_5505;
 wire n_5506;
 wire n_5507;
 wire n_5508;
 wire n_5509;
 wire n_551;
 wire n_5510;
 wire n_5511;
 wire n_5512;
 wire n_5513;
 wire n_5514;
 wire n_5515;
 wire n_5516;
 wire n_5517;
 wire n_5518;
 wire n_5519;
 wire n_552;
 wire n_5520;
 wire n_5521;
 wire n_5522;
 wire n_5523;
 wire n_5524;
 wire n_5525;
 wire n_5526;
 wire n_5527;
 wire n_5528;
 wire n_5529;
 wire n_553;
 wire n_5530;
 wire n_5531;
 wire n_5532;
 wire n_5533;
 wire n_5534;
 wire n_5535;
 wire n_5536;
 wire n_5537;
 wire n_5538;
 wire n_5539;
 wire n_554;
 wire n_5540;
 wire n_5541;
 wire n_5542;
 wire n_5543;
 wire n_5544;
 wire n_5545;
 wire n_5546;
 wire n_5547;
 wire n_5548;
 wire n_5549;
 wire n_555;
 wire n_5550;
 wire n_5551;
 wire n_5552;
 wire n_5553;
 wire n_5554;
 wire n_5555;
 wire n_5556;
 wire n_5557;
 wire n_5558;
 wire n_5559;
 wire n_556;
 wire n_5560;
 wire n_5561;
 wire n_5562;
 wire n_5563;
 wire n_5564;
 wire n_5565;
 wire n_5566;
 wire n_5567;
 wire n_5568;
 wire n_5569;
 wire n_557;
 wire n_5570;
 wire n_5571;
 wire n_5572;
 wire n_5573;
 wire n_5574;
 wire n_5575;
 wire n_5576;
 wire n_5577;
 wire n_5578;
 wire n_5579;
 wire n_558;
 wire n_5580;
 wire n_5581;
 wire n_5582;
 wire n_5583;
 wire n_5584;
 wire n_5585;
 wire n_5586;
 wire n_5587;
 wire n_5588;
 wire n_5589;
 wire n_559;
 wire n_5590;
 wire n_5591;
 wire n_5592;
 wire n_5593;
 wire n_5594;
 wire n_5595;
 wire n_5596;
 wire n_5597;
 wire n_5598;
 wire n_5599;
 wire n_560;
 wire n_5600;
 wire n_5601;
 wire n_5602;
 wire n_5603;
 wire n_5604;
 wire n_5605;
 wire n_5606;
 wire n_5607;
 wire n_5608;
 wire n_5609;
 wire n_561;
 wire n_5610;
 wire n_5611;
 wire n_5612;
 wire n_5613;
 wire n_5614;
 wire n_5615;
 wire n_5616;
 wire n_5617;
 wire n_5618;
 wire n_5619;
 wire n_562;
 wire n_5620;
 wire n_5621;
 wire n_5622;
 wire n_5623;
 wire n_5624;
 wire n_5625;
 wire n_5626;
 wire n_5627;
 wire n_5628;
 wire n_5629;
 wire n_563;
 wire n_5630;
 wire n_5631;
 wire n_5632;
 wire n_5633;
 wire n_5634;
 wire n_5635;
 wire n_5636;
 wire n_5637;
 wire n_5638;
 wire n_5639;
 wire n_564;
 wire n_5640;
 wire n_5641;
 wire n_5642;
 wire n_5643;
 wire n_5644;
 wire n_5645;
 wire n_5646;
 wire n_5647;
 wire n_5648;
 wire n_5649;
 wire n_565;
 wire n_5650;
 wire n_5651;
 wire n_5652;
 wire n_5653;
 wire n_5654;
 wire n_5655;
 wire n_5656;
 wire n_5657;
 wire n_5658;
 wire n_5659;
 wire n_566;
 wire n_5660;
 wire n_5661;
 wire n_5662;
 wire n_5663;
 wire n_5664;
 wire n_5665;
 wire n_5666;
 wire n_5667;
 wire n_5668;
 wire n_5669;
 wire n_5670;
 wire n_5671;
 wire n_5672;
 wire n_5673;
 wire n_5674;
 wire n_5675;
 wire n_5676;
 wire n_5677;
 wire n_5678;
 wire n_5679;
 wire n_568;
 wire n_5680;
 wire n_5681;
 wire n_5682;
 wire n_5683;
 wire n_5684;
 wire n_5685;
 wire n_5686;
 wire n_5687;
 wire n_5688;
 wire n_5689;
 wire n_569;
 wire n_5690;
 wire n_5691;
 wire n_5692;
 wire n_5693;
 wire n_5694;
 wire n_5695;
 wire n_5696;
 wire n_5697;
 wire n_5698;
 wire n_5699;
 wire n_57;
 wire n_570;
 wire n_5700;
 wire n_5701;
 wire n_5702;
 wire n_5703;
 wire n_5704;
 wire n_5705;
 wire n_5706;
 wire n_5707;
 wire n_5708;
 wire n_5709;
 wire n_571;
 wire n_5710;
 wire n_5711;
 wire n_5712;
 wire n_5713;
 wire n_5714;
 wire n_5715;
 wire n_5716;
 wire n_5717;
 wire n_5718;
 wire n_5719;
 wire n_572;
 wire n_5720;
 wire n_5721;
 wire n_5722;
 wire n_5723;
 wire n_5724;
 wire n_5725;
 wire n_5726;
 wire n_5727;
 wire n_5728;
 wire n_5729;
 wire n_573;
 wire n_5730;
 wire n_5731;
 wire n_5732;
 wire n_5733;
 wire n_5734;
 wire n_5735;
 wire n_5736;
 wire n_5737;
 wire n_5738;
 wire n_5739;
 wire n_574;
 wire n_5740;
 wire n_5741;
 wire n_5742;
 wire n_5743;
 wire n_5744;
 wire n_5745;
 wire n_5746;
 wire n_5747;
 wire n_5748;
 wire n_5749;
 wire n_575;
 wire n_5750;
 wire n_5751;
 wire n_5752;
 wire n_5753;
 wire n_5754;
 wire n_5755;
 wire n_5756;
 wire n_5757;
 wire n_5758;
 wire n_5759;
 wire n_576;
 wire n_5760;
 wire n_5761;
 wire n_5762;
 wire n_5763;
 wire n_5764;
 wire n_5765;
 wire n_5766;
 wire n_5767;
 wire n_5768;
 wire n_5769;
 wire n_577;
 wire n_5770;
 wire n_5771;
 wire n_5772;
 wire n_5773;
 wire n_5774;
 wire n_5775;
 wire n_5776;
 wire n_5777;
 wire n_5778;
 wire n_5779;
 wire n_578;
 wire n_5780;
 wire n_5781;
 wire n_5782;
 wire n_5783;
 wire n_5784;
 wire n_5785;
 wire n_5786;
 wire n_5787;
 wire n_5788;
 wire n_5789;
 wire n_579;
 wire n_5790;
 wire n_5791;
 wire n_5792;
 wire n_5793;
 wire n_5794;
 wire n_5795;
 wire n_5796;
 wire n_5797;
 wire n_5798;
 wire n_5799;
 wire n_58;
 wire n_5800;
 wire n_5801;
 wire n_5802;
 wire n_5803;
 wire n_5804;
 wire n_5805;
 wire n_5806;
 wire n_5807;
 wire n_5808;
 wire n_5809;
 wire n_581;
 wire n_5810;
 wire n_5811;
 wire n_5812;
 wire n_5813;
 wire n_5814;
 wire n_5815;
 wire n_5816;
 wire n_5817;
 wire n_5818;
 wire n_5819;
 wire n_582;
 wire n_5820;
 wire n_5821;
 wire n_5822;
 wire n_5823;
 wire n_5824;
 wire n_5825;
 wire n_5826;
 wire n_5827;
 wire n_5828;
 wire n_5829;
 wire n_583;
 wire n_5830;
 wire n_5831;
 wire n_5832;
 wire n_5833;
 wire n_5834;
 wire n_5835;
 wire n_5836;
 wire n_5837;
 wire n_5838;
 wire n_5839;
 wire n_584;
 wire n_5840;
 wire n_5841;
 wire n_5842;
 wire n_5843;
 wire n_5844;
 wire n_5845;
 wire n_5846;
 wire n_5847;
 wire n_5848;
 wire n_5849;
 wire n_585;
 wire n_5850;
 wire n_5851;
 wire n_5852;
 wire n_5853;
 wire n_5854;
 wire n_5855;
 wire n_5856;
 wire n_5857;
 wire n_5858;
 wire n_5859;
 wire n_586;
 wire n_5860;
 wire n_5861;
 wire n_5862;
 wire n_5863;
 wire n_5864;
 wire n_5865;
 wire n_5866;
 wire n_5867;
 wire n_5868;
 wire n_5869;
 wire n_587;
 wire n_5870;
 wire n_5871;
 wire n_5872;
 wire n_5873;
 wire n_5874;
 wire n_5875;
 wire n_5876;
 wire n_5877;
 wire n_5878;
 wire n_5879;
 wire n_588;
 wire n_5880;
 wire n_5881;
 wire n_5882;
 wire n_5884;
 wire n_5885;
 wire n_5886;
 wire n_5887;
 wire n_5888;
 wire n_5889;
 wire n_589;
 wire n_5890;
 wire n_5891;
 wire n_5892;
 wire n_5893;
 wire n_5894;
 wire n_5895;
 wire n_5896;
 wire n_5897;
 wire n_5898;
 wire n_5899;
 wire n_59;
 wire n_590;
 wire n_5900;
 wire n_5901;
 wire n_5902;
 wire n_5903;
 wire n_5904;
 wire n_5905;
 wire n_5906;
 wire n_5907;
 wire n_5908;
 wire n_5909;
 wire n_591;
 wire n_5910;
 wire n_5911;
 wire n_5912;
 wire n_5913;
 wire n_5914;
 wire n_5915;
 wire n_5916;
 wire n_5917;
 wire n_5918;
 wire n_5919;
 wire n_592;
 wire n_5920;
 wire n_5921;
 wire n_5922;
 wire n_5923;
 wire n_5924;
 wire n_5925;
 wire n_5926;
 wire n_5927;
 wire n_5928;
 wire n_5929;
 wire n_593;
 wire n_5930;
 wire n_5931;
 wire n_5932;
 wire n_5933;
 wire n_5934;
 wire n_5935;
 wire n_5936;
 wire n_5937;
 wire n_5938;
 wire n_5939;
 wire n_594;
 wire n_5940;
 wire n_5941;
 wire n_5942;
 wire n_5943;
 wire n_5944;
 wire n_5945;
 wire n_5946;
 wire n_5947;
 wire n_5948;
 wire n_5949;
 wire n_595;
 wire n_5950;
 wire n_5951;
 wire n_5952;
 wire n_5953;
 wire n_5954;
 wire n_5955;
 wire n_5956;
 wire n_5957;
 wire n_5958;
 wire n_5959;
 wire n_596;
 wire n_5960;
 wire n_5961;
 wire n_5962;
 wire n_5963;
 wire n_5964;
 wire n_5965;
 wire n_5966;
 wire n_5967;
 wire n_5968;
 wire n_5969;
 wire n_597;
 wire n_5970;
 wire n_5971;
 wire n_5972;
 wire n_5973;
 wire n_5974;
 wire n_5975;
 wire n_5976;
 wire n_5977;
 wire n_5978;
 wire n_5979;
 wire n_598;
 wire n_5980;
 wire n_5981;
 wire n_5982;
 wire n_5983;
 wire n_5984;
 wire n_5985;
 wire n_5986;
 wire n_5987;
 wire n_5988;
 wire n_5989;
 wire n_599;
 wire n_5990;
 wire n_5991;
 wire n_5992;
 wire n_5993;
 wire n_5994;
 wire n_5995;
 wire n_5996;
 wire n_5997;
 wire n_5998;
 wire n_5999;
 wire n_6;
 wire n_60;
 wire n_6000;
 wire n_6001;
 wire n_6002;
 wire n_6003;
 wire n_6004;
 wire n_6005;
 wire n_6006;
 wire n_6007;
 wire n_6008;
 wire n_6009;
 wire n_601;
 wire n_6010;
 wire n_6011;
 wire n_6012;
 wire n_6013;
 wire n_6014;
 wire n_6015;
 wire n_6016;
 wire n_6017;
 wire n_6018;
 wire n_6019;
 wire n_602;
 wire n_6020;
 wire n_6021;
 wire n_6022;
 wire n_6023;
 wire n_6024;
 wire n_6025;
 wire n_6026;
 wire n_6027;
 wire n_6028;
 wire n_6029;
 wire n_603;
 wire n_6030;
 wire n_6031;
 wire n_6032;
 wire n_6033;
 wire n_6034;
 wire n_6035;
 wire n_6036;
 wire n_6037;
 wire n_6038;
 wire n_6039;
 wire n_604;
 wire n_6040;
 wire n_6041;
 wire n_6042;
 wire n_6043;
 wire n_6044;
 wire n_6045;
 wire n_6046;
 wire n_6047;
 wire n_6048;
 wire n_6049;
 wire n_605;
 wire n_6050;
 wire n_6051;
 wire n_6052;
 wire n_6053;
 wire n_6054;
 wire n_6055;
 wire n_6056;
 wire n_6057;
 wire n_6058;
 wire n_6059;
 wire n_606;
 wire n_6060;
 wire n_6061;
 wire n_6062;
 wire n_6063;
 wire n_6064;
 wire n_6065;
 wire n_6066;
 wire n_6067;
 wire n_6068;
 wire n_6069;
 wire n_607;
 wire n_6070;
 wire n_6071;
 wire n_6072;
 wire n_6073;
 wire n_6074;
 wire n_6075;
 wire n_6076;
 wire n_6077;
 wire n_6078;
 wire n_6079;
 wire n_608;
 wire n_6080;
 wire n_6081;
 wire n_6082;
 wire n_6083;
 wire n_6084;
 wire n_6085;
 wire n_6086;
 wire n_6087;
 wire n_6088;
 wire n_6089;
 wire n_609;
 wire n_6090;
 wire n_6091;
 wire n_6092;
 wire n_6093;
 wire n_6094;
 wire n_6095;
 wire n_6096;
 wire n_6097;
 wire n_6098;
 wire n_6099;
 wire n_61;
 wire n_610;
 wire n_6100;
 wire n_6101;
 wire n_6102;
 wire n_6103;
 wire n_6104;
 wire n_6105;
 wire n_6106;
 wire n_6107;
 wire n_6108;
 wire n_6109;
 wire n_611;
 wire n_6110;
 wire n_6111;
 wire n_6112;
 wire n_6113;
 wire n_6114;
 wire n_6115;
 wire n_6116;
 wire n_6117;
 wire n_6118;
 wire n_6119;
 wire n_612;
 wire n_6120;
 wire n_6121;
 wire n_6122;
 wire n_6123;
 wire n_6124;
 wire n_6125;
 wire n_6126;
 wire n_6127;
 wire n_6128;
 wire n_6129;
 wire n_613;
 wire n_6130;
 wire n_6131;
 wire n_6132;
 wire n_6133;
 wire n_6134;
 wire n_6135;
 wire n_6136;
 wire n_6137;
 wire n_6138;
 wire n_6139;
 wire n_614;
 wire n_6140;
 wire n_6141;
 wire n_6142;
 wire n_6143;
 wire n_6144;
 wire n_6145;
 wire n_6146;
 wire n_6147;
 wire n_6148;
 wire n_6149;
 wire n_615;
 wire n_6150;
 wire n_6151;
 wire n_6152;
 wire n_6153;
 wire n_6154;
 wire n_6155;
 wire n_6156;
 wire n_6157;
 wire n_6158;
 wire n_6159;
 wire n_616;
 wire n_6160;
 wire n_6161;
 wire n_6162;
 wire n_6163;
 wire n_6164;
 wire n_6165;
 wire n_6166;
 wire n_6167;
 wire n_6168;
 wire n_6169;
 wire n_617;
 wire n_6170;
 wire n_6171;
 wire n_6172;
 wire n_6173;
 wire n_6174;
 wire n_6175;
 wire n_6176;
 wire n_6177;
 wire n_6178;
 wire n_6179;
 wire n_618;
 wire n_6180;
 wire n_6181;
 wire n_6182;
 wire n_6183;
 wire n_6184;
 wire n_6185;
 wire n_6186;
 wire n_6187;
 wire n_6188;
 wire n_6189;
 wire n_619;
 wire n_6190;
 wire n_6191;
 wire n_6192;
 wire n_6193;
 wire n_6194;
 wire n_6195;
 wire n_6196;
 wire n_6197;
 wire n_6198;
 wire n_6199;
 wire n_62;
 wire n_620;
 wire n_6200;
 wire n_6201;
 wire n_6202;
 wire n_6203;
 wire n_6204;
 wire n_6205;
 wire n_6206;
 wire n_6207;
 wire n_6208;
 wire n_6209;
 wire n_621;
 wire n_6210;
 wire n_6211;
 wire n_6212;
 wire n_6213;
 wire n_6214;
 wire n_6215;
 wire n_6216;
 wire n_6217;
 wire n_6218;
 wire n_6219;
 wire n_622;
 wire n_6220;
 wire n_6221;
 wire n_6222;
 wire n_6223;
 wire n_6224;
 wire n_6225;
 wire n_6226;
 wire n_6227;
 wire n_6228;
 wire n_6229;
 wire n_623;
 wire n_6230;
 wire n_6231;
 wire n_6232;
 wire n_6233;
 wire n_6234;
 wire n_6235;
 wire n_6236;
 wire n_6237;
 wire n_6238;
 wire n_6239;
 wire n_624;
 wire n_6240;
 wire n_6241;
 wire n_6242;
 wire n_6243;
 wire n_6244;
 wire n_6245;
 wire n_6246;
 wire n_6247;
 wire n_6248;
 wire n_6249;
 wire n_625;
 wire n_6250;
 wire n_6251;
 wire n_6252;
 wire n_6253;
 wire n_6254;
 wire n_6255;
 wire n_6256;
 wire n_6257;
 wire n_6258;
 wire n_6259;
 wire n_626;
 wire n_6260;
 wire n_6261;
 wire n_6262;
 wire n_6263;
 wire n_6264;
 wire n_6265;
 wire n_6266;
 wire n_6267;
 wire n_6268;
 wire n_6269;
 wire n_627;
 wire n_6270;
 wire n_6271;
 wire n_6272;
 wire n_6273;
 wire n_6274;
 wire n_6275;
 wire n_6276;
 wire n_6277;
 wire n_6278;
 wire n_6279;
 wire n_628;
 wire n_6280;
 wire n_6281;
 wire n_6282;
 wire n_6283;
 wire n_6284;
 wire n_6285;
 wire n_6286;
 wire n_6287;
 wire n_6288;
 wire n_6289;
 wire n_629;
 wire n_6290;
 wire n_6291;
 wire n_6292;
 wire n_6293;
 wire n_6294;
 wire n_6295;
 wire n_6296;
 wire n_6297;
 wire n_6298;
 wire n_6299;
 wire n_63;
 wire n_630;
 wire n_6300;
 wire n_6301;
 wire n_6302;
 wire n_6303;
 wire n_6304;
 wire n_6305;
 wire n_6306;
 wire n_6307;
 wire n_6308;
 wire n_6309;
 wire n_631;
 wire n_6310;
 wire n_6311;
 wire n_6312;
 wire n_6313;
 wire n_6314;
 wire n_6315;
 wire n_6316;
 wire n_6317;
 wire n_6318;
 wire n_6319;
 wire n_632;
 wire n_6320;
 wire n_6321;
 wire n_6322;
 wire n_6323;
 wire n_6324;
 wire n_6325;
 wire n_6326;
 wire n_6327;
 wire n_6328;
 wire n_6329;
 wire n_633;
 wire n_6330;
 wire n_6331;
 wire n_6332;
 wire n_6333;
 wire n_6334;
 wire n_6335;
 wire n_6336;
 wire n_6337;
 wire n_6338;
 wire n_6339;
 wire n_634;
 wire n_6340;
 wire n_6341;
 wire n_6342;
 wire n_6343;
 wire n_6344;
 wire n_6345;
 wire n_6346;
 wire n_6347;
 wire n_6348;
 wire n_6349;
 wire n_635;
 wire n_6350;
 wire n_6351;
 wire n_6352;
 wire n_6353;
 wire n_6354;
 wire n_6355;
 wire n_6356;
 wire n_6357;
 wire n_6358;
 wire n_6359;
 wire n_636;
 wire n_6360;
 wire n_6361;
 wire n_6362;
 wire n_6363;
 wire n_6364;
 wire n_6365;
 wire n_6366;
 wire n_6367;
 wire n_6368;
 wire n_6369;
 wire n_637;
 wire n_6370;
 wire n_6371;
 wire n_6372;
 wire n_6373;
 wire n_6374;
 wire n_6375;
 wire n_6376;
 wire n_6377;
 wire n_6378;
 wire n_6379;
 wire n_638;
 wire n_6380;
 wire n_6381;
 wire n_6382;
 wire n_6383;
 wire n_6384;
 wire n_6385;
 wire n_6386;
 wire n_6387;
 wire n_6388;
 wire n_6389;
 wire n_639;
 wire n_6390;
 wire n_6391;
 wire n_6392;
 wire n_6393;
 wire n_6394;
 wire n_6395;
 wire n_6396;
 wire n_6397;
 wire n_6398;
 wire n_6399;
 wire n_640;
 wire n_6400;
 wire n_6401;
 wire n_6402;
 wire n_6403;
 wire n_6404;
 wire n_6405;
 wire n_6406;
 wire n_6407;
 wire n_6408;
 wire n_6409;
 wire n_641;
 wire n_6410;
 wire n_6411;
 wire n_6412;
 wire n_6413;
 wire n_6414;
 wire n_6415;
 wire n_6416;
 wire n_6417;
 wire n_6418;
 wire n_6419;
 wire n_642;
 wire n_6420;
 wire n_6421;
 wire n_6422;
 wire n_6423;
 wire n_6424;
 wire n_6425;
 wire n_6426;
 wire n_6427;
 wire n_6428;
 wire n_6429;
 wire n_643;
 wire n_6430;
 wire n_6431;
 wire n_6432;
 wire n_6433;
 wire n_6434;
 wire n_6435;
 wire n_6436;
 wire n_6437;
 wire n_6438;
 wire n_6439;
 wire n_644;
 wire n_6440;
 wire n_6441;
 wire n_6442;
 wire n_6443;
 wire n_6444;
 wire n_6445;
 wire n_6446;
 wire n_6447;
 wire n_6448;
 wire n_6449;
 wire n_645;
 wire n_6450;
 wire n_6451;
 wire n_6452;
 wire n_6453;
 wire n_6454;
 wire n_6455;
 wire n_6456;
 wire n_6457;
 wire n_6458;
 wire n_6459;
 wire n_646;
 wire n_6460;
 wire n_6461;
 wire n_6462;
 wire n_6463;
 wire n_6464;
 wire n_6465;
 wire n_6466;
 wire n_6467;
 wire n_6468;
 wire n_6469;
 wire n_647;
 wire n_6470;
 wire n_6471;
 wire n_6472;
 wire n_6473;
 wire n_6474;
 wire n_6475;
 wire n_6476;
 wire n_6477;
 wire n_6478;
 wire n_6479;
 wire n_648;
 wire n_6480;
 wire n_6481;
 wire n_6482;
 wire n_6483;
 wire n_6484;
 wire n_6485;
 wire n_6486;
 wire n_6487;
 wire n_6488;
 wire n_6489;
 wire n_649;
 wire n_6490;
 wire n_6491;
 wire n_6492;
 wire n_6493;
 wire n_6494;
 wire n_6495;
 wire n_6496;
 wire n_6497;
 wire n_6498;
 wire n_6499;
 wire n_650;
 wire n_6500;
 wire n_6501;
 wire n_6502;
 wire n_6503;
 wire n_6504;
 wire n_6505;
 wire n_6506;
 wire n_6507;
 wire n_6508;
 wire n_6509;
 wire n_651;
 wire n_6510;
 wire n_6511;
 wire n_6512;
 wire n_6513;
 wire n_6514;
 wire n_6515;
 wire n_6516;
 wire n_6517;
 wire n_6518;
 wire n_6519;
 wire n_652;
 wire n_6520;
 wire n_6521;
 wire n_6522;
 wire n_6523;
 wire n_6524;
 wire n_6525;
 wire n_6526;
 wire n_6527;
 wire n_6528;
 wire n_6529;
 wire n_653;
 wire n_6530;
 wire n_6531;
 wire n_6532;
 wire n_6533;
 wire n_6534;
 wire n_6535;
 wire n_6536;
 wire n_6537;
 wire n_6538;
 wire n_6539;
 wire n_654;
 wire n_6540;
 wire n_6541;
 wire n_6542;
 wire n_6543;
 wire n_6544;
 wire n_6545;
 wire n_6546;
 wire n_6547;
 wire n_6548;
 wire n_6549;
 wire n_655;
 wire n_6550;
 wire n_6551;
 wire n_6552;
 wire n_6553;
 wire n_6554;
 wire n_6555;
 wire n_6556;
 wire n_6557;
 wire n_6558;
 wire n_6559;
 wire n_656;
 wire n_6560;
 wire n_6561;
 wire n_6562;
 wire n_6563;
 wire n_6564;
 wire n_6565;
 wire n_6566;
 wire n_6567;
 wire n_6568;
 wire n_6569;
 wire n_657;
 wire n_6570;
 wire n_6571;
 wire n_6572;
 wire n_6573;
 wire n_6574;
 wire n_6575;
 wire n_6576;
 wire n_6577;
 wire n_6578;
 wire n_6579;
 wire n_658;
 wire n_6580;
 wire n_6581;
 wire n_6582;
 wire n_6583;
 wire n_6584;
 wire n_6585;
 wire n_6586;
 wire n_6587;
 wire n_6588;
 wire n_6589;
 wire n_659;
 wire n_6590;
 wire n_6591;
 wire n_6592;
 wire n_6593;
 wire n_6594;
 wire n_6595;
 wire n_6596;
 wire n_6597;
 wire n_6598;
 wire n_6599;
 wire n_660;
 wire n_6600;
 wire n_6601;
 wire n_6602;
 wire n_6603;
 wire n_6604;
 wire n_6605;
 wire n_6606;
 wire n_6607;
 wire n_6608;
 wire n_6609;
 wire n_661;
 wire n_6610;
 wire n_6611;
 wire n_6612;
 wire n_6613;
 wire n_6614;
 wire n_6615;
 wire n_6616;
 wire n_6617;
 wire n_6618;
 wire n_6619;
 wire n_662;
 wire n_6620;
 wire n_6621;
 wire n_6622;
 wire n_6623;
 wire n_6624;
 wire n_6625;
 wire n_6626;
 wire n_6627;
 wire n_6628;
 wire n_6629;
 wire n_663;
 wire n_6630;
 wire n_6631;
 wire n_6632;
 wire n_6633;
 wire n_6634;
 wire n_6635;
 wire n_6636;
 wire n_6637;
 wire n_6638;
 wire n_6639;
 wire n_664;
 wire n_6640;
 wire n_6641;
 wire n_6642;
 wire n_6643;
 wire n_6644;
 wire n_6645;
 wire n_6646;
 wire n_6647;
 wire n_6648;
 wire n_6649;
 wire n_665;
 wire n_6650;
 wire n_6651;
 wire n_6652;
 wire n_6653;
 wire n_6654;
 wire n_6655;
 wire n_6656;
 wire n_6657;
 wire n_6658;
 wire n_6659;
 wire n_666;
 wire n_6660;
 wire n_6661;
 wire n_6662;
 wire n_6663;
 wire n_6664;
 wire n_6665;
 wire n_6666;
 wire n_6667;
 wire n_6668;
 wire n_6669;
 wire n_667;
 wire n_6670;
 wire n_6671;
 wire n_6672;
 wire n_6673;
 wire n_6674;
 wire n_6675;
 wire n_6676;
 wire n_6677;
 wire n_6678;
 wire n_6679;
 wire n_668;
 wire n_6680;
 wire n_6681;
 wire n_6682;
 wire n_6683;
 wire n_6684;
 wire n_6685;
 wire n_6686;
 wire n_6687;
 wire n_6688;
 wire n_6689;
 wire n_669;
 wire n_6690;
 wire n_6691;
 wire n_6692;
 wire n_6693;
 wire n_6694;
 wire n_6695;
 wire n_6696;
 wire n_6697;
 wire n_6698;
 wire n_6699;
 wire n_67;
 wire n_670;
 wire n_6700;
 wire n_6701;
 wire n_6702;
 wire n_6703;
 wire n_6704;
 wire n_6705;
 wire n_6706;
 wire n_6707;
 wire n_6708;
 wire n_6709;
 wire n_671;
 wire n_6710;
 wire n_6711;
 wire n_6712;
 wire n_6713;
 wire n_6714;
 wire n_6715;
 wire n_6716;
 wire n_6717;
 wire n_6718;
 wire n_6719;
 wire n_672;
 wire n_6720;
 wire n_6721;
 wire n_6722;
 wire n_6723;
 wire n_6724;
 wire n_6725;
 wire n_6726;
 wire n_6727;
 wire n_6728;
 wire n_6729;
 wire n_673;
 wire n_6730;
 wire n_6731;
 wire n_6732;
 wire n_6733;
 wire n_6734;
 wire n_6735;
 wire n_6736;
 wire n_6737;
 wire n_6738;
 wire n_6739;
 wire n_674;
 wire n_6740;
 wire n_6741;
 wire n_6742;
 wire n_6743;
 wire n_6744;
 wire n_6745;
 wire n_6746;
 wire n_6747;
 wire n_6748;
 wire n_6749;
 wire n_675;
 wire n_6750;
 wire n_6751;
 wire n_6752;
 wire n_6753;
 wire n_6754;
 wire n_6755;
 wire n_6756;
 wire n_6757;
 wire n_6758;
 wire n_6759;
 wire n_676;
 wire n_6760;
 wire n_6761;
 wire n_6762;
 wire n_6763;
 wire n_6764;
 wire n_6765;
 wire n_6766;
 wire n_6767;
 wire n_6768;
 wire n_6769;
 wire n_677;
 wire n_6770;
 wire n_6771;
 wire n_6772;
 wire n_6773;
 wire n_6774;
 wire n_6775;
 wire n_6776;
 wire n_6777;
 wire n_6778;
 wire n_6779;
 wire n_678;
 wire n_6780;
 wire n_6781;
 wire n_6782;
 wire n_6783;
 wire n_6784;
 wire n_6785;
 wire n_6786;
 wire n_6787;
 wire n_6788;
 wire n_6789;
 wire n_679;
 wire n_6790;
 wire n_6791;
 wire n_6792;
 wire n_6793;
 wire n_6794;
 wire n_6795;
 wire n_6796;
 wire n_6797;
 wire n_6798;
 wire n_6799;
 wire n_68;
 wire n_680;
 wire n_6800;
 wire n_6801;
 wire n_6802;
 wire n_6803;
 wire n_6804;
 wire n_6805;
 wire n_6806;
 wire n_6807;
 wire n_6808;
 wire n_6809;
 wire n_681;
 wire n_6810;
 wire n_6811;
 wire n_6812;
 wire n_6813;
 wire n_6814;
 wire n_6815;
 wire n_6816;
 wire n_6817;
 wire n_6818;
 wire n_6819;
 wire n_682;
 wire n_6820;
 wire n_6821;
 wire n_6822;
 wire n_6823;
 wire n_6824;
 wire n_6825;
 wire n_6826;
 wire n_6827;
 wire n_6828;
 wire n_6829;
 wire n_683;
 wire n_6830;
 wire n_6832;
 wire n_6833;
 wire n_6834;
 wire n_6835;
 wire n_6836;
 wire n_6837;
 wire n_6838;
 wire n_6839;
 wire n_684;
 wire n_6840;
 wire n_6841;
 wire n_6842;
 wire n_6843;
 wire n_6844;
 wire n_6845;
 wire n_6846;
 wire n_6847;
 wire n_6848;
 wire n_6849;
 wire n_685;
 wire n_6850;
 wire n_6851;
 wire n_6852;
 wire n_6853;
 wire n_6854;
 wire n_6855;
 wire n_6856;
 wire n_6857;
 wire n_6858;
 wire n_6859;
 wire n_686;
 wire n_6860;
 wire n_6861;
 wire n_6862;
 wire n_6863;
 wire n_6864;
 wire n_6865;
 wire n_6866;
 wire n_6867;
 wire n_6868;
 wire n_6869;
 wire n_687;
 wire n_6870;
 wire n_6871;
 wire n_6872;
 wire n_6873;
 wire n_6874;
 wire n_6875;
 wire n_6876;
 wire n_6877;
 wire n_6878;
 wire n_6879;
 wire n_688;
 wire n_6880;
 wire n_6881;
 wire n_6882;
 wire n_6883;
 wire n_6884;
 wire n_6885;
 wire n_6886;
 wire n_6887;
 wire n_6888;
 wire n_6889;
 wire n_689;
 wire n_6890;
 wire n_6891;
 wire n_6892;
 wire n_6893;
 wire n_6894;
 wire n_6895;
 wire n_6896;
 wire n_6897;
 wire n_6898;
 wire n_6899;
 wire n_69;
 wire n_690;
 wire n_6900;
 wire n_6901;
 wire n_6902;
 wire n_6903;
 wire n_6904;
 wire n_6905;
 wire n_6906;
 wire n_6907;
 wire n_6908;
 wire n_6909;
 wire n_691;
 wire n_6910;
 wire n_6911;
 wire n_6912;
 wire n_6913;
 wire n_6914;
 wire n_6915;
 wire n_6916;
 wire n_6917;
 wire n_6918;
 wire n_6919;
 wire n_692;
 wire n_6920;
 wire n_6921;
 wire n_6922;
 wire n_6923;
 wire n_6924;
 wire n_6925;
 wire n_6926;
 wire n_6927;
 wire n_6928;
 wire n_6929;
 wire n_693;
 wire n_6930;
 wire n_6931;
 wire n_6932;
 wire n_6933;
 wire n_6934;
 wire n_6935;
 wire n_6936;
 wire n_6937;
 wire n_6938;
 wire n_6939;
 wire n_6940;
 wire n_6941;
 wire n_6942;
 wire n_6943;
 wire n_6944;
 wire n_6945;
 wire n_6946;
 wire n_6947;
 wire n_6948;
 wire n_6949;
 wire n_695;
 wire n_6950;
 wire n_6951;
 wire n_6952;
 wire n_6953;
 wire n_6954;
 wire n_6955;
 wire n_6956;
 wire n_6957;
 wire n_6958;
 wire n_6959;
 wire n_696;
 wire n_6960;
 wire n_6961;
 wire n_6962;
 wire n_6963;
 wire n_6964;
 wire n_6965;
 wire n_6966;
 wire n_6967;
 wire n_6968;
 wire n_6969;
 wire n_697;
 wire n_6970;
 wire n_6971;
 wire n_6972;
 wire n_6973;
 wire n_6974;
 wire n_6975;
 wire n_6976;
 wire n_6977;
 wire n_6978;
 wire n_6979;
 wire n_698;
 wire n_6980;
 wire n_6981;
 wire n_6982;
 wire n_6983;
 wire n_6984;
 wire n_6985;
 wire n_6986;
 wire n_6987;
 wire n_6988;
 wire n_6989;
 wire n_699;
 wire n_6990;
 wire n_6991;
 wire n_6992;
 wire n_6993;
 wire n_6994;
 wire n_6995;
 wire n_6996;
 wire n_6997;
 wire n_6998;
 wire n_6999;
 wire n_7;
 wire n_70;
 wire n_700;
 wire n_7000;
 wire n_7001;
 wire n_7002;
 wire n_7003;
 wire n_7004;
 wire n_7005;
 wire n_7006;
 wire n_7007;
 wire n_7008;
 wire n_7009;
 wire n_701;
 wire n_7010;
 wire n_7011;
 wire n_7012;
 wire n_7013;
 wire n_7014;
 wire n_7015;
 wire n_7016;
 wire n_7017;
 wire n_7018;
 wire n_7019;
 wire n_702;
 wire n_7020;
 wire n_7021;
 wire n_7022;
 wire n_7023;
 wire n_7024;
 wire n_7025;
 wire n_7026;
 wire n_7027;
 wire n_7028;
 wire n_7029;
 wire n_703;
 wire n_7030;
 wire n_7031;
 wire n_7032;
 wire n_7033;
 wire n_7034;
 wire n_7035;
 wire n_7036;
 wire n_7037;
 wire n_7038;
 wire n_7039;
 wire n_704;
 wire n_7040;
 wire n_7041;
 wire n_7042;
 wire n_7043;
 wire n_7044;
 wire n_7045;
 wire n_7046;
 wire n_7047;
 wire n_7048;
 wire n_7049;
 wire n_705;
 wire n_7050;
 wire n_7051;
 wire n_7052;
 wire n_7053;
 wire n_7054;
 wire n_7055;
 wire n_7056;
 wire n_7057;
 wire n_7058;
 wire n_7059;
 wire n_706;
 wire n_7060;
 wire n_7061;
 wire n_7062;
 wire n_7063;
 wire n_7064;
 wire n_7065;
 wire n_7066;
 wire n_7067;
 wire n_7068;
 wire n_7069;
 wire n_707;
 wire n_7070;
 wire n_7071;
 wire n_7072;
 wire n_7073;
 wire n_7074;
 wire n_7075;
 wire n_7076;
 wire n_7077;
 wire n_7078;
 wire n_7079;
 wire n_708;
 wire n_7080;
 wire n_7082;
 wire n_7083;
 wire n_7084;
 wire n_7085;
 wire n_7086;
 wire n_7087;
 wire n_7088;
 wire n_7089;
 wire n_709;
 wire n_7090;
 wire n_7091;
 wire n_7092;
 wire n_7093;
 wire n_7094;
 wire n_7095;
 wire n_7096;
 wire n_7097;
 wire n_7098;
 wire n_7099;
 wire n_71;
 wire n_710;
 wire n_7100;
 wire n_7101;
 wire n_7102;
 wire n_7103;
 wire n_7104;
 wire n_7105;
 wire n_7106;
 wire n_7107;
 wire n_7108;
 wire n_7109;
 wire n_711;
 wire n_7110;
 wire n_7111;
 wire n_7112;
 wire n_7113;
 wire n_7114;
 wire n_7115;
 wire n_7116;
 wire n_7117;
 wire n_7118;
 wire n_7119;
 wire n_712;
 wire n_7120;
 wire n_7121;
 wire n_7122;
 wire n_7123;
 wire n_7124;
 wire n_7125;
 wire n_7126;
 wire n_7127;
 wire n_7128;
 wire n_7129;
 wire n_713;
 wire n_7130;
 wire n_7131;
 wire n_7132;
 wire n_7133;
 wire n_7134;
 wire n_7135;
 wire n_7136;
 wire n_7137;
 wire n_7138;
 wire n_7139;
 wire n_714;
 wire n_7140;
 wire n_7141;
 wire n_7142;
 wire n_7143;
 wire n_7144;
 wire n_7145;
 wire n_7146;
 wire n_7147;
 wire n_7148;
 wire n_7149;
 wire n_715;
 wire n_7150;
 wire n_7151;
 wire n_7152;
 wire n_7153;
 wire n_7154;
 wire n_7155;
 wire n_7156;
 wire n_7157;
 wire n_7158;
 wire n_7159;
 wire n_716;
 wire n_7160;
 wire n_7161;
 wire n_7162;
 wire n_7163;
 wire n_7164;
 wire n_7165;
 wire n_7166;
 wire n_7167;
 wire n_7168;
 wire n_7169;
 wire n_717;
 wire n_7170;
 wire n_7171;
 wire n_7172;
 wire n_7173;
 wire n_7174;
 wire n_7175;
 wire n_7176;
 wire n_7177;
 wire n_7178;
 wire n_7179;
 wire n_718;
 wire n_7180;
 wire n_7181;
 wire n_7182;
 wire n_7183;
 wire n_7184;
 wire n_7185;
 wire n_7186;
 wire n_7187;
 wire n_7188;
 wire n_7189;
 wire n_719;
 wire n_7190;
 wire n_7191;
 wire n_7192;
 wire n_7193;
 wire n_7194;
 wire n_7195;
 wire n_7196;
 wire n_7197;
 wire n_7198;
 wire n_7199;
 wire n_72;
 wire n_720;
 wire n_7200;
 wire n_7201;
 wire n_7202;
 wire n_7203;
 wire n_7204;
 wire n_7205;
 wire n_7206;
 wire n_7207;
 wire n_7208;
 wire n_7209;
 wire n_721;
 wire n_7210;
 wire n_7211;
 wire n_7212;
 wire n_7213;
 wire n_7214;
 wire n_7215;
 wire n_7216;
 wire n_7217;
 wire n_7218;
 wire n_7219;
 wire n_722;
 wire n_7220;
 wire n_7221;
 wire n_7222;
 wire n_7223;
 wire n_7224;
 wire n_7225;
 wire n_7226;
 wire n_7227;
 wire n_7228;
 wire n_7229;
 wire n_723;
 wire n_7230;
 wire n_7231;
 wire n_7232;
 wire n_7233;
 wire n_7234;
 wire n_7235;
 wire n_7236;
 wire n_7237;
 wire n_7238;
 wire n_7239;
 wire n_724;
 wire n_7240;
 wire n_7241;
 wire n_7242;
 wire n_7243;
 wire n_7244;
 wire n_7245;
 wire n_7246;
 wire n_7247;
 wire n_7248;
 wire n_7249;
 wire n_725;
 wire n_7250;
 wire n_7251;
 wire n_7252;
 wire n_7253;
 wire n_7254;
 wire n_7255;
 wire n_7256;
 wire n_7258;
 wire n_7259;
 wire n_726;
 wire n_7260;
 wire n_7261;
 wire n_7262;
 wire n_7263;
 wire n_7264;
 wire n_7265;
 wire n_7266;
 wire n_7267;
 wire n_7268;
 wire n_7269;
 wire n_727;
 wire n_7270;
 wire n_7271;
 wire n_7272;
 wire n_7273;
 wire n_7274;
 wire n_7275;
 wire n_7276;
 wire n_7277;
 wire n_7278;
 wire n_7279;
 wire n_728;
 wire n_7280;
 wire n_7281;
 wire n_7282;
 wire n_7283;
 wire n_7284;
 wire n_7285;
 wire n_7286;
 wire n_7287;
 wire n_7288;
 wire n_7289;
 wire n_729;
 wire n_7290;
 wire n_7291;
 wire n_7292;
 wire n_7293;
 wire n_7294;
 wire n_7295;
 wire n_7296;
 wire n_7297;
 wire n_7298;
 wire n_7299;
 wire n_73;
 wire n_7300;
 wire n_7301;
 wire n_7302;
 wire n_7303;
 wire n_7304;
 wire n_7305;
 wire n_7306;
 wire n_7307;
 wire n_7308;
 wire n_7309;
 wire n_731;
 wire n_7310;
 wire n_7311;
 wire n_7312;
 wire n_7313;
 wire n_7314;
 wire n_7315;
 wire n_7316;
 wire n_7317;
 wire n_7318;
 wire n_7319;
 wire n_732;
 wire n_7320;
 wire n_7321;
 wire n_7322;
 wire n_7323;
 wire n_7324;
 wire n_7325;
 wire n_7326;
 wire n_7327;
 wire n_7328;
 wire n_7329;
 wire n_733;
 wire n_7330;
 wire n_7331;
 wire n_7332;
 wire n_7333;
 wire n_7334;
 wire n_7335;
 wire n_7336;
 wire n_7337;
 wire n_7338;
 wire n_7339;
 wire n_734;
 wire n_7340;
 wire n_7341;
 wire n_7342;
 wire n_7343;
 wire n_7344;
 wire n_7345;
 wire n_7346;
 wire n_7347;
 wire n_7348;
 wire n_7349;
 wire n_735;
 wire n_7350;
 wire n_7351;
 wire n_7352;
 wire n_7353;
 wire n_7354;
 wire n_7355;
 wire n_7356;
 wire n_7357;
 wire n_7358;
 wire n_7359;
 wire n_736;
 wire n_7360;
 wire n_7361;
 wire n_7362;
 wire n_7363;
 wire n_7364;
 wire n_7365;
 wire n_7366;
 wire n_7367;
 wire n_7368;
 wire n_7369;
 wire n_737;
 wire n_7370;
 wire n_7371;
 wire n_7372;
 wire n_7373;
 wire n_7374;
 wire n_7375;
 wire n_7376;
 wire n_7377;
 wire n_7378;
 wire n_7379;
 wire n_738;
 wire n_7380;
 wire n_7381;
 wire n_7382;
 wire n_7383;
 wire n_7384;
 wire n_7385;
 wire n_7386;
 wire n_7387;
 wire n_7388;
 wire n_7389;
 wire n_739;
 wire n_7390;
 wire n_7391;
 wire n_7392;
 wire n_7393;
 wire n_7394;
 wire n_7395;
 wire n_7396;
 wire n_7397;
 wire n_7398;
 wire n_7399;
 wire n_74;
 wire n_740;
 wire n_7400;
 wire n_7401;
 wire n_7402;
 wire n_7403;
 wire n_7404;
 wire n_7405;
 wire n_7406;
 wire n_7407;
 wire n_7408;
 wire n_741;
 wire n_7410;
 wire n_7411;
 wire n_7412;
 wire n_7413;
 wire n_7414;
 wire n_7415;
 wire n_7416;
 wire n_7417;
 wire n_7418;
 wire n_7419;
 wire n_742;
 wire n_7420;
 wire n_7421;
 wire n_7422;
 wire n_7423;
 wire n_7424;
 wire n_7425;
 wire n_7426;
 wire n_7427;
 wire n_7428;
 wire n_7429;
 wire n_743;
 wire n_7430;
 wire n_7431;
 wire n_7432;
 wire n_7433;
 wire n_7434;
 wire n_7435;
 wire n_7436;
 wire n_7437;
 wire n_7438;
 wire n_7439;
 wire n_744;
 wire n_7440;
 wire n_7441;
 wire n_7442;
 wire n_7443;
 wire n_7444;
 wire n_7445;
 wire n_7446;
 wire n_7447;
 wire n_7448;
 wire n_745;
 wire n_7450;
 wire n_7451;
 wire n_7453;
 wire n_7454;
 wire n_7455;
 wire n_7456;
 wire n_7457;
 wire n_7458;
 wire n_7459;
 wire n_746;
 wire n_7460;
 wire n_7461;
 wire n_7462;
 wire n_7463;
 wire n_7464;
 wire n_7465;
 wire n_7466;
 wire n_7467;
 wire n_7468;
 wire n_7469;
 wire n_747;
 wire n_7470;
 wire n_7471;
 wire n_7472;
 wire n_7474;
 wire n_7475;
 wire n_7477;
 wire n_7479;
 wire n_748;
 wire n_7480;
 wire n_7481;
 wire n_7482;
 wire n_749;
 wire n_7491;
 wire n_7492;
 wire n_7494;
 wire n_7495;
 wire n_75;
 wire n_750;
 wire n_7502;
 wire n_7503;
 wire n_7507;
 wire n_751;
 wire n_7513;
 wire n_7514;
 wire n_7518;
 wire n_7519;
 wire n_752;
 wire n_7522;
 wire n_7523;
 wire n_7524;
 wire n_7525;
 wire n_7526;
 wire n_7527;
 wire n_7528;
 wire n_7529;
 wire n_753;
 wire n_7533;
 wire n_7537;
 wire n_7539;
 wire n_754;
 wire n_7540;
 wire n_7541;
 wire n_7542;
 wire n_7546;
 wire n_7547;
 wire n_7548;
 wire n_7549;
 wire n_755;
 wire n_7550;
 wire n_7554;
 wire n_7555;
 wire n_7556;
 wire n_756;
 wire n_7560;
 wire n_7564;
 wire n_7565;
 wire n_757;
 wire n_7573;
 wire n_7574;
 wire n_758;
 wire n_7584;
 wire n_7585;
 wire n_7588;
 wire n_7589;
 wire n_759;
 wire n_7592;
 wire n_7593;
 wire n_76;
 wire n_760;
 wire n_7602;
 wire n_7605;
 wire n_7606;
 wire n_7607;
 wire n_7608;
 wire n_7609;
 wire n_761;
 wire n_7610;
 wire n_7611;
 wire n_7612;
 wire n_7613;
 wire n_7614;
 wire n_7615;
 wire n_7616;
 wire n_7617;
 wire n_7618;
 wire n_7619;
 wire n_762;
 wire n_7620;
 wire n_7621;
 wire n_7622;
 wire n_7623;
 wire n_7624;
 wire n_7625;
 wire n_7626;
 wire n_7627;
 wire n_7628;
 wire n_7629;
 wire n_763;
 wire n_7630;
 wire n_7631;
 wire n_7632;
 wire n_7633;
 wire n_7634;
 wire n_7635;
 wire n_7636;
 wire n_7637;
 wire n_7638;
 wire n_7639;
 wire n_764;
 wire n_7640;
 wire n_7641;
 wire n_7642;
 wire n_7643;
 wire n_7644;
 wire n_7645;
 wire n_7646;
 wire n_7647;
 wire n_7648;
 wire n_7649;
 wire n_765;
 wire n_7650;
 wire n_7651;
 wire n_7652;
 wire n_7653;
 wire n_7654;
 wire n_7657;
 wire n_7658;
 wire n_7659;
 wire n_766;
 wire n_7660;
 wire n_7661;
 wire n_7662;
 wire n_7663;
 wire n_7664;
 wire n_7665;
 wire n_7666;
 wire n_7667;
 wire n_7668;
 wire n_7669;
 wire n_767;
 wire n_7670;
 wire n_7671;
 wire n_7672;
 wire n_7673;
 wire n_7674;
 wire n_7675;
 wire n_7676;
 wire n_7677;
 wire n_7678;
 wire n_7679;
 wire n_768;
 wire n_7680;
 wire n_7681;
 wire n_7682;
 wire n_7683;
 wire n_7684;
 wire n_7685;
 wire n_7686;
 wire n_7687;
 wire n_7688;
 wire n_7689;
 wire n_769;
 wire n_7690;
 wire n_7691;
 wire n_7692;
 wire n_7693;
 wire n_7694;
 wire n_7695;
 wire n_7696;
 wire n_7697;
 wire n_7698;
 wire n_7699;
 wire n_77;
 wire n_770;
 wire n_7700;
 wire n_7701;
 wire n_7702;
 wire n_7703;
 wire n_7704;
 wire n_7705;
 wire n_7706;
 wire n_7707;
 wire n_7708;
 wire n_7709;
 wire n_771;
 wire n_7710;
 wire n_7711;
 wire n_7712;
 wire n_7713;
 wire n_7716;
 wire n_7717;
 wire n_7718;
 wire n_7719;
 wire n_772;
 wire n_7720;
 wire n_7721;
 wire n_7722;
 wire n_7723;
 wire n_7724;
 wire n_7725;
 wire n_7726;
 wire n_7727;
 wire n_7728;
 wire n_7729;
 wire n_773;
 wire n_7730;
 wire n_7731;
 wire n_7732;
 wire n_7733;
 wire n_7734;
 wire n_7735;
 wire n_7736;
 wire n_7737;
 wire n_7738;
 wire n_7739;
 wire n_774;
 wire n_7740;
 wire n_7741;
 wire n_7742;
 wire n_7743;
 wire n_7744;
 wire n_7745;
 wire n_7746;
 wire n_7747;
 wire n_7748;
 wire n_7749;
 wire n_775;
 wire n_7750;
 wire n_7751;
 wire n_7752;
 wire n_7753;
 wire n_7754;
 wire n_7755;
 wire n_7756;
 wire n_7757;
 wire n_7758;
 wire n_7759;
 wire n_776;
 wire n_7760;
 wire n_7761;
 wire n_7762;
 wire n_7763;
 wire n_7764;
 wire n_7765;
 wire n_7766;
 wire n_7767;
 wire n_7768;
 wire n_7769;
 wire n_777;
 wire n_7770;
 wire n_7771;
 wire n_7772;
 wire n_7773;
 wire n_7774;
 wire n_7775;
 wire n_7776;
 wire n_7777;
 wire n_7778;
 wire n_7779;
 wire n_778;
 wire n_7780;
 wire n_7781;
 wire n_7782;
 wire n_7783;
 wire n_7784;
 wire n_7785;
 wire n_7786;
 wire n_7787;
 wire n_7788;
 wire n_7789;
 wire n_779;
 wire n_7790;
 wire n_7791;
 wire n_7792;
 wire n_7793;
 wire n_7794;
 wire n_7795;
 wire n_7796;
 wire n_7797;
 wire n_7798;
 wire n_7799;
 wire n_78;
 wire n_780;
 wire n_7800;
 wire n_7801;
 wire n_7802;
 wire n_7803;
 wire n_7804;
 wire n_7805;
 wire n_7806;
 wire n_7807;
 wire n_7808;
 wire n_7809;
 wire n_781;
 wire n_7810;
 wire n_7811;
 wire n_7812;
 wire n_7813;
 wire n_7814;
 wire n_7815;
 wire n_7816;
 wire n_7817;
 wire n_7818;
 wire n_7819;
 wire n_782;
 wire n_7820;
 wire n_7821;
 wire n_7822;
 wire n_7823;
 wire n_7824;
 wire n_7825;
 wire n_7826;
 wire n_7827;
 wire n_7828;
 wire n_7829;
 wire n_783;
 wire n_7830;
 wire n_7831;
 wire n_7832;
 wire n_7833;
 wire n_7834;
 wire n_7835;
 wire n_7836;
 wire n_7837;
 wire n_7838;
 wire n_7839;
 wire n_784;
 wire n_7840;
 wire n_7841;
 wire n_7842;
 wire n_7843;
 wire n_7844;
 wire n_7845;
 wire n_7846;
 wire n_7847;
 wire n_7848;
 wire n_7849;
 wire n_785;
 wire n_7850;
 wire n_7851;
 wire n_7852;
 wire n_7853;
 wire n_7854;
 wire n_7855;
 wire n_7856;
 wire n_7857;
 wire n_7858;
 wire n_7859;
 wire n_786;
 wire n_7860;
 wire n_7861;
 wire n_7862;
 wire n_7863;
 wire n_7864;
 wire n_7865;
 wire n_7866;
 wire n_7867;
 wire n_7869;
 wire n_787;
 wire n_7870;
 wire n_7871;
 wire n_7872;
 wire n_7873;
 wire n_7874;
 wire n_7875;
 wire n_7876;
 wire n_7877;
 wire n_7878;
 wire n_788;
 wire n_7880;
 wire n_7881;
 wire n_7882;
 wire n_7883;
 wire n_7884;
 wire n_7885;
 wire n_7886;
 wire n_7887;
 wire n_7888;
 wire n_7889;
 wire n_789;
 wire n_7890;
 wire n_7891;
 wire n_7892;
 wire n_7893;
 wire n_7894;
 wire n_7895;
 wire n_7896;
 wire n_7897;
 wire n_7898;
 wire n_79;
 wire n_790;
 wire n_7900;
 wire n_7901;
 wire n_7902;
 wire n_7903;
 wire n_7904;
 wire n_7905;
 wire n_7906;
 wire n_7907;
 wire n_7908;
 wire n_7909;
 wire n_791;
 wire n_7911;
 wire n_7912;
 wire n_7913;
 wire n_7914;
 wire n_7915;
 wire n_7916;
 wire n_7917;
 wire n_7918;
 wire n_7919;
 wire n_792;
 wire n_7921;
 wire n_7922;
 wire n_7923;
 wire n_7924;
 wire n_7925;
 wire n_7926;
 wire n_7927;
 wire n_793;
 wire n_7931;
 wire n_7932;
 wire n_7935;
 wire n_7936;
 wire n_794;
 wire n_7943;
 wire n_7945;
 wire n_7946;
 wire n_7947;
 wire n_7948;
 wire n_7949;
 wire n_795;
 wire n_7950;
 wire n_7951;
 wire n_7952;
 wire n_7953;
 wire n_7954;
 wire n_7955;
 wire n_7956;
 wire n_7957;
 wire n_7958;
 wire n_7959;
 wire n_796;
 wire n_7960;
 wire n_7961;
 wire n_7962;
 wire n_7963;
 wire n_7964;
 wire n_7965;
 wire n_7966;
 wire n_7967;
 wire n_7968;
 wire n_7969;
 wire n_797;
 wire n_7970;
 wire n_7971;
 wire n_7972;
 wire n_7973;
 wire n_7974;
 wire n_7975;
 wire n_7976;
 wire n_7977;
 wire n_7978;
 wire n_7979;
 wire n_798;
 wire n_7980;
 wire n_7981;
 wire n_7982;
 wire n_7983;
 wire n_7984;
 wire n_7985;
 wire n_7986;
 wire n_7987;
 wire n_7988;
 wire n_7989;
 wire n_799;
 wire n_7990;
 wire n_7991;
 wire n_7992;
 wire n_7993;
 wire n_7994;
 wire n_7995;
 wire n_7996;
 wire n_7997;
 wire n_7998;
 wire n_7999;
 wire n_8;
 wire n_80;
 wire n_800;
 wire n_8000;
 wire n_8001;
 wire n_8002;
 wire n_8003;
 wire n_8004;
 wire n_8005;
 wire n_8006;
 wire n_8007;
 wire n_8008;
 wire n_8009;
 wire n_801;
 wire n_8010;
 wire n_8011;
 wire n_8012;
 wire n_8013;
 wire n_8014;
 wire n_8015;
 wire n_8016;
 wire n_8017;
 wire n_8018;
 wire n_8019;
 wire n_802;
 wire n_8020;
 wire n_8021;
 wire n_8022;
 wire n_8023;
 wire n_8024;
 wire n_8025;
 wire n_8026;
 wire n_8027;
 wire n_8028;
 wire n_8029;
 wire n_803;
 wire n_8030;
 wire n_8031;
 wire n_8032;
 wire n_8033;
 wire n_8034;
 wire n_8035;
 wire n_8036;
 wire n_8037;
 wire n_8038;
 wire n_8039;
 wire n_804;
 wire n_8040;
 wire n_8041;
 wire n_8042;
 wire n_8043;
 wire n_8044;
 wire n_8045;
 wire n_8046;
 wire n_8047;
 wire n_8048;
 wire n_8049;
 wire n_805;
 wire n_8050;
 wire n_8051;
 wire n_8052;
 wire n_8053;
 wire n_8054;
 wire n_8055;
 wire n_8056;
 wire n_8057;
 wire n_8058;
 wire n_8059;
 wire n_806;
 wire n_8060;
 wire n_8061;
 wire n_8062;
 wire n_8063;
 wire n_8064;
 wire n_8065;
 wire n_8066;
 wire n_8067;
 wire n_8068;
 wire n_8069;
 wire n_807;
 wire n_8070;
 wire n_8071;
 wire n_8072;
 wire n_8073;
 wire n_8074;
 wire n_8075;
 wire n_8076;
 wire n_8077;
 wire n_8078;
 wire n_8079;
 wire n_808;
 wire n_8080;
 wire n_8081;
 wire n_8082;
 wire n_8083;
 wire n_8084;
 wire n_8085;
 wire n_8086;
 wire n_8087;
 wire n_8088;
 wire n_8089;
 wire n_809;
 wire n_8090;
 wire n_8091;
 wire n_8092;
 wire n_8093;
 wire n_8094;
 wire n_8095;
 wire n_8096;
 wire n_8097;
 wire n_8098;
 wire n_8099;
 wire n_81;
 wire n_810;
 wire n_8100;
 wire n_8101;
 wire n_8102;
 wire n_8103;
 wire n_8104;
 wire n_8105;
 wire n_8106;
 wire n_8107;
 wire n_8108;
 wire n_8109;
 wire n_811;
 wire n_8110;
 wire n_8111;
 wire n_8112;
 wire n_8113;
 wire n_8114;
 wire n_8115;
 wire n_8116;
 wire n_8117;
 wire n_8118;
 wire n_8119;
 wire n_812;
 wire n_8120;
 wire n_8121;
 wire n_8122;
 wire n_8123;
 wire n_8124;
 wire n_8125;
 wire n_8126;
 wire n_8127;
 wire n_8128;
 wire n_8129;
 wire n_813;
 wire n_8130;
 wire n_8131;
 wire n_8132;
 wire n_8133;
 wire n_8134;
 wire n_8135;
 wire n_8136;
 wire n_8137;
 wire n_8138;
 wire n_8139;
 wire n_814;
 wire n_8140;
 wire n_8141;
 wire n_8142;
 wire n_8143;
 wire n_8144;
 wire n_8145;
 wire n_8146;
 wire n_8147;
 wire n_8148;
 wire n_8149;
 wire n_815;
 wire n_8150;
 wire n_8151;
 wire n_8152;
 wire n_8153;
 wire n_8154;
 wire n_8155;
 wire n_8156;
 wire n_8157;
 wire n_8158;
 wire n_8159;
 wire n_816;
 wire n_8160;
 wire n_8161;
 wire n_8162;
 wire n_8163;
 wire n_8164;
 wire n_8165;
 wire n_8166;
 wire n_8167;
 wire n_8169;
 wire n_817;
 wire n_8177;
 wire n_8178;
 wire n_8179;
 wire n_818;
 wire n_8180;
 wire n_8181;
 wire n_8182;
 wire n_8183;
 wire n_8184;
 wire n_8186;
 wire n_8187;
 wire n_8188;
 wire n_8189;
 wire n_819;
 wire n_8190;
 wire n_8191;
 wire n_8192;
 wire n_8195;
 wire n_8196;
 wire n_8197;
 wire n_8198;
 wire n_8199;
 wire n_82;
 wire n_820;
 wire n_8200;
 wire n_8202;
 wire n_8203;
 wire n_8204;
 wire n_8205;
 wire n_8206;
 wire n_8207;
 wire n_8208;
 wire n_8209;
 wire n_821;
 wire n_8210;
 wire n_8211;
 wire n_8212;
 wire n_8213;
 wire n_8214;
 wire n_8215;
 wire n_8217;
 wire n_8218;
 wire n_8219;
 wire n_822;
 wire n_8220;
 wire n_8221;
 wire n_8222;
 wire n_8224;
 wire n_8225;
 wire n_8226;
 wire n_8227;
 wire n_8228;
 wire n_8229;
 wire n_823;
 wire n_8230;
 wire n_8231;
 wire n_8232;
 wire n_8234;
 wire n_8235;
 wire n_8236;
 wire n_8238;
 wire n_8239;
 wire n_824;
 wire n_8240;
 wire n_8241;
 wire n_8242;
 wire n_8243;
 wire n_8244;
 wire n_8245;
 wire n_8246;
 wire n_8247;
 wire n_8248;
 wire n_8249;
 wire n_825;
 wire n_8250;
 wire n_8252;
 wire n_8253;
 wire n_8254;
 wire n_8255;
 wire n_8256;
 wire n_8258;
 wire n_8259;
 wire n_826;
 wire n_8260;
 wire n_8261;
 wire n_8262;
 wire n_8263;
 wire n_8264;
 wire n_8265;
 wire n_8266;
 wire n_8267;
 wire n_8268;
 wire n_8269;
 wire n_827;
 wire n_8270;
 wire n_8271;
 wire n_8272;
 wire n_8273;
 wire n_8274;
 wire n_8275;
 wire n_8276;
 wire n_8277;
 wire n_8278;
 wire n_8279;
 wire n_828;
 wire n_8280;
 wire n_8281;
 wire n_8282;
 wire n_8283;
 wire n_8284;
 wire n_8285;
 wire n_8286;
 wire n_8287;
 wire n_8289;
 wire n_829;
 wire n_8290;
 wire n_8291;
 wire n_8293;
 wire n_8294;
 wire n_8295;
 wire n_8296;
 wire n_8298;
 wire n_8299;
 wire n_83;
 wire n_830;
 wire n_8300;
 wire n_8301;
 wire n_8302;
 wire n_8303;
 wire n_8304;
 wire n_8305;
 wire n_8307;
 wire n_8308;
 wire n_8309;
 wire n_831;
 wire n_8310;
 wire n_8311;
 wire n_8312;
 wire n_8313;
 wire n_8314;
 wire n_8315;
 wire n_8316;
 wire n_8317;
 wire n_8318;
 wire n_8319;
 wire n_832;
 wire n_8320;
 wire n_8321;
 wire n_8322;
 wire n_8323;
 wire n_8324;
 wire n_8325;
 wire n_8326;
 wire n_8327;
 wire n_8328;
 wire n_8329;
 wire n_833;
 wire n_8330;
 wire n_8331;
 wire n_8332;
 wire n_8333;
 wire n_8334;
 wire n_8335;
 wire n_8336;
 wire n_8337;
 wire n_8338;
 wire n_8339;
 wire n_834;
 wire n_8340;
 wire n_8342;
 wire n_8343;
 wire n_8344;
 wire n_8345;
 wire n_8346;
 wire n_835;
 wire n_836;
 wire n_837;
 wire n_838;
 wire n_839;
 wire n_84;
 wire n_840;
 wire n_841;
 wire n_842;
 wire n_843;
 wire n_844;
 wire n_845;
 wire n_846;
 wire n_847;
 wire n_848;
 wire n_849;
 wire n_85;
 wire n_850;
 wire n_851;
 wire n_852;
 wire n_853;
 wire n_854;
 wire n_855;
 wire n_856;
 wire n_857;
 wire n_858;
 wire n_859;
 wire n_86;
 wire n_860;
 wire n_861;
 wire n_862;
 wire n_8623;
 wire n_8625;
 wire n_8629;
 wire n_863;
 wire n_864;
 wire n_865;
 wire n_8652;
 wire n_8656;
 wire n_866;
 wire n_8668;
 wire n_867;
 wire n_8678;
 wire n_8679;
 wire n_868;
 wire n_8687;
 wire n_8688;
 wire n_869;
 wire n_8690;
 wire n_8691;
 wire n_87;
 wire n_870;
 wire n_8702;
 wire n_8703;
 wire n_871;
 wire n_8719;
 wire n_872;
 wire n_8720;
 wire n_8723;
 wire n_873;
 wire n_8732;
 wire n_8733;
 wire n_8738;
 wire n_874;
 wire n_8742;
 wire n_8747;
 wire n_8748;
 wire n_875;
 wire n_876;
 wire n_8760;
 wire n_8766;
 wire n_877;
 wire n_8770;
 wire n_8771;
 wire n_8779;
 wire n_878;
 wire n_8780;
 wire n_8783;
 wire n_8785;
 wire n_8789;
 wire n_879;
 wire n_8792;
 wire n_88;
 wire n_880;
 wire n_8801;
 wire n_881;
 wire n_882;
 wire n_8820;
 wire n_883;
 wire n_8831;
 wire n_8833;
 wire n_884;
 wire n_8847;
 wire n_885;
 wire n_8851;
 wire n_8856;
 wire n_886;
 wire n_887;
 wire n_8872;
 wire n_8877;
 wire n_8879;
 wire n_888;
 wire n_8881;
 wire n_8884;
 wire n_8887;
 wire n_889;
 wire n_8894;
 wire n_8896;
 wire n_8899;
 wire n_89;
 wire n_890;
 wire n_8908;
 wire n_891;
 wire n_8912;
 wire n_892;
 wire n_8922;
 wire n_8923;
 wire n_893;
 wire n_8932;
 wire n_8933;
 wire n_894;
 wire n_8942;
 wire n_8946;
 wire n_895;
 wire n_896;
 wire n_8963;
 wire n_8964;
 wire n_897;
 wire n_898;
 wire n_899;
 wire n_8992;
 wire n_8993;
 wire n_8994;
 wire n_8995;
 wire n_8996;
 wire n_8997;
 wire n_8998;
 wire n_8999;
 wire n_9;
 wire n_90;
 wire n_900;
 wire n_9000;
 wire n_9001;
 wire n_9002;
 wire n_9005;
 wire n_9008;
 wire n_901;
 wire n_9011;
 wire n_9014;
 wire n_9017;
 wire n_902;
 wire n_9020;
 wire n_9023;
 wire n_9026;
 wire n_9029;
 wire n_903;
 wire n_9032;
 wire n_9035;
 wire n_9038;
 wire n_904;
 wire n_9041;
 wire n_9044;
 wire n_9047;
 wire n_905;
 wire n_9050;
 wire n_9053;
 wire n_9056;
 wire n_9059;
 wire n_906;
 wire n_9062;
 wire n_9065;
 wire n_9068;
 wire n_907;
 wire n_9071;
 wire n_9074;
 wire n_9077;
 wire n_908;
 wire n_9080;
 wire n_9083;
 wire n_9086;
 wire n_9089;
 wire n_909;
 wire n_9092;
 wire n_9095;
 wire n_9098;
 wire n_91;
 wire n_910;
 wire n_9101;
 wire n_9104;
 wire n_9107;
 wire n_911;
 wire n_9110;
 wire n_9113;
 wire n_9116;
 wire n_9119;
 wire n_912;
 wire n_9122;
 wire n_9125;
 wire n_9128;
 wire n_913;
 wire n_9131;
 wire n_9134;
 wire n_9137;
 wire n_914;
 wire n_9140;
 wire n_9143;
 wire n_9146;
 wire n_9149;
 wire n_915;
 wire n_9152;
 wire n_9155;
 wire n_9158;
 wire n_916;
 wire n_9161;
 wire n_9164;
 wire n_9167;
 wire n_917;
 wire n_9170;
 wire n_9173;
 wire n_9176;
 wire n_9179;
 wire n_918;
 wire n_9182;
 wire n_9185;
 wire n_9188;
 wire n_919;
 wire n_9191;
 wire n_9194;
 wire n_9197;
 wire n_92;
 wire n_920;
 wire n_9200;
 wire n_9203;
 wire n_9206;
 wire n_9209;
 wire n_921;
 wire n_9212;
 wire n_9215;
 wire n_9218;
 wire n_922;
 wire n_9221;
 wire n_9224;
 wire n_9227;
 wire n_923;
 wire n_9230;
 wire n_9233;
 wire n_9236;
 wire n_9239;
 wire n_924;
 wire n_9242;
 wire n_9245;
 wire n_9248;
 wire n_925;
 wire n_9251;
 wire n_9254;
 wire n_9257;
 wire n_926;
 wire n_9260;
 wire n_9263;
 wire n_9266;
 wire n_9269;
 wire n_927;
 wire n_9272;
 wire n_9275;
 wire n_9278;
 wire n_928;
 wire n_9281;
 wire n_9284;
 wire n_9287;
 wire n_929;
 wire n_9290;
 wire n_9293;
 wire n_9296;
 wire n_9299;
 wire n_93;
 wire n_930;
 wire n_9302;
 wire n_9305;
 wire n_9308;
 wire n_931;
 wire n_9311;
 wire n_9314;
 wire n_9317;
 wire n_932;
 wire n_9320;
 wire n_9323;
 wire n_9326;
 wire n_9329;
 wire n_933;
 wire n_9332;
 wire n_9335;
 wire n_9338;
 wire n_934;
 wire n_9341;
 wire n_9344;
 wire n_9347;
 wire n_935;
 wire n_9350;
 wire n_9353;
 wire n_9356;
 wire n_9359;
 wire n_936;
 wire n_9362;
 wire n_9365;
 wire n_9368;
 wire n_937;
 wire n_9371;
 wire n_9374;
 wire n_9377;
 wire n_938;
 wire n_9380;
 wire n_9383;
 wire n_9386;
 wire n_939;
 wire n_9393;
 wire n_9398;
 wire n_94;
 wire n_940;
 wire n_9403;
 wire n_9408;
 wire n_941;
 wire n_9413;
 wire n_9418;
 wire n_942;
 wire n_9423;
 wire n_9428;
 wire n_943;
 wire n_9433;
 wire n_9438;
 wire n_944;
 wire n_9443;
 wire n_9448;
 wire n_945;
 wire n_9453;
 wire n_9458;
 wire n_946;
 wire n_9463;
 wire n_9468;
 wire n_947;
 wire n_9473;
 wire n_9478;
 wire n_948;
 wire n_9483;
 wire n_9488;
 wire n_9493;
 wire n_9498;
 wire n_95;
 wire n_950;
 wire n_9503;
 wire n_9508;
 wire n_951;
 wire n_9513;
 wire n_9518;
 wire n_952;
 wire n_9523;
 wire n_9528;
 wire n_953;
 wire n_9533;
 wire n_9538;
 wire n_954;
 wire n_9543;
 wire n_9548;
 wire n_955;
 wire n_9553;
 wire n_9558;
 wire n_956;
 wire n_9563;
 wire n_9568;
 wire n_9573;
 wire n_9578;
 wire n_958;
 wire n_9583;
 wire n_9588;
 wire n_959;
 wire n_9593;
 wire n_9598;
 wire n_96;
 wire n_960;
 wire n_9603;
 wire n_9608;
 wire n_961;
 wire n_9613;
 wire n_9618;
 wire n_962;
 wire n_9623;
 wire n_9628;
 wire n_963;
 wire n_9633;
 wire n_9638;
 wire n_964;
 wire n_9643;
 wire n_9648;
 wire n_965;
 wire n_9653;
 wire n_9658;
 wire n_9663;
 wire n_9668;
 wire n_967;
 wire n_9673;
 wire n_9678;
 wire n_968;
 wire n_9683;
 wire n_9688;
 wire n_969;
 wire n_9693;
 wire n_9698;
 wire n_97;
 wire n_970;
 wire n_9703;
 wire n_9708;
 wire n_971;
 wire n_9713;
 wire n_9718;
 wire n_972;
 wire n_9723;
 wire n_9728;
 wire n_973;
 wire n_9733;
 wire n_9738;
 wire n_974;
 wire n_9743;
 wire n_9748;
 wire n_975;
 wire n_9753;
 wire n_9758;
 wire n_976;
 wire n_9763;
 wire n_9768;
 wire n_977;
 wire n_9773;
 wire n_9778;
 wire n_978;
 wire n_9783;
 wire n_9788;
 wire n_979;
 wire n_9793;
 wire n_9798;
 wire n_98;
 wire n_980;
 wire n_9803;
 wire n_9808;
 wire n_981;
 wire n_9813;
 wire n_9818;
 wire n_982;
 wire n_9823;
 wire n_9828;
 wire n_983;
 wire n_9833;
 wire n_9838;
 wire n_984;
 wire n_9843;
 wire n_9848;
 wire n_985;
 wire n_9853;
 wire n_9858;
 wire n_986;
 wire n_9863;
 wire n_9868;
 wire n_987;
 wire n_9873;
 wire n_9878;
 wire n_988;
 wire n_9883;
 wire n_9888;
 wire n_989;
 wire n_9893;
 wire n_9898;
 wire n_99;
 wire n_990;
 wire n_9903;
 wire n_9908;
 wire n_991;
 wire n_9913;
 wire n_9918;
 wire n_992;
 wire n_9923;
 wire n_9928;
 wire n_993;
 wire n_9933;
 wire n_9938;
 wire n_994;
 wire n_9943;
 wire n_9948;
 wire n_995;
 wire n_9953;
 wire n_9958;
 wire n_996;
 wire n_9963;
 wire n_9968;
 wire n_997;
 wire n_9973;
 wire n_9978;
 wire n_998;
 wire n_9983;
 wire n_9988;
 wire n_999;
 wire n_9993;
 wire n_9998;
 wire \text_out[0]_3160 ;
 wire \text_out[100]_3140 ;
 wire \text_out[101]_3141 ;
 wire \text_out[102]_3142 ;
 wire \text_out[103]_3143 ;
 wire \text_out[104]_3104 ;
 wire \text_out[105]_3105 ;
 wire \text_out[106]_3106 ;
 wire \text_out[107]_3107 ;
 wire \text_out[108]_3108 ;
 wire \text_out[109]_3109 ;
 wire \text_out[10]_3130 ;
 wire \text_out[110]_3110 ;
 wire \text_out[111]_3111 ;
 wire \text_out[112]_3072 ;
 wire \text_out[113]_3073 ;
 wire \text_out[114]_3074 ;
 wire \text_out[115]_3075 ;
 wire \text_out[116]_3076 ;
 wire \text_out[117]_3077 ;
 wire \text_out[118]_3078 ;
 wire \text_out[119]_3079 ;
 wire \text_out[11]_3131 ;
 wire \text_out[120]_3040 ;
 wire \text_out[121]_3041 ;
 wire \text_out[122]_3042 ;
 wire \text_out[123]_3043 ;
 wire \text_out[124]_3044 ;
 wire \text_out[125]_3045 ;
 wire \text_out[126]_3046 ;
 wire \text_out[127]_3047 ;
 wire \text_out[12]_3132 ;
 wire \text_out[13]_3133 ;
 wire \text_out[14]_3134 ;
 wire \text_out[15]_3135 ;
 wire \text_out[16]_3096 ;
 wire \text_out[17]_3097 ;
 wire \text_out[18]_3098 ;
 wire \text_out[19]_3099 ;
 wire \text_out[1]_3161 ;
 wire \text_out[20]_3100 ;
 wire \text_out[21]_3101 ;
 wire \text_out[22]_3102 ;
 wire \text_out[23]_3103 ;
 wire \text_out[24]_3064 ;
 wire \text_out[25]_3065 ;
 wire \text_out[26]_3066 ;
 wire \text_out[27]_3067 ;
 wire \text_out[28]_3068 ;
 wire \text_out[29]_3069 ;
 wire \text_out[2]_3162 ;
 wire \text_out[30]_3070 ;
 wire \text_out[31]_3071 ;
 wire \text_out[32]_3152 ;
 wire \text_out[33]_3153 ;
 wire \text_out[34]_3154 ;
 wire \text_out[35]_3155 ;
 wire \text_out[36]_3156 ;
 wire \text_out[37]_3157 ;
 wire \text_out[38]_3158 ;
 wire \text_out[39]_3159 ;
 wire \text_out[3]_3163 ;
 wire \text_out[40]_3120 ;
 wire \text_out[41]_3121 ;
 wire \text_out[42]_3122 ;
 wire \text_out[43]_3123 ;
 wire \text_out[44]_3124 ;
 wire \text_out[45]_3125 ;
 wire \text_out[46]_3126 ;
 wire \text_out[47]_3127 ;
 wire \text_out[48]_3088 ;
 wire \text_out[49]_3089 ;
 wire \text_out[4]_3164 ;
 wire \text_out[50]_3090 ;
 wire \text_out[51]_3091 ;
 wire \text_out[52]_3092 ;
 wire \text_out[53]_3093 ;
 wire \text_out[54]_3094 ;
 wire \text_out[55]_3095 ;
 wire \text_out[56]_3056 ;
 wire \text_out[57]_3057 ;
 wire \text_out[58]_3058 ;
 wire \text_out[59]_3059 ;
 wire \text_out[5]_3165 ;
 wire \text_out[60]_3060 ;
 wire \text_out[61]_3061 ;
 wire \text_out[62]_3062 ;
 wire \text_out[63]_3063 ;
 wire \text_out[64]_3144 ;
 wire \text_out[65]_3145 ;
 wire \text_out[66]_3146 ;
 wire \text_out[67]_3147 ;
 wire \text_out[68]_3148 ;
 wire \text_out[69]_3149 ;
 wire \text_out[6]_3166 ;
 wire \text_out[70]_3150 ;
 wire \text_out[71]_3151 ;
 wire \text_out[72]_3112 ;
 wire \text_out[73]_3113 ;
 wire \text_out[74]_3114 ;
 wire \text_out[75]_3115 ;
 wire \text_out[76]_3116 ;
 wire \text_out[77]_3117 ;
 wire \text_out[78]_3118 ;
 wire \text_out[79]_3119 ;
 wire \text_out[7]_3167 ;
 wire \text_out[80]_3080 ;
 wire \text_out[81]_3081 ;
 wire \text_out[82]_3082 ;
 wire \text_out[83]_3083 ;
 wire \text_out[84]_3084 ;
 wire \text_out[85]_3085 ;
 wire \text_out[86]_3086 ;
 wire \text_out[87]_3087 ;
 wire \text_out[88]_3048 ;
 wire \text_out[89]_3049 ;
 wire \text_out[8]_3128 ;
 wire \text_out[90]_3050 ;
 wire \text_out[91]_3051 ;
 wire \text_out[92]_3052 ;
 wire \text_out[93]_3053 ;
 wire \text_out[94]_3054 ;
 wire \text_out[95]_3055 ;
 wire \text_out[96]_3136 ;
 wire \text_out[97]_3137 ;
 wire \text_out[98]_3138 ;
 wire \text_out[99]_3139 ;
 wire \text_out[9]_3129 ;
 wire u0_n_29279;
 wire u0_n_29280;
 wire u0_n_29281;
 wire u0_n_29283;
 wire u0_n_29284;
 wire u0_n_29285;
 wire u0_n_29286;
 wire u0_n_29287;
 wire u0_n_29288;
 wire u0_n_29289;
 wire u0_n_29290;
 wire u0_n_29291;
 wire u0_n_29292;
 wire u0_n_29293;
 wire u0_n_29294;
 wire u0_n_29295;
 wire u0_n_29296;
 wire u0_n_29297;
 wire u0_n_29298;
 wire u0_n_29299;
 wire u0_n_29300;
 wire u0_n_29301;
 wire u0_n_29302;
 wire u0_n_29303;
 wire u0_n_29305;
 wire u0_n_29308;
 wire u0_n_29311;
 wire u0_n_29314;
 wire u0_n_29317;
 wire u0_n_29320;
 wire u0_n_29321;
 wire u0_n_29322;
 wire u0_n_29324;
 wire u0_n_29326;
 wire u0_n_29328;
 wire u0_n_29329;
 wire u0_n_29330;
 wire u0_n_29331;
 wire u0_n_29332;
 wire u0_n_29334;
 wire u0_n_29335;
 wire u0_n_29336;
 wire u0_n_29337;
 wire u0_n_29338;
 wire u0_n_29339;
 wire u0_n_29341;
 wire u0_n_29342;
 wire u0_n_29343;
 wire u0_n_29344;
 wire u0_n_29345;
 wire u0_n_29348;
 wire u0_n_29350;
 wire u0_n_29353;
 wire u0_n_29355;
 wire u0_n_29356;
 wire u0_n_29357;
 wire u0_n_29360;
 wire u0_n_29363;
 wire u0_n_29364;
 wire u0_n_29368;
 wire u0_n_29369;
 wire u0_n_29371;
 wire u0_n_29372;
 wire u0_n_29373;
 wire u0_n_29374;
 wire u0_n_29375;
 wire u0_n_29376;
 wire u0_n_29377;
 wire u0_n_29378;
 wire u0_n_29379;
 wire u0_n_29380;
 wire u0_n_29381;
 wire u0_n_29382;
 wire u0_n_29383;
 wire u0_n_29384;
 wire u0_n_29385;
 wire u0_n_29386;
 wire u0_n_29387;
 wire u0_n_29388;
 wire u0_n_29390;
 wire u0_n_29391;
 wire u0_n_29392;
 wire u0_n_29393;
 wire u0_n_29394;
 wire u0_n_29395;
 wire u0_n_29396;
 wire u0_n_29397;
 wire u0_n_29398;
 wire u0_n_29399;
 wire u0_n_29400;
 wire u0_n_29402;
 wire u0_n_29403;
 wire u0_n_29404;
 wire u0_n_29406;
 wire u0_n_29407;
 wire u0_n_29408;
 wire u0_n_29409;
 wire u0_n_29410;
 wire u0_n_29411;
 wire u0_n_29414;
 wire u0_n_29417;
 wire u0_n_29418;
 wire u0_n_29421;
 wire u0_n_29424;
 wire u0_n_29426;
 wire u0_n_29429;
 wire u0_n_29431;
 wire u0_n_29432;
 wire u0_n_29434;
 wire u0_n_29435;
 wire u0_n_29436;
 wire u0_n_29440;
 wire u0_n_29441;
 wire u0_n_29444;
 wire u0_n_29459;
 wire u0_n_29460;
 wire u0_n_29461;
 wire u0_n_29462;
 wire u0_n_29463;
 wire u0_n_29465;
 wire u0_n_29467;
 wire u0_n_29468;
 wire u0_n_29469;
 wire u0_n_29470;
 wire u0_n_29471;
 wire u0_n_29472;
 wire u0_n_29473;
 wire u0_n_29474;
 wire u0_n_29475;
 wire u0_n_29476;
 wire u0_n_29477;
 wire u0_n_29478;
 wire u0_n_29479;
 wire u0_n_29480;
 wire u0_n_29481;
 wire u0_n_29482;
 wire u0_n_29483;
 wire u0_n_29484;
 wire u0_n_29485;
 wire u0_n_29486;
 wire u0_n_29487;
 wire u0_n_29488;
 wire u0_n_29489;
 wire u0_n_29490;
 wire u0_n_29491;
 wire u0_n_29492;
 wire u0_n_29493;
 wire u0_n_29494;
 wire u0_n_29496;
 wire u0_n_29498;
 wire u0_n_29500;
 wire u0_n_29503;
 wire u0_n_29506;
 wire u0_n_29520;
 wire u0_n_29521;
 wire u0_n_29522;
 wire u0_n_29523;
 wire u0_n_29524;
 wire u0_n_29526;
 wire u0_n_29527;
 wire u0_n_29528;
 wire u0_n_29529;
 wire u0_n_29530;
 wire u0_n_29531;
 wire u0_n_29532;
 wire u0_n_29533;
 wire u0_n_29534;
 wire u0_n_29535;
 wire u0_n_29536;
 wire u0_n_29537;
 wire u0_n_29538;
 wire u0_n_29539;
 wire u0_n_29540;
 wire u0_n_29541;
 wire u0_n_29542;
 wire u0_n_29543;
 wire u0_n_29544;
 wire u0_n_29547;
 wire u0_n_29548;
 wire u0_n_29549;
 wire u0_n_29550;
 wire u0_n_29551;
 wire u0_n_29552;
 wire u0_n_29553;
 wire u0_n_29554;
 wire u0_n_29555;
 wire u0_n_29556;
 wire u0_n_29557;
 wire u0_n_29558;
 wire u0_n_29559;
 wire u0_n_29560;
 wire u0_n_29561;
 wire u0_n_29562;
 wire u0_n_29563;
 wire u0_n_29564;
 wire u0_n_29565;
 wire u0_n_29566;
 wire u0_n_29567;
 wire u0_n_29568;
 wire u0_n_29569;
 wire u0_n_29570;
 wire u0_n_29571;
 wire u0_n_29574;
 wire u0_n_29579;
 wire u0_n_29582;
 wire u0_n_29584;
 wire u0_n_29587;
 wire u0_n_29590;
 wire u0_n_29616;
 wire u0_n_29617;
 wire u0_n_29618;
 wire u0_n_29619;
 wire u0_n_29620;
 wire u0_n_29621;
 wire u0_n_29623;
 wire u0_n_29624;
 wire u0_n_29625;
 wire u0_n_29627;
 wire u0_n_29632;
 wire u0_n_29633;
 wire u0_n_29634;
 wire u0_n_29635;
 wire u0_n_29636;
 wire u0_n_29637;
 wire u0_n_29638;
 wire u0_n_29639;
 wire u0_n_29640;
 wire u0_n_29641;
 wire u0_n_29642;
 wire u0_n_29643;
 wire u0_n_29646;
 wire u0_n_29649;
 wire u0_n_29657;
 wire u0_n_29658;
 wire u0_n_29659;
 wire u0_n_29660;
 wire u0_n_29661;
 wire u0_n_29662;
 wire u0_n_29663;
 wire u0_n_29664;
 wire u0_n_29665;
 wire u0_n_29666;
 wire u0_n_29667;
 wire u0_n_29668;
 wire u0_n_29669;
 wire u0_n_29676;
 wire u0_n_29677;
 wire u0_n_29678;
 wire u0_n_29679;
 wire u0_n_29680;
 wire u0_n_29681;
 wire u0_n_29682;
 wire u0_n_29683;
 wire u0_n_29684;
 wire u0_n_29687;
 wire u0_n_29688;
 wire u0_n_29690;
 wire u0_n_29700;
 wire u0_n_29701;
 wire u0_n_29702;
 wire u0_n_29703;
 wire u0_n_29704;
 wire u0_n_29706;
 wire u0_n_29708;
 wire u0_n_29709;
 wire u0_n_29710;
 wire u0_n_29711;
 wire u0_n_29712;
 wire u0_n_29714;
 wire u0_n_29717;
 wire u0_n_29718;
 wire u0_n_29719;
 wire u0_n_29720;
 wire u0_n_29721;
 wire u0_n_29722;
 wire u0_n_29723;
 wire u0_n_29724;
 wire u0_n_29725;
 wire u0_n_29726;
 wire u0_n_29727;
 wire u0_n_29728;
 wire u0_n_29729;
 wire u0_n_29730;
 wire u0_n_29731;
 wire u0_n_29733;
 wire u0_n_29734;
 wire u0_n_29735;
 wire u0_n_29736;
 wire u0_n_29738;
 wire u0_n_29739;
 wire u0_n_29742;
 wire u0_n_29744;
 wire u0_n_29745;
 wire u0_n_29746;
 wire u0_n_29747;
 wire u0_n_29748;
 wire u0_n_29750;
 wire u0_n_29751;
 wire u0_n_29752;
 wire u0_n_29753;
 wire u0_n_29754;
 wire u0_n_29755;
 wire u0_n_29756;
 wire u0_n_29757;
 wire u0_n_29759;
 wire u0_n_29761;
 wire u0_n_29763;
 wire u0_n_29765;
 wire u0_n_29767;
 wire u0_n_29770;
 wire u0_n_29772;
 wire u0_n_29773;
 wire u0_n_29774;
 wire u0_n_29775;
 wire u0_n_29776;
 wire u0_n_29777;
 wire u0_n_29778;
 wire u0_n_29780;
 wire u0_n_29781;
 wire u0_n_29782;
 wire u0_n_29783;
 wire u0_n_29785;
 wire u0_n_29786;
 wire u0_n_29787;
 wire u0_n_29789;
 wire u0_n_29790;
 wire u0_n_29791;
 wire u0_n_29794;
 wire u0_n_29795;
 wire u0_n_29796;
 wire u0_n_29797;
 wire u0_n_29798;
 wire u0_n_29800;
 wire u0_n_29801;
 wire u0_n_29802;
 wire u0_n_29804;
 wire u0_n_29806;
 wire u0_n_29807;
 wire u0_n_29808;
 wire u0_n_29810;
 wire u0_n_29811;
 wire u0_n_29813;
 wire u0_n_29815;
 wire u0_n_29817;
 wire u0_n_29818;
 wire u0_n_29819;
 wire u0_n_29821;
 wire u0_n_29822;
 wire u0_n_29824;
 wire u0_n_29825;
 wire u0_n_29826;
 wire u0_n_29828;
 wire u0_n_29831;
 wire u0_n_29832;
 wire u0_n_29833;
 wire u0_n_29835;
 wire u0_n_29837;
 wire u0_n_29838;
 wire u0_n_29840;
 wire u0_n_29842;
 wire u0_n_29844;
 wire u0_n_29845;
 wire u0_n_29846;
 wire u0_n_29848;
 wire u0_n_29850;
 wire u0_n_29852;
 wire u0_n_29853;
 wire u0_n_29855;
 wire u0_n_29857;
 wire u0_n_29859;
 wire u0_n_29861;
 wire u0_n_29863;
 wire u0_n_29864;
 wire u0_n_29866;
 wire u0_n_29868;
 wire u0_n_29869;
 wire u0_n_29870;
 wire u0_n_29871;
 wire u0_n_29872;
 wire u0_n_29874;
 wire u0_n_29877;
 wire u0_n_29878;
 wire u0_n_29881;
 wire u0_n_29883;
 wire u0_n_29886;
 wire u0_n_29887;
 wire u0_n_29889;
 wire u0_n_29890;
 wire u0_n_29891;
 wire u0_n_29892;
 wire u0_n_29894;
 wire u0_n_29896;
 wire u0_n_29898;
 wire u0_n_29900;
 wire u0_n_29901;
 wire u0_n_29903;
 wire u0_n_29904;
 wire u0_n_29908;
 wire u0_n_29909;
 wire u0_n_29910;
 wire u0_n_29911;
 wire u0_n_29912;
 wire u0_n_29913;
 wire u0_n_29916;
 wire u0_n_29919;
 wire u0_n_29922;
 wire u0_n_29923;
 wire u0_n_29924;
 wire u0_n_29926;
 wire u0_n_29928;
 wire u0_n_29929;
 wire u0_n_29930;
 wire u0_n_29931;
 wire u0_n_29932;
 wire u0_n_29933;
 wire u0_n_29934;
 wire u0_n_29935;
 wire u0_n_29936;
 wire u0_n_29937;
 wire u0_n_29938;
 wire u0_n_29940;
 wire u0_n_29941;
 wire u0_n_29944;
 wire u0_n_29946;
 wire u0_n_29948;
 wire u0_n_29950;
 wire u0_n_29951;
 wire u0_n_29952;
 wire u0_n_29957;
 wire u0_n_29958;
 wire u0_n_29959;
 wire u0_n_29960;
 wire u0_n_29962;
 wire u0_n_29963;
 wire u0_n_29964;
 wire u0_n_29966;
 wire u0_n_29968;
 wire u0_n_29969;
 wire u0_n_29970;
 wire u0_n_29971;
 wire u0_n_29972;
 wire u0_n_29973;
 wire u0_n_29975;
 wire u0_n_29976;
 wire u0_n_29978;
 wire u0_n_29980;
 wire u0_n_29981;
 wire u0_n_29983;
 wire u0_n_29984;
 wire u0_n_29986;
 wire u0_n_29987;
 wire u0_n_29988;
 wire u0_n_29989;
 wire u0_n_29990;
 wire u0_n_29991;
 wire u0_n_29992;
 wire u0_n_29994;
 wire u0_n_29997;
 wire u0_n_29999;
 wire u0_n_30001;
 wire u0_n_30003;
 wire u0_n_30004;
 wire u0_n_30006;
 wire u0_n_30008;
 wire u0_n_30009;
 wire u0_n_30011;
 wire u0_n_30013;
 wire u0_n_30014;
 wire u0_n_30016;
 wire u0_n_30017;
 wire u0_n_30018;
 wire u0_n_30020;
 wire u0_n_30021;
 wire u0_n_30022;
 wire u0_n_30024;
 wire u0_n_30027;
 wire u0_n_30028;
 wire u0_n_30029;
 wire u0_n_30031;
 wire u0_n_30032;
 wire u0_n_30033;
 wire u0_n_30035;
 wire u0_n_30037;
 wire u0_n_30039;
 wire u0_n_30041;
 wire u0_n_30043;
 wire u0_n_30044;
 wire u0_n_30046;
 wire u0_n_30047;
 wire u0_n_30049;
 wire u0_n_30051;
 wire u0_n_30052;
 wire u0_n_30054;
 wire u0_n_30056;
 wire u0_n_30058;
 wire u0_n_30059;
 wire u0_n_30062;
 wire u0_n_30064;
 wire u0_n_30066;
 wire u0_n_30068;
 wire u0_n_30070;
 wire u0_n_30072;
 wire u0_n_30076;
 wire u0_n_30078;
 wire u0_n_30080;
 wire u0_n_30081;
 wire u0_n_30082;
 wire u0_n_30083;
 wire u0_n_30087;
 wire u0_n_30090;
 wire u0_n_30092;
 wire u0_n_30094;
 wire u0_n_30096;
 wire u0_n_30098;
 wire u0_n_30099;
 wire u0_n_30101;
 wire u0_n_30102;
 wire u0_n_30104;
 wire u0_n_30105;
 wire u0_n_30108;
 wire u0_n_30109;
 wire u0_n_30111;
 wire u0_n_30114;
 wire u0_n_30115;
 wire u0_n_30119;
 wire u0_n_30120;
 wire u0_n_30121;
 wire u0_n_30122;
 wire u0_n_30123;
 wire u0_n_30124;
 wire u0_n_30126;
 wire u0_n_30128;
 wire u0_n_30129;
 wire u0_n_30131;
 wire u0_n_30132;
 wire u0_n_30133;
 wire u0_n_30134;
 wire u0_n_30136;
 wire u0_n_30137;
 wire u0_n_30138;
 wire u0_n_30140;
 wire u0_n_30141;
 wire u0_n_30144;
 wire u0_n_30146;
 wire u0_n_30148;
 wire u0_n_30150;
 wire u0_n_30153;
 wire u0_n_30155;
 wire u0_n_30156;
 wire u0_n_30158;
 wire u0_n_30159;
 wire u0_n_30160;
 wire u0_n_30161;
 wire u0_n_30163;
 wire u0_n_30165;
 wire u0_n_30166;
 wire u0_n_30168;
 wire u0_n_30169;
 wire u0_n_30170;
 wire u0_n_30172;
 wire u0_n_30176;
 wire u0_n_30178;
 wire u0_n_30180;
 wire u0_n_30182;
 wire u0_n_30183;
 wire u0_n_30185;
 wire u0_n_30187;
 wire u0_n_30189;
 wire u0_n_30190;
 wire u0_n_30191;
 wire u0_n_30192;
 wire u0_n_30193;
 wire u0_n_30194;
 wire u0_n_30195;
 wire u0_n_30196;
 wire u0_n_30197;
 wire u0_n_30198;
 wire u0_n_30199;
 wire u0_n_30200;
 wire u0_n_30201;
 wire u0_n_30204;
 wire u0_n_30207;
 wire u0_n_30209;
 wire u0_n_30211;
 wire u0_n_30214;
 wire u0_n_30215;
 wire u0_n_30217;
 wire u0_n_30218;
 wire u0_n_30221;
 wire u0_n_30223;
 wire u0_n_30224;
 wire u0_n_30229;
 wire u0_n_30232;
 wire u0_n_30233;
 wire u0_n_30235;
 wire u0_n_30237;
 wire u0_n_30240;
 wire u0_n_30242;
 wire u0_n_30244;
 wire u0_n_30247;
 wire u0_n_30249;
 wire u0_n_30250;
 wire u0_n_30252;
 wire u0_n_30255;
 wire u0_n_30257;
 wire u0_n_30258;
 wire u0_n_30261;
 wire u0_n_30263;
 wire u0_n_30266;
 wire u0_n_30267;
 wire u0_n_30268;
 wire u0_n_30269;
 wire u0_n_30270;
 wire u0_n_30271;
 wire u0_n_30273;
 wire u0_n_30274;
 wire u0_n_30276;
 wire u0_n_30277;
 wire u0_n_30279;
 wire u0_n_30280;
 wire u0_n_30283;
 wire u0_n_30284;
 wire u0_n_30286;
 wire u0_n_30289;
 wire u0_n_30290;
 wire u0_n_30292;
 wire u0_n_30293;
 wire u0_n_30296;
 wire u0_n_30298;
 wire u0_n_30299;
 wire u0_n_30302;
 wire u0_n_30304;
 wire u0_n_30309;
 wire u0_n_30310;
 wire u0_n_30314;
 wire u0_n_30317;
 wire u0_n_30321;
 wire u0_n_30323;
 wire u0_n_30324;
 wire u0_n_30326;
 wire u0_n_30330;
 wire u0_n_30332;
 wire u0_n_30334;
 wire u0_n_30337;
 wire u0_n_30339;
 wire u0_n_30341;
 wire u0_n_30343;
 wire u0_n_30346;
 wire u0_n_30348;
 wire u0_n_30349;
 wire u0_n_30350;
 wire u0_n_30351;
 wire u0_n_30352;
 wire u0_n_30353;
 wire u0_n_30354;
 wire u0_n_30355;
 wire u0_n_30356;
 wire u0_n_30357;
 wire u0_n_30358;
 wire u0_n_30359;
 wire u0_n_30360;
 wire u0_n_30361;
 wire u0_n_30362;
 wire u0_n_30363;
 wire u0_n_30364;
 wire u0_n_30365;
 wire u0_n_30366;
 wire u0_n_30367;
 wire u0_n_30368;
 wire u0_n_30369;
 wire u0_n_30370;
 wire u0_n_30371;
 wire u0_n_30372;
 wire u0_n_30373;
 wire u0_n_30375;
 wire u0_n_30377;
 wire u0_n_30380;
 wire u0_n_30382;
 wire u0_n_30383;
 wire u0_n_30385;
 wire u0_n_30388;
 wire u0_n_30390;
 wire u0_n_30391;
 wire u0_n_30392;
 wire u0_n_30395;
 wire u0_n_30396;
 wire u0_n_30398;
 wire u0_n_30400;
 wire u0_n_30402;
 wire u0_n_30404;
 wire u0_n_30405;
 wire u0_n_30406;
 wire u0_n_30408;
 wire u0_n_30409;
 wire u0_n_30411;
 wire u0_n_30413;
 wire u0_n_30415;
 wire u0_n_30418;
 wire u0_n_30419;
 wire u0_n_30420;
 wire u0_n_30422;
 wire u0_n_30423;
 wire u0_n_30425;
 wire u0_n_30427;
 wire u0_n_30428;
 wire u0_n_30431;
 wire u0_n_30435;
 wire u0_n_30438;
 wire u0_n_30441;
 wire u0_n_30443;
 wire u0_n_30445;
 wire u0_n_30449;
 wire u0_n_30450;
 wire u0_n_30452;
 wire u0_n_30453;
 wire u0_n_30454;
 wire u0_n_30457;
 wire u0_n_30459;
 wire u0_n_30460;
 wire u0_n_30461;
 wire u0_n_30463;
 wire u0_n_30464;
 wire u0_n_30465;
 wire u0_n_30467;
 wire u0_n_30469;
 wire u0_n_30471;
 wire u0_n_30472;
 wire u0_n_30474;
 wire u0_n_30476;
 wire u0_n_30477;
 wire u0_n_30478;
 wire u0_n_30480;
 wire u0_n_30482;
 wire u0_n_30484;
 wire u0_n_30486;
 wire u0_n_30488;
 wire u0_n_30489;
 wire u0_n_30491;
 wire u0_n_30492;
 wire u0_n_30493;
 wire u0_n_30495;
 wire u0_n_30498;
 wire u0_n_30501;
 wire u0_n_30503;
 wire u0_n_30504;
 wire u0_n_30506;
 wire u0_n_30514;
 wire u0_n_30520;
 wire u0_n_30521;
 wire u0_n_30522;
 wire u0_n_30524;
 wire u0_n_30525;
 wire u0_n_30527;
 wire u0_n_30529;
 wire u0_n_30530;
 wire u0_n_30531;
 wire u0_n_30532;
 wire u0_n_30535;
 wire u0_n_30536;
 wire u0_n_30538;
 wire u0_n_30540;
 wire u0_n_30541;
 wire u0_n_30542;
 wire u0_n_30543;
 wire u0_n_30544;
 wire u0_n_30546;
 wire u0_n_30549;
 wire u0_n_30550;
 wire u0_n_30551;
 wire u0_n_30553;
 wire u0_n_30555;
 wire u0_n_30557;
 wire u0_n_30558;
 wire u0_n_30560;
 wire u0_n_30561;
 wire u0_n_30563;
 wire u0_n_30565;
 wire u0_n_30567;
 wire u0_n_30569;
 wire u0_n_30570;
 wire u0_n_30572;
 wire u0_n_30573;
 wire u0_n_30575;
 wire u0_n_30576;
 wire u0_n_30577;
 wire u0_n_30578;
 wire u0_n_30582;
 wire u0_n_30584;
 wire u0_n_30586;
 wire u0_n_30589;
 wire u0_n_30591;
 wire u0_n_30592;
 wire u0_n_30594;
 wire u0_n_30595;
 wire u0_n_30597;
 wire u0_n_30598;
 wire u0_n_30599;
 wire u0_n_30602;
 wire u0_n_30605;
 wire u0_n_30606;
 wire u0_n_30608;
 wire u0_n_30611;
 wire u0_n_30614;
 wire u0_n_30615;
 wire u0_n_30618;
 wire u0_n_30623;
 wire u0_n_30626;
 wire u0_n_30629;
 wire u0_n_30632;
 wire u0_n_30635;
 wire u0_n_30640;
 wire u0_n_30644;
 wire u0_n_30647;
 wire u0_n_30648;
 wire u0_n_30650;
 wire u0_n_30652;
 wire u0_n_30653;
 wire u0_n_30654;
 wire u0_n_30658;
 wire u0_n_30659;
 wire u0_n_30663;
 wire u0_n_30667;
 wire u0_n_30668;
 wire u0_n_30670;
 wire u0_n_30672;
 wire u0_n_30674;
 wire u0_n_30676;
 wire u0_n_30679;
 wire u0_n_30680;
 wire u0_n_30683;
 wire u0_n_30685;
 wire u0_n_30686;
 wire u0_n_30688;
 wire u0_n_30690;
 wire u0_n_30692;
 wire u0_n_30695;
 wire u0_n_30697;
 wire u0_n_30698;
 wire u0_n_30700;
 wire u0_n_30702;
 wire u0_n_30704;
 wire u0_n_30705;
 wire u0_n_30708;
 wire u0_n_30711;
 wire u0_n_30715;
 wire u0_n_30717;
 wire u0_n_30718;
 wire u0_n_30719;
 wire u0_n_30720;
 wire u0_n_30721;
 wire u0_n_30722;
 wire u0_n_30723;
 wire u0_n_30724;
 wire u0_n_30725;
 wire u0_n_30726;
 wire u0_n_30727;
 wire u0_n_30728;
 wire u0_n_30729;
 wire u0_n_30730;
 wire u0_n_30731;
 wire u0_n_30732;
 wire u0_n_30733;
 wire u0_n_30734;
 wire u0_n_30735;
 wire u0_n_30736;
 wire u0_n_30737;
 wire u0_n_30738;
 wire u0_n_30739;
 wire u0_n_30740;
 wire u0_n_30741;
 wire u0_n_30742;
 wire u0_n_30743;
 wire u0_n_30744;
 wire u0_n_30745;
 wire u0_n_30746;
 wire u0_n_30747;
 wire u0_n_30748;
 wire u0_n_30749;
 wire u0_n_30750;
 wire u0_n_30751;
 wire u0_n_30752;
 wire u0_n_30753;
 wire u0_n_30754;
 wire u0_n_30755;
 wire u0_n_30756;
 wire u0_n_30757;
 wire u0_n_30758;
 wire u0_n_30759;
 wire u0_n_30760;
 wire u0_n_30761;
 wire u0_n_30762;
 wire u0_n_30763;
 wire u0_n_30764;
 wire u0_n_30765;
 wire u0_n_30766;
 wire u0_n_30767;
 wire u0_n_30768;
 wire u0_n_30769;
 wire u0_n_30770;
 wire u0_n_30771;
 wire u0_n_30772;
 wire u0_n_30773;
 wire u0_n_30774;
 wire u0_n_30775;
 wire u0_n_30776;
 wire u0_n_30777;
 wire u0_n_30778;
 wire u0_n_30779;
 wire u0_n_30782;
 wire u0_n_30784;
 wire u0_n_30785;
 wire u0_n_30786;
 wire u0_n_30788;
 wire u0_n_30789;
 wire u0_n_30791;
 wire u0_n_30793;
 wire u0_n_30796;
 wire u0_n_30798;
 wire u0_n_30799;
 wire u0_n_30802;
 wire u0_n_30804;
 wire u0_n_30806;
 wire u0_n_30808;
 wire u0_n_30810;
 wire u0_n_30811;
 wire u0_n_30814;
 wire u0_n_30817;
 wire u0_n_30820;
 wire u0_n_30822;
 wire u0_n_30824;
 wire u0_n_30825;
 wire u0_n_30826;
 wire u0_n_30828;
 wire u0_n_30831;
 wire u0_n_30833;
 wire u0_n_30835;
 wire u0_n_30837;
 wire u0_n_30840;
 wire u0_n_30843;
 wire u0_n_30845;
 wire u0_n_30847;
 wire u0_n_30849;
 wire u0_n_30851;
 wire u0_n_30853;
 wire u0_n_30854;
 wire u0_n_30857;
 wire u0_n_30858;
 wire u0_n_30859;
 wire u0_n_30861;
 wire u0_n_30864;
 wire u0_n_30867;
 wire u0_n_30868;
 wire u0_n_30869;
 wire u0_n_30871;
 wire u0_n_30872;
 wire u0_n_30873;
 wire u0_n_30875;
 wire u0_n_30876;
 wire u0_n_30890;
 wire u0_n_30899;
 wire u0_n_30900;
 wire u0_n_30901;
 wire u0_n_30902;
 wire u0_n_30903;
 wire u0_n_30904;
 wire u0_n_30905;
 wire u0_n_30906;
 wire u0_n_30907;
 wire u0_n_30908;
 wire u0_n_30909;
 wire u0_n_30910;
 wire u0_n_30911;
 wire u0_n_30912;
 wire u0_n_30913;
 wire u0_n_30914;
 wire u0_n_30915;
 wire u0_n_30918;
 wire u0_n_30921;
 wire u0_n_30922;
 wire u0_n_30926;
 wire u0_n_30928;
 wire u0_n_30931;
 wire u0_n_30932;
 wire u0_n_30934;
 wire u0_n_30935;
 wire u0_n_30936;
 wire u0_n_30938;
 wire u0_n_30941;
 wire u0_n_30943;
 wire u0_n_30946;
 wire u0_n_30949;
 wire u0_n_30950;
 wire u0_n_30952;
 wire u0_n_30953;
 wire u0_n_30956;
 wire u0_n_30958;
 wire u0_n_30959;
 wire u0_n_30960;
 wire u0_n_30961;
 wire u0_n_30963;
 wire u0_n_30964;
 wire u0_n_30967;
 wire u0_n_30969;
 wire u0_n_30971;
 wire u0_n_30972;
 wire u0_n_30975;
 wire u0_n_30976;
 wire u0_n_30977;
 wire u0_n_30978;
 wire u0_n_30980;
 wire u0_n_30983;
 wire u0_n_30985;
 wire u0_n_30986;
 wire u0_n_30987;
 wire u0_n_30988;
 wire u0_n_30990;
 wire u0_n_30992;
 wire u0_n_30994;
 wire u0_n_30996;
 wire u0_n_30997;
 wire u0_n_30998;
 wire u0_n_31000;
 wire u0_n_31001;
 wire u0_n_31002;
 wire u0_n_31004;
 wire u0_n_31005;
 wire u0_n_31006;
 wire u0_n_31009;
 wire u0_n_31011;
 wire u0_n_31012;
 wire u0_n_31014;
 wire u0_n_31016;
 wire u0_n_31017;
 wire u0_n_31019;
 wire u0_n_31021;
 wire u0_n_31023;
 wire u0_n_31026;
 wire u0_n_31027;
 wire u0_n_31028;
 wire u0_n_31030;
 wire u0_n_31033;
 wire u0_n_31036;
 wire u0_n_31038;
 wire u0_n_31040;
 wire u0_n_31041;
 wire u0_n_31043;
 wire u0_n_31045;
 wire u0_n_31048;
 wire u0_n_31050;
 wire u0_n_31051;
 wire u0_n_31053;
 wire u0_n_31054;
 wire u0_n_31055;
 wire u0_n_31056;
 wire u0_n_31057;
 wire u0_n_31059;
 wire u0_n_31061;
 wire u0_n_31063;
 wire u0_n_31064;
 wire u0_n_31065;
 wire u0_n_31066;
 wire u0_n_31068;
 wire u0_n_31069;
 wire u0_n_31070;
 wire u0_n_31072;
 wire u0_n_31073;
 wire u0_n_31076;
 wire u0_n_31081;
 wire u0_n_31082;
 wire u0_n_31083;
 wire u0_n_31084;
 wire u0_n_31085;
 wire u0_n_31086;
 wire u0_n_31087;
 wire u0_n_31088;
 wire u0_n_31089;
 wire u0_n_31090;
 wire u0_n_31091;
 wire u0_n_31092;
 wire u0_n_31093;
 wire u0_n_31094;
 wire u0_n_31095;
 wire u0_n_31096;
 wire u0_n_31097;
 wire u0_n_31098;
 wire u0_n_31099;
 wire u0_n_31100;
 wire u0_n_31101;
 wire u0_n_31102;
 wire u0_n_31103;
 wire u0_n_31104;
 wire u0_n_31105;
 wire u0_n_31106;
 wire u0_n_31107;
 wire u0_n_31108;
 wire u0_n_31109;
 wire u0_n_31110;
 wire u0_n_31111;
 wire u0_n_31112;
 wire u0_n_31113;
 wire u0_n_31114;
 wire u0_n_31115;
 wire u0_n_31116;
 wire u0_n_31117;
 wire u0_n_31118;
 wire u0_n_31119;
 wire u0_n_31120;
 wire u0_n_31121;
 wire u0_n_31122;
 wire u0_n_31123;
 wire u0_n_31124;
 wire u0_n_31125;
 wire u0_n_31126;
 wire u0_n_31127;
 wire u0_n_31128;
 wire u0_n_31129;
 wire u0_n_31130;
 wire u0_n_31131;
 wire u0_n_31132;
 wire u0_n_31133;
 wire u0_n_31134;
 wire u0_n_31135;
 wire u0_n_31136;
 wire u0_n_31137;
 wire u0_n_31138;
 wire u0_n_31139;
 wire u0_n_31140;
 wire u0_n_31141;
 wire u0_n_31142;
 wire u0_n_31143;
 wire u0_n_31144;
 wire u0_n_31145;
 wire u0_n_31146;
 wire u0_n_31147;
 wire u0_n_31148;
 wire u0_n_31149;
 wire u0_n_31150;
 wire u0_n_31151;
 wire u0_n_31152;
 wire u0_n_31153;
 wire u0_n_31154;
 wire u0_n_31155;
 wire u0_n_31156;
 wire u0_n_31157;
 wire u0_n_31158;
 wire u0_n_31159;
 wire u0_n_31160;
 wire u0_n_31161;
 wire u0_n_31162;
 wire u0_n_31163;
 wire u0_n_31164;
 wire u0_n_31165;
 wire u0_n_31166;
 wire u0_n_31167;
 wire u0_n_31168;
 wire u0_n_31169;
 wire u0_n_31170;
 wire u0_n_31172;
 wire u0_n_31173;
 wire u0_n_31174;
 wire u0_n_31175;
 wire u0_n_31176;
 wire u0_n_31177;
 wire u0_n_31178;
 wire u0_n_31179;
 wire u0_n_31180;
 wire u0_n_31181;
 wire u0_n_31182;
 wire u0_n_31183;
 wire u0_n_31184;
 wire u0_n_31185;
 wire u0_n_31186;
 wire u0_n_31187;
 wire u0_n_31188;
 wire u0_n_31190;
 wire u0_n_31191;
 wire u0_n_31192;
 wire u0_n_31193;
 wire u0_n_31195;
 wire u0_n_31196;
 wire u0_n_31198;
 wire u0_n_31200;
 wire u0_n_31202;
 wire u0_n_31231;
 wire u0_n_31232;
 wire u0_n_31233;
 wire u0_n_31234;
 wire u0_n_31235;
 wire u0_n_31236;
 wire u0_n_31237;
 wire u0_n_31238;
 wire u0_n_31239;
 wire u0_n_31240;
 wire u0_n_31241;
 wire u0_n_31242;
 wire u0_n_31243;
 wire u0_n_31244;
 wire u0_n_31245;
 wire u0_n_31246;
 wire u0_n_31247;
 wire u0_n_31248;
 wire u0_n_31249;
 wire u0_n_31250;
 wire u0_n_31251;
 wire u0_n_31252;
 wire u0_n_31253;
 wire u0_n_31254;
 wire u0_n_31255;
 wire u0_n_31256;
 wire u0_n_31257;
 wire u0_n_31258;
 wire u0_n_31259;
 wire u0_n_31260;
 wire u0_n_31261;
 wire u0_n_31262;
 wire u0_n_31263;
 wire u0_n_31264;
 wire u0_n_31265;
 wire u0_n_31266;
 wire u0_n_31267;
 wire u0_n_31268;
 wire u0_n_31269;
 wire u0_n_31270;
 wire u0_n_31271;
 wire u0_n_31272;
 wire u0_n_31273;
 wire u0_n_31274;
 wire u0_n_31275;
 wire u0_n_31276;
 wire u0_n_31277;
 wire u0_n_31278;
 wire u0_n_31279;
 wire u0_n_31280;
 wire u0_n_31281;
 wire u0_n_31282;
 wire u0_n_31283;
 wire u0_n_31284;
 wire u0_n_31285;
 wire u0_n_31286;
 wire u0_n_31287;
 wire u0_n_31288;
 wire u0_n_31289;
 wire u0_n_31290;
 wire u0_n_31291;
 wire u0_n_31292;
 wire u0_n_31293;
 wire u0_n_31294;
 wire u0_n_31295;
 wire u0_n_31296;
 wire u0_n_31297;
 wire u0_n_31298;
 wire u0_n_31299;
 wire u0_n_31300;
 wire u0_n_31301;
 wire u0_n_31302;
 wire u0_n_31303;
 wire u0_n_31304;
 wire u0_n_31305;
 wire u0_n_31306;
 wire u0_n_31307;
 wire u0_n_31308;
 wire u0_n_31309;
 wire u0_n_31310;
 wire u0_n_31311;
 wire u0_n_31312;
 wire u0_n_31313;
 wire u0_n_31314;
 wire u0_n_31316;
 wire u0_n_31317;
 wire u0_n_31318;
 wire u0_n_31319;
 wire u0_n_31320;
 wire u0_n_31322;
 wire u0_n_31323;
 wire u0_n_31324;
 wire u0_n_31325;
 wire u0_n_31326;
 wire u0_n_31327;
 wire u0_n_31328;
 wire u0_n_31329;
 wire u0_n_31330;
 wire u0_n_31331;
 wire u0_n_31332;
 wire u0_n_31333;
 wire u0_n_31334;
 wire u0_n_31335;
 wire u0_n_31336;
 wire u0_n_31337;
 wire u0_n_31339;
 wire u0_n_31340;
 wire u0_n_31342;
 wire u0_n_31344;
 wire u0_n_31346;
 wire u0_n_31347;
 wire u0_n_31349;
 wire u0_n_31350;
 wire u0_n_31352;
 wire u0_n_31353;
 wire u0_n_31354;
 wire u0_n_31355;
 wire u0_n_31356;
 wire u0_n_31358;
 wire u0_n_31360;
 wire u0_n_31361;
 wire u0_n_31363;
 wire u0_n_31370;
 wire u0_n_31388;
 wire u0_n_31389;
 wire u0_n_31390;
 wire u0_n_31391;
 wire u0_n_31392;
 wire u0_n_31393;
 wire u0_n_31394;
 wire u0_n_31395;
 wire u0_n_31396;
 wire u0_n_31397;
 wire u0_n_31398;
 wire u0_n_31399;
 wire u0_n_31400;
 wire u0_n_31401;
 wire u0_n_31402;
 wire u0_n_31403;
 wire u0_n_31404;
 wire u0_n_31405;
 wire u0_n_31406;
 wire u0_n_31407;
 wire u0_n_31408;
 wire u0_n_31409;
 wire u0_n_31410;
 wire u0_n_31411;
 wire u0_n_31412;
 wire u0_n_31413;
 wire u0_n_31414;
 wire u0_n_31415;
 wire u0_n_31416;
 wire u0_n_31417;
 wire u0_n_31418;
 wire u0_n_31419;
 wire u0_n_31420;
 wire u0_n_31421;
 wire u0_n_31422;
 wire u0_n_31423;
 wire u0_n_31424;
 wire u0_n_31425;
 wire u0_n_31426;
 wire u0_n_31427;
 wire u0_n_31428;
 wire u0_n_31429;
 wire u0_n_31430;
 wire u0_n_31431;
 wire u0_n_31432;
 wire u0_n_31433;
 wire u0_n_31434;
 wire u0_n_31435;
 wire u0_n_31436;
 wire u0_n_31437;
 wire u0_n_31438;
 wire u0_n_31439;
 wire u0_n_31440;
 wire u0_n_31441;
 wire u0_n_31442;
 wire u0_n_31443;
 wire u0_n_31444;
 wire u0_n_31445;
 wire u0_n_31446;
 wire u0_n_31447;
 wire u0_n_31448;
 wire u0_n_31449;
 wire u0_n_31450;
 wire u0_n_31451;
 wire u0_n_31452;
 wire u0_n_31454;
 wire u0_n_31455;
 wire u0_n_31456;
 wire u0_n_31457;
 wire u0_n_31458;
 wire u0_n_31459;
 wire u0_n_31460;
 wire u0_n_31461;
 wire u0_n_31462;
 wire u0_n_31463;
 wire u0_n_31464;
 wire u0_n_31465;
 wire u0_n_31466;
 wire u0_n_31467;
 wire u0_n_31468;
 wire u0_n_31469;
 wire u0_n_31470;
 wire u0_n_31471;
 wire u0_n_31473;
 wire u0_n_31474;
 wire u0_n_31475;
 wire u0_n_31477;
 wire u0_n_31478;
 wire u0_n_31479;
 wire u0_n_31480;
 wire u0_n_31481;
 wire u0_n_31482;
 wire u0_n_31483;
 wire u0_n_31484;
 wire u0_n_31485;
 wire u0_n_31486;
 wire u0_n_31487;
 wire u0_n_31488;
 wire u0_n_31489;
 wire u0_n_31491;
 wire u0_n_31492;
 wire u0_n_31493;
 wire u0_n_31494;
 wire u0_n_31495;
 wire u0_n_31496;
 wire u0_n_31497;
 wire u0_n_31498;
 wire u0_n_31499;
 wire u0_n_31500;
 wire u0_n_31501;
 wire u0_n_31502;
 wire u0_n_31503;
 wire u0_n_31504;
 wire u0_n_31507;
 wire u0_n_31508;
 wire u0_n_31509;
 wire u0_n_31510;
 wire u0_n_31512;
 wire u0_n_31513;
 wire u0_n_31514;
 wire u0_n_31515;
 wire u0_n_31516;
 wire u0_n_31517;
 wire u0_n_31518;
 wire u0_n_31519;
 wire u0_n_31520;
 wire u0_n_31521;
 wire u0_n_31522;
 wire u0_n_31523;
 wire u0_n_31524;
 wire u0_n_31525;
 wire u0_n_31526;
 wire u0_n_31527;
 wire u0_n_31528;
 wire u0_n_31529;
 wire u0_n_31530;
 wire u0_n_31531;
 wire u0_n_31532;
 wire u0_n_31533;
 wire u0_n_31534;
 wire u0_n_31535;
 wire u0_n_31536;
 wire u0_n_31537;
 wire u0_n_31538;
 wire u0_n_31539;
 wire u0_n_31540;
 wire u0_n_31541;
 wire u0_n_31542;
 wire u0_n_31543;
 wire u0_n_31544;
 wire u0_n_31545;
 wire u0_n_31546;
 wire u0_n_31547;
 wire u0_n_31548;
 wire u0_n_31549;
 wire u0_n_31550;
 wire u0_n_31551;
 wire u0_n_31552;
 wire u0_n_31553;
 wire u0_n_31568;
 wire u0_n_31569;
 wire u0_n_31570;
 wire u0_n_31571;
 wire u0_n_31572;
 wire u0_n_31573;
 wire u0_n_31574;
 wire u0_n_31575;
 wire u0_n_31576;
 wire u0_n_31577;
 wire u0_n_31578;
 wire u0_n_31579;
 wire u0_n_31580;
 wire u0_n_31581;
 wire u0_n_31582;
 wire u0_n_31583;
 wire u0_n_31584;
 wire u0_n_31585;
 wire u0_n_31586;
 wire u0_n_31587;
 wire u0_n_31588;
 wire u0_n_31589;
 wire u0_n_31590;
 wire u0_n_31591;
 wire u0_n_31592;
 wire u0_n_31593;
 wire u0_n_31594;
 wire u0_n_31595;
 wire u0_n_31596;
 wire u0_n_31597;
 wire u0_n_31598;
 wire u0_n_31599;
 wire u0_n_31600;
 wire u0_n_31601;
 wire u0_n_31602;
 wire u0_n_31603;
 wire u0_n_31604;
 wire u0_n_31605;
 wire u0_n_31606;
 wire u0_n_31607;
 wire u0_n_31608;
 wire u0_n_31609;
 wire u0_n_31610;
 wire u0_n_31611;
 wire u0_n_31612;
 wire u0_n_31613;
 wire u0_n_31614;
 wire u0_n_31615;
 wire u0_n_31616;
 wire u0_n_31617;
 wire u0_n_31618;
 wire u0_n_31619;
 wire u0_n_31620;
 wire u0_n_31621;
 wire u0_n_31622;
 wire u0_n_31623;
 wire u0_n_31624;
 wire u0_n_31625;
 wire u0_n_31626;
 wire u0_n_31627;
 wire u0_n_31628;
 wire u0_n_31629;
 wire u0_n_31630;
 wire u0_n_31631;
 wire u0_n_31632;
 wire u0_n_31633;
 wire u0_n_31634;
 wire u0_n_31635;
 wire u0_n_31636;
 wire u0_n_31637;
 wire u0_n_31638;
 wire u0_n_31639;
 wire u0_n_31640;
 wire u0_n_31642;
 wire u0_n_31643;
 wire u0_n_31644;
 wire u0_n_31645;
 wire u0_n_31646;
 wire u0_n_31647;
 wire u0_n_31648;
 wire u0_n_31649;
 wire u0_n_31650;
 wire u0_n_31651;
 wire u0_n_31653;
 wire u0_n_31654;
 wire u0_n_31655;
 wire u0_n_31656;
 wire u0_n_31657;
 wire u0_n_31659;
 wire u0_n_31660;
 wire u0_n_31661;
 wire u0_n_31662;
 wire u0_n_31664;
 wire u0_n_31665;
 wire u0_n_31666;
 wire u0_n_31667;
 wire u0_n_31668;
 wire u0_n_31669;
 wire u0_n_31670;
 wire u0_n_31671;
 wire u0_n_31672;
 wire u0_n_31673;
 wire u0_n_31674;
 wire u0_n_31675;
 wire u0_n_31676;
 wire u0_n_31677;
 wire u0_n_31678;
 wire u0_n_31679;
 wire u0_n_31680;
 wire u0_n_31681;
 wire u0_n_31682;
 wire u0_n_31683;
 wire u0_n_31684;
 wire u0_n_31685;
 wire u0_n_31686;
 wire u0_n_31687;
 wire u0_n_31688;
 wire u0_n_31689;
 wire u0_n_31690;
 wire u0_n_31691;
 wire u0_n_31692;
 wire u0_n_31693;
 wire u0_n_31694;
 wire u0_n_31696;
 wire u0_n_31698;
 wire u0_n_31700;
 wire u0_n_31702;
 wire u0_n_31704;
 wire u0_n_31706;
 wire u0_n_31707;
 wire u0_n_31709;
 wire u0_n_31712;
 wire u0_n_31714;
 wire u0_n_31715;
 wire u0_n_31717;
 wire u0_n_31718;
 wire u0_n_31720;
 wire u0_n_31721;
 wire u0_n_31722;
 wire u0_n_31723;
 wire u0_n_31724;
 wire u0_n_31726;
 wire u0_n_31727;
 wire u0_n_31729;
 wire u0_n_31730;
 wire u0_n_31733;
 wire u0_n_31734;
 wire u0_n_31736;
 wire u0_n_31738;
 wire u0_n_31740;
 wire u0_n_31747;
 wire u0_n_31748;
 wire u0_n_31749;
 wire u0_n_31751;
 wire u0_n_31752;
 wire u0_n_31753;
 wire u0_n_31754;
 wire u0_n_31755;
 wire u0_n_31756;
 wire u0_n_31757;
 wire u0_n_31758;
 wire u0_n_31759;
 wire u0_n_31760;
 wire u0_n_31761;
 wire u0_n_31762;
 wire u0_n_31763;
 wire u0_n_31764;
 wire u0_n_31765;
 wire u0_n_31766;
 wire u0_n_31767;
 wire u0_n_31768;
 wire u0_n_31769;
 wire u0_n_31770;
 wire u0_n_31771;
 wire u0_n_31772;
 wire u0_n_31773;
 wire u0_n_31774;
 wire u0_n_31775;
 wire u0_n_31776;
 wire u0_n_31777;
 wire u0_n_31778;
 wire u0_n_31779;
 wire u0_n_31780;
 wire u0_n_31781;
 wire u0_n_31782;
 wire u0_n_31783;
 wire u0_n_31784;
 wire u0_n_31785;
 wire u0_n_31786;
 wire u0_n_31787;
 wire u0_n_31788;
 wire u0_n_31789;
 wire u0_n_31790;
 wire u0_n_31791;
 wire u0_n_31792;
 wire u0_n_31793;
 wire u0_n_31794;
 wire u0_n_31795;
 wire u0_n_31796;
 wire u0_n_31797;
 wire u0_n_31798;
 wire u0_n_31799;
 wire u0_n_31800;
 wire u0_n_31801;
 wire u0_n_31802;
 wire u0_n_31803;
 wire u0_n_31804;
 wire u0_n_31805;
 wire u0_n_31806;
 wire u0_n_31807;
 wire u0_n_31808;
 wire u0_n_31809;
 wire u0_n_31810;
 wire u0_n_31811;
 wire u0_n_31812;
 wire u0_n_31813;
 wire u0_n_31814;
 wire u0_n_31815;
 wire u0_n_31816;
 wire u0_n_31817;
 wire u0_n_31818;
 wire u0_n_31819;
 wire u0_n_31820;
 wire u0_n_31821;
 wire u0_n_31822;
 wire u0_n_31823;
 wire u0_n_31824;
 wire u0_n_31825;
 wire u0_n_31826;
 wire u0_n_31827;
 wire u0_n_31830;
 wire u0_n_31835;
 wire u0_n_31837;
 wire u0_n_31838;
 wire u0_n_31839;
 wire u0_n_31840;
 wire u0_n_31841;
 wire u0_n_31842;
 wire u0_n_31846;
 wire u0_n_31850;
 wire u0_n_31874;
 wire u0_n_31875;
 wire u0_n_31886;
 wire u0_n_31895;
 wire u0_n_31900;
 wire u0_n_31905;
 wire u0_n_31906;
 wire u0_n_31909;
 wire u0_n_31910;
 wire u0_n_31911;
 wire u0_n_31912;
 wire u0_n_31913;
 wire u0_n_31914;
 wire u0_n_31915;
 wire u0_n_31916;
 wire u0_n_31917;
 wire u0_n_31918;
 wire u0_n_31919;
 wire u0_n_31920;
 wire u0_n_31921;
 wire u0_n_31922;
 wire u0_n_31923;
 wire u0_n_31924;
 wire u0_n_31926;
 wire u0_n_31927;
 wire u0_n_31928;
 wire u0_n_31929;
 wire u0_n_31930;
 wire u0_n_31931;
 wire u0_n_31932;
 wire u0_n_31933;
 wire u0_n_31934;
 wire u0_n_31935;
 wire u0_n_31936;
 wire u0_n_31937;
 wire u0_n_31938;
 wire u0_n_31939;
 wire u0_n_31940;
 wire u0_n_31941;
 wire u0_n_31942;
 wire u0_n_31943;
 wire u0_n_31944;
 wire u0_n_31945;
 wire u0_n_31946;
 wire u0_n_31949;
 wire u0_n_31950;
 wire u0_n_31951;
 wire u0_n_31952;
 wire u0_n_31953;
 wire u0_n_31954;
 wire u0_n_31955;
 wire u0_n_31956;
 wire u0_n_31957;
 wire u0_n_31958;
 wire u0_n_31959;
 wire u0_n_31960;
 wire u0_n_31961;
 wire u0_n_31962;
 wire u0_n_31963;
 wire u0_n_31964;
 wire u0_n_31965;
 wire u0_n_31966;
 wire u0_n_31967;
 wire u0_n_31968;
 wire u0_n_31969;
 wire u0_n_31970;
 wire u0_n_31971;
 wire u0_n_31972;
 wire u0_n_31973;
 wire u0_n_31974;
 wire u0_n_31975;
 wire u0_n_31976;
 wire u0_n_31977;
 wire u0_n_31981;
 wire u0_n_31982;
 wire u0_n_31983;
 wire u0_n_31984;
 wire u0_n_31985;
 wire u0_n_31986;
 wire u0_n_31988;
 wire u0_n_31998;
 wire u0_n_32011;
 wire u0_n_32012;
 wire u0_n_32017;
 wire u0_n_32021;
 wire u0_n_32023;
 wire u0_n_32040;
 wire u0_n_32042;
 wire u0_n_32052;
 wire u0_n_32053;
 wire u0_n_32063;
 wire u0_n_32073;
 wire u0_n_32075;
 wire u0_n_32080;
 wire u0_n_32083;
 wire u0_n_32084;
 wire u0_n_32108;
 wire u0_n_32109;
 wire u0_n_32113;
 wire u0_n_32121;
 wire u0_n_32122;
 wire u0_n_32141;
 wire u0_n_32142;
 wire u0_n_32160;
 wire u0_n_32165;
 wire u0_n_32166;
 wire u0_n_32174;
 wire u0_n_32175;
 wire u0_n_32184;
 wire u0_n_32185;
 wire u0_n_32193;
 wire u0_n_32194;
 wire u0_n_32208;
 wire u0_n_32209;
 wire u0_n_32221;
 wire u0_n_32226;
 wire u0_n_32241;
 wire u0_n_32242;
 wire u0_n_32248;
 wire u0_n_32249;
 wire u0_n_32254;
 wire u0_n_32260;
 wire u0_n_32272;
 wire u0_n_32273;
 wire u0_n_32289;
 wire u0_n_32290;
 wire u0_n_32304;
 wire u0_n_32306;
 wire u0_n_32308;
 wire u0_n_32315;
 wire u0_n_32320;
 wire u0_n_32321;
 wire u0_n_32338;
 wire u0_n_32339;
 wire u0_n_32344;
 wire u0_n_32353;
 wire u0_n_32372;
 wire u0_n_32373;
 wire u0_n_32385;
 wire u0_n_32386;
 wire u0_n_32387;
 wire u0_n_32407;
 wire u0_n_32409;
 wire u0_n_32410;
 wire u0_n_32416;
 wire u0_n_32425;
 wire u0_n_32528;
 wire u0_n_32571;
 wire u0_n_32673;
 wire u0_n_32675;
 wire u0_n_32676;
 wire u0_n_32683;
 wire u0_n_32685;
 wire u0_n_32687;
 wire u0_n_32689;
 wire u0_n_32691;
 wire u0_n_32695;
 wire u0_n_32697;
 wire u0_n_32698;
 wire u0_n_32704;
 wire u0_n_32706;
 wire u0_n_32714;
 wire u0_n_32715;
 wire u0_n_32716;
 wire u0_n_32717;
 wire u0_n_32731;
 wire u0_n_32735;
 wire u0_n_32737;
 wire u0_n_32741;
 wire u0_n_32743;
 wire u0_n_32745;
 wire u0_n_32747;
 wire u0_n_32749;
 wire u0_n_32751;
 wire u0_n_32753;
 wire u0_n_32759;
 wire u0_n_32761;
 wire u0_n_32763;
 wire u0_n_32766;
 wire u0_n_32773;
 wire u0_n_32774;
 wire u0_n_32793;
 wire u0_n_32795;
 wire u0_n_32796;
 wire u0_n_32797;
 wire u0_n_32798;
 wire u0_n_32799;
 wire u0_n_32800;
 wire u0_n_32801;
 wire u0_n_32802;
 wire u0_n_32803;
 wire u0_n_32804;
 wire u0_n_32805;
 wire u0_n_32806;
 wire u0_n_32807;
 wire u0_n_32808;
 wire u0_n_32809;
 wire u0_n_32810;
 wire u0_n_32811;
 wire u0_n_32812;
 wire u0_n_32813;
 wire u0_n_32814;
 wire u0_n_32815;
 wire u0_n_32816;
 wire u0_n_32817;
 wire u0_n_32818;
 wire u0_n_32819;
 wire u0_n_32820;
 wire u0_n_32821;
 wire u0_n_32822;
 wire u0_n_32825;
 wire u0_n_32834;
 wire u0_n_32835;
 wire u0_n_32836;
 wire u0_n_32839;
 wire u0_n_32843;
 wire u0_n_32845;
 wire u0_n_32851;
 wire u0_n_32875;
 wire u0_n_32877;
 wire u0_n_32879;
 wire u0_n_32924;
 wire u0_n_32934;
 wire u0_n_32942;
 wire u0_n_32966;
 wire u0_n_32967;
 wire u0_n_32971;
 wire u0_n_32983;
 wire u0_n_32990;
 wire u0_n_32991;
 wire u0_n_33001;
 wire u0_n_33004;
 wire u0_n_33008;
 wire u0_n_33030;
 wire u0_n_33033;
 wire u0_n_33110;
 wire u0_n_33138;
 wire u0_n_33149;
 wire u0_n_33150;
 wire [3:0] dcnt;
 wire [7:0] sa00;
 wire [7:0] sa01;
 wire [7:0] sa02;
 wire [7:0] sa03;
 wire [7:0] sa10;
 wire [7:0] sa11;
 wire [7:0] sa12;
 wire [7:0] sa13;
 wire [7:0] sa20;
 wire [7:0] sa21;
 wire [7:0] sa22;
 wire [7:0] sa23;
 wire [7:0] sa30;
 wire [7:0] sa31;
 wire [7:0] sa32;
 wire [7:0] sa33;
 wire [127:0] text_in_r;
 wire [3:0] u0_r0_rcnt;
 wire [31:0] u0_rcon;
 wire [30:0] \u0_w[3] ;
 wire [31:0] w0;
 wire [31:0] w1;
 wire [31:0] w2;
 wire [31:0] w3;

 DFFHQNx1_ASAP7_75t_R \dcnt_reg[0]  (.CLK(clk),
    .D(n_1272),
    .QN(dcnt[0]));
 DFFHQNx1_ASAP7_75t_R \dcnt_reg[1]  (.CLK(clk),
    .D(n_1245),
    .QN(dcnt[1]));
 DFFHQNx1_ASAP7_75t_R \dcnt_reg[2]  (.CLK(clk),
    .D(n_1147),
    .QN(dcnt[2]));
 DFFHQNx1_ASAP7_75t_R \dcnt_reg[3]  (.CLK(clk),
    .D(n_1271),
    .QN(dcnt[3]));
 DFFHQNx1_ASAP7_75t_R done_reg (.CLK(clk),
    .D(n_3832),
    .QN(done_3039));
 INVxp33_ASAP7_75t_R drc_bufs (.A(n_95),
    .Y(n_36));
 INVxp33_ASAP7_75t_R drc_bufs111232 (.A(n_95),
    .Y(n_35));
 INVxp33_ASAP7_75t_R drc_bufs111233 (.A(n_95),
    .Y(n_34));
 INVxp33_ASAP7_75t_R drc_bufs111234 (.A(n_95),
    .Y(n_33));
 INVxp33_ASAP7_75t_R drc_bufs111235 (.A(n_95),
    .Y(n_32));
 INVxp33_ASAP7_75t_R drc_bufs111236 (.A(n_95),
    .Y(n_31));
 INVxp33_ASAP7_75t_R drc_bufs111237 (.A(n_95),
    .Y(n_30));
 INVxp33_ASAP7_75t_R drc_bufs111238 (.A(n_95),
    .Y(n_29));
 INVxp33_ASAP7_75t_R drc_bufs111251 (.A(n_95),
    .Y(n_28));
 INVxp33_ASAP7_75t_R drc_bufs111259 (.A(n_95),
    .Y(n_27));
 HB1xp67_ASAP7_75t_L drc_bufs220670 (.A(n_2061),
    .Y(n_1380));
 HB1xp67_ASAP7_75t_R drc_bufs220676 (.A(n_2395),
    .Y(n_1379));
 BUFx2_ASAP7_75t_SL drc_bufs220682 (.A(n_2047),
    .Y(n_1378));
 HB1xp67_ASAP7_75t_R drc_bufs220688 (.A(sa11[6]),
    .Y(n_1377));
 HB1xp67_ASAP7_75t_R drc_bufs220729 (.A(n_2084),
    .Y(n_1372));
 BUFx2_ASAP7_75t_SL drc_bufs220735 (.A(n_8180),
    .Y(n_1371));
 HB1xp67_ASAP7_75t_R drc_bufs220752 (.A(n_2064),
    .Y(n_1370));
 HB1xp67_ASAP7_75t_SL drc_bufs220758 (.A(n_2059),
    .Y(n_1369));
 HB1xp67_ASAP7_75t_R drc_bufs220764 (.A(n_8189),
    .Y(n_1368));
 BUFx2_ASAP7_75t_L drc_bufs220777 (.A(n_2089),
    .Y(n_1366));
 HB1xp67_ASAP7_75t_L drc_bufs220788 (.A(sa02[0]),
    .Y(n_1365));
 HB1xp67_ASAP7_75t_SL drc_bufs220794 (.A(n_2066),
    .Y(n_1364));
 HB1xp67_ASAP7_75t_R drc_bufs220814 (.A(n_8200),
    .Y(n_1361));
 HB1xp67_ASAP7_75t_R drc_bufs220820 (.A(sa20[4]),
    .Y(n_1360));
 HB1xp67_ASAP7_75t_R drc_bufs220826 (.A(n_8212),
    .Y(n_1359));
 HB1xp67_ASAP7_75t_L drc_bufs220832 (.A(n_2057),
    .Y(n_1358));
 HB1xp67_ASAP7_75t_SL drc_bufs220838 (.A(n_2415),
    .Y(n_1357));
 INVxp67_ASAP7_75t_R drc_bufs220882 (.A(n_2411),
    .Y(n_1406));
 HB1xp67_ASAP7_75t_SL drc_bufs220892 (.A(n_2092),
    .Y(n_1374));
 HB1xp67_ASAP7_75t_L drc_bufs220899 (.A(n_2399),
    .Y(n_1389));
 HB1xp67_ASAP7_75t_R drc_bufs220943 (.A(sa30[6]),
    .Y(n_1367));
 HB1xp67_ASAP7_75t_R drc_bufs220950 (.A(n_1938),
    .Y(n_1353));
 BUFx2_ASAP7_75t_L drc_bufs220957 (.A(n_2065),
    .Y(n_1432));
 HB1xp67_ASAP7_75t_SL drc_bufs221271 (.A(\text_out[0]_3160 ),
    .Y(n_9002));
 HB1xp67_ASAP7_75t_SL drc_bufs221274 (.A(\text_out[127]_3047 ),
    .Y(n_9005));
 HB1xp67_ASAP7_75t_SL drc_bufs221277 (.A(\text_out[2]_3162 ),
    .Y(n_9008));
 HB1xp67_ASAP7_75t_SL drc_bufs221280 (.A(\text_out[125]_3045 ),
    .Y(n_9011));
 HB1xp67_ASAP7_75t_SL drc_bufs221283 (.A(\text_out[124]_3044 ),
    .Y(n_9014));
 HB1xp67_ASAP7_75t_SL drc_bufs221286 (.A(\text_out[123]_3043 ),
    .Y(n_9017));
 HB1xp67_ASAP7_75t_SL drc_bufs221289 (.A(\text_out[122]_3042 ),
    .Y(n_9020));
 HB1xp67_ASAP7_75t_SL drc_bufs221292 (.A(\text_out[121]_3041 ),
    .Y(n_9023));
 HB1xp67_ASAP7_75t_SL drc_bufs221295 (.A(\text_out[120]_3040 ),
    .Y(n_9026));
 HB1xp67_ASAP7_75t_SL drc_bufs221298 (.A(\text_out[119]_3079 ),
    .Y(n_9029));
 HB1xp67_ASAP7_75t_SL drc_bufs221301 (.A(\text_out[118]_3078 ),
    .Y(n_9032));
 HB1xp67_ASAP7_75t_SL drc_bufs221304 (.A(\text_out[117]_3077 ),
    .Y(n_9035));
 HB1xp67_ASAP7_75t_SL drc_bufs221307 (.A(\text_out[116]_3076 ),
    .Y(n_9038));
 HB1xp67_ASAP7_75t_SL drc_bufs221310 (.A(\text_out[115]_3075 ),
    .Y(n_9041));
 HB1xp67_ASAP7_75t_SL drc_bufs221313 (.A(\text_out[114]_3074 ),
    .Y(n_9044));
 HB1xp67_ASAP7_75t_SL drc_bufs221316 (.A(\text_out[113]_3073 ),
    .Y(n_9047));
 HB1xp67_ASAP7_75t_SL drc_bufs221319 (.A(\text_out[112]_3072 ),
    .Y(n_9050));
 HB1xp67_ASAP7_75t_SL drc_bufs221322 (.A(\text_out[111]_3111 ),
    .Y(n_9053));
 HB1xp67_ASAP7_75t_SL drc_bufs221325 (.A(\text_out[110]_3110 ),
    .Y(n_9056));
 HB1xp67_ASAP7_75t_SL drc_bufs221328 (.A(\text_out[109]_3109 ),
    .Y(n_9059));
 HB1xp67_ASAP7_75t_SL drc_bufs221331 (.A(\text_out[108]_3108 ),
    .Y(n_9062));
 HB1xp67_ASAP7_75t_SL drc_bufs221334 (.A(\text_out[107]_3107 ),
    .Y(n_9065));
 HB1xp67_ASAP7_75t_SL drc_bufs221337 (.A(\text_out[106]_3106 ),
    .Y(n_9068));
 HB1xp67_ASAP7_75t_SL drc_bufs221340 (.A(\text_out[105]_3105 ),
    .Y(n_9071));
 HB1xp67_ASAP7_75t_SL drc_bufs221343 (.A(\text_out[104]_3104 ),
    .Y(n_9074));
 HB1xp67_ASAP7_75t_SL drc_bufs221346 (.A(\text_out[103]_3143 ),
    .Y(n_9077));
 HB1xp67_ASAP7_75t_SL drc_bufs221349 (.A(\text_out[102]_3142 ),
    .Y(n_9080));
 HB1xp67_ASAP7_75t_SL drc_bufs221352 (.A(\text_out[101]_3141 ),
    .Y(n_9083));
 HB1xp67_ASAP7_75t_SL drc_bufs221355 (.A(\text_out[100]_3140 ),
    .Y(n_9086));
 HB1xp67_ASAP7_75t_SL drc_bufs221358 (.A(\text_out[99]_3139 ),
    .Y(n_9089));
 HB1xp67_ASAP7_75t_SL drc_bufs221361 (.A(\text_out[98]_3138 ),
    .Y(n_9092));
 HB1xp67_ASAP7_75t_SL drc_bufs221364 (.A(\text_out[97]_3137 ),
    .Y(n_9095));
 HB1xp67_ASAP7_75t_SL drc_bufs221367 (.A(\text_out[96]_3136 ),
    .Y(n_9098));
 HB1xp67_ASAP7_75t_SL drc_bufs221370 (.A(\text_out[95]_3055 ),
    .Y(n_9101));
 HB1xp67_ASAP7_75t_SL drc_bufs221373 (.A(\text_out[94]_3054 ),
    .Y(n_9104));
 HB1xp67_ASAP7_75t_SL drc_bufs221376 (.A(\text_out[93]_3053 ),
    .Y(n_9107));
 HB1xp67_ASAP7_75t_SL drc_bufs221379 (.A(\text_out[92]_3052 ),
    .Y(n_9110));
 HB1xp67_ASAP7_75t_SL drc_bufs221382 (.A(\text_out[91]_3051 ),
    .Y(n_9113));
 HB1xp67_ASAP7_75t_SL drc_bufs221385 (.A(\text_out[90]_3050 ),
    .Y(n_9116));
 HB1xp67_ASAP7_75t_SL drc_bufs221388 (.A(\text_out[89]_3049 ),
    .Y(n_9119));
 HB1xp67_ASAP7_75t_SL drc_bufs221391 (.A(\text_out[88]_3048 ),
    .Y(n_9122));
 HB1xp67_ASAP7_75t_SL drc_bufs221394 (.A(\text_out[87]_3087 ),
    .Y(n_9125));
 HB1xp67_ASAP7_75t_SL drc_bufs221397 (.A(\text_out[86]_3086 ),
    .Y(n_9128));
 HB1xp67_ASAP7_75t_SL drc_bufs221400 (.A(\text_out[85]_3085 ),
    .Y(n_9131));
 HB1xp67_ASAP7_75t_SL drc_bufs221403 (.A(\text_out[84]_3084 ),
    .Y(n_9134));
 HB1xp67_ASAP7_75t_SL drc_bufs221406 (.A(\text_out[83]_3083 ),
    .Y(n_9137));
 HB1xp67_ASAP7_75t_SL drc_bufs221409 (.A(\text_out[82]_3082 ),
    .Y(n_9140));
 HB1xp67_ASAP7_75t_SL drc_bufs221412 (.A(\text_out[81]_3081 ),
    .Y(n_9143));
 HB1xp67_ASAP7_75t_SL drc_bufs221415 (.A(\text_out[80]_3080 ),
    .Y(n_9146));
 HB1xp67_ASAP7_75t_SL drc_bufs221418 (.A(\text_out[79]_3119 ),
    .Y(n_9149));
 HB1xp67_ASAP7_75t_SL drc_bufs221421 (.A(\text_out[78]_3118 ),
    .Y(n_9152));
 HB1xp67_ASAP7_75t_SL drc_bufs221424 (.A(\text_out[77]_3117 ),
    .Y(n_9155));
 HB1xp67_ASAP7_75t_SL drc_bufs221427 (.A(\text_out[76]_3116 ),
    .Y(n_9158));
 HB1xp67_ASAP7_75t_SL drc_bufs221430 (.A(\text_out[75]_3115 ),
    .Y(n_9161));
 HB1xp67_ASAP7_75t_SL drc_bufs221433 (.A(\text_out[74]_3114 ),
    .Y(n_9164));
 HB1xp67_ASAP7_75t_SL drc_bufs221436 (.A(\text_out[73]_3113 ),
    .Y(n_9167));
 HB1xp67_ASAP7_75t_SL drc_bufs221439 (.A(\text_out[72]_3112 ),
    .Y(n_9170));
 HB1xp67_ASAP7_75t_SL drc_bufs221442 (.A(\text_out[71]_3151 ),
    .Y(n_9173));
 HB1xp67_ASAP7_75t_SL drc_bufs221445 (.A(\text_out[70]_3150 ),
    .Y(n_9176));
 HB1xp67_ASAP7_75t_SL drc_bufs221448 (.A(\text_out[69]_3149 ),
    .Y(n_9179));
 HB1xp67_ASAP7_75t_SL drc_bufs221451 (.A(\text_out[68]_3148 ),
    .Y(n_9182));
 HB1xp67_ASAP7_75t_SL drc_bufs221454 (.A(\text_out[67]_3147 ),
    .Y(n_9185));
 HB1xp67_ASAP7_75t_SL drc_bufs221457 (.A(\text_out[66]_3146 ),
    .Y(n_9188));
 HB1xp67_ASAP7_75t_SL drc_bufs221460 (.A(\text_out[65]_3145 ),
    .Y(n_9191));
 HB1xp67_ASAP7_75t_SL drc_bufs221463 (.A(\text_out[64]_3144 ),
    .Y(n_9194));
 HB1xp67_ASAP7_75t_SL drc_bufs221466 (.A(\text_out[63]_3063 ),
    .Y(n_9197));
 HB1xp67_ASAP7_75t_SL drc_bufs221469 (.A(\text_out[6]_3166 ),
    .Y(n_9200));
 HB1xp67_ASAP7_75t_SL drc_bufs221472 (.A(\text_out[61]_3061 ),
    .Y(n_9203));
 HB1xp67_ASAP7_75t_SL drc_bufs221475 (.A(\text_out[60]_3060 ),
    .Y(n_9206));
 HB1xp67_ASAP7_75t_SL drc_bufs221478 (.A(\text_out[59]_3059 ),
    .Y(n_9209));
 HB1xp67_ASAP7_75t_SL drc_bufs221481 (.A(\text_out[58]_3058 ),
    .Y(n_9212));
 HB1xp67_ASAP7_75t_SL drc_bufs221484 (.A(\text_out[57]_3057 ),
    .Y(n_9215));
 HB1xp67_ASAP7_75t_SL drc_bufs221487 (.A(\text_out[56]_3056 ),
    .Y(n_9218));
 HB1xp67_ASAP7_75t_SL drc_bufs221490 (.A(\text_out[55]_3095 ),
    .Y(n_9221));
 HB1xp67_ASAP7_75t_SL drc_bufs221493 (.A(\text_out[54]_3094 ),
    .Y(n_9224));
 HB1xp67_ASAP7_75t_SL drc_bufs221496 (.A(\text_out[53]_3093 ),
    .Y(n_9227));
 HB1xp67_ASAP7_75t_SL drc_bufs221499 (.A(\text_out[52]_3092 ),
    .Y(n_9230));
 HB1xp67_ASAP7_75t_SL drc_bufs221502 (.A(\text_out[51]_3091 ),
    .Y(n_9233));
 HB1xp67_ASAP7_75t_SL drc_bufs221505 (.A(\text_out[50]_3090 ),
    .Y(n_9236));
 HB1xp67_ASAP7_75t_SL drc_bufs221508 (.A(\text_out[49]_3089 ),
    .Y(n_9239));
 HB1xp67_ASAP7_75t_SL drc_bufs221511 (.A(\text_out[48]_3088 ),
    .Y(n_9242));
 HB1xp67_ASAP7_75t_SL drc_bufs221514 (.A(\text_out[47]_3127 ),
    .Y(n_9245));
 HB1xp67_ASAP7_75t_SL drc_bufs221517 (.A(\text_out[46]_3126 ),
    .Y(n_9248));
 HB1xp67_ASAP7_75t_SL drc_bufs221520 (.A(\text_out[45]_3125 ),
    .Y(n_9251));
 HB1xp67_ASAP7_75t_SL drc_bufs221523 (.A(\text_out[44]_3124 ),
    .Y(n_9254));
 HB1xp67_ASAP7_75t_SL drc_bufs221526 (.A(\text_out[43]_3123 ),
    .Y(n_9257));
 HB1xp67_ASAP7_75t_SL drc_bufs221529 (.A(\text_out[42]_3122 ),
    .Y(n_9260));
 HB1xp67_ASAP7_75t_SL drc_bufs221532 (.A(\text_out[41]_3121 ),
    .Y(n_9263));
 HB1xp67_ASAP7_75t_SL drc_bufs221535 (.A(\text_out[40]_3120 ),
    .Y(n_9266));
 HB1xp67_ASAP7_75t_SL drc_bufs221538 (.A(\text_out[39]_3159 ),
    .Y(n_9269));
 HB1xp67_ASAP7_75t_SL drc_bufs221541 (.A(\text_out[38]_3158 ),
    .Y(n_9272));
 HB1xp67_ASAP7_75t_SL drc_bufs221544 (.A(\text_out[37]_3157 ),
    .Y(n_9275));
 HB1xp67_ASAP7_75t_SL drc_bufs221547 (.A(\text_out[36]_3156 ),
    .Y(n_9278));
 HB1xp67_ASAP7_75t_SL drc_bufs221550 (.A(\text_out[35]_3155 ),
    .Y(n_9281));
 HB1xp67_ASAP7_75t_SL drc_bufs221553 (.A(\text_out[34]_3154 ),
    .Y(n_9284));
 HB1xp67_ASAP7_75t_SL drc_bufs221556 (.A(\text_out[33]_3153 ),
    .Y(n_9287));
 HB1xp67_ASAP7_75t_SL drc_bufs221559 (.A(\text_out[32]_3152 ),
    .Y(n_9290));
 HB1xp67_ASAP7_75t_SL drc_bufs221562 (.A(\text_out[31]_3071 ),
    .Y(n_9293));
 HB1xp67_ASAP7_75t_SL drc_bufs221565 (.A(\text_out[14]_3134 ),
    .Y(n_9296));
 HB1xp67_ASAP7_75t_SL drc_bufs221568 (.A(\text_out[29]_3069 ),
    .Y(n_9299));
 HB1xp67_ASAP7_75t_SL drc_bufs221571 (.A(\text_out[28]_3068 ),
    .Y(n_9302));
 HB1xp67_ASAP7_75t_SL drc_bufs221574 (.A(\text_out[27]_3067 ),
    .Y(n_9305));
 HB1xp67_ASAP7_75t_SL drc_bufs221577 (.A(\text_out[26]_3066 ),
    .Y(n_9308));
 HB1xp67_ASAP7_75t_SL drc_bufs221580 (.A(\text_out[25]_3065 ),
    .Y(n_9311));
 HB1xp67_ASAP7_75t_SL drc_bufs221583 (.A(\text_out[24]_3064 ),
    .Y(n_9314));
 HB1xp67_ASAP7_75t_SL drc_bufs221586 (.A(\text_out[23]_3103 ),
    .Y(n_9317));
 HB1xp67_ASAP7_75t_SL drc_bufs221589 (.A(\text_out[22]_3102 ),
    .Y(n_9320));
 HB1xp67_ASAP7_75t_SL drc_bufs221592 (.A(\text_out[21]_3101 ),
    .Y(n_9323));
 HB1xp67_ASAP7_75t_SL drc_bufs221595 (.A(\text_out[20]_3100 ),
    .Y(n_9326));
 HB1xp67_ASAP7_75t_SL drc_bufs221598 (.A(\text_out[19]_3099 ),
    .Y(n_9329));
 HB1xp67_ASAP7_75t_SL drc_bufs221601 (.A(\text_out[18]_3098 ),
    .Y(n_9332));
 HB1xp67_ASAP7_75t_SL drc_bufs221604 (.A(\text_out[17]_3097 ),
    .Y(n_9335));
 HB1xp67_ASAP7_75t_SL drc_bufs221607 (.A(\text_out[16]_3096 ),
    .Y(n_9338));
 HB1xp67_ASAP7_75t_SL drc_bufs221610 (.A(\text_out[15]_3135 ),
    .Y(n_9341));
 HB1xp67_ASAP7_75t_SL drc_bufs221613 (.A(\text_out[30]_3070 ),
    .Y(n_9344));
 HB1xp67_ASAP7_75t_SL drc_bufs221616 (.A(\text_out[13]_3133 ),
    .Y(n_9347));
 HB1xp67_ASAP7_75t_SL drc_bufs221619 (.A(\text_out[12]_3132 ),
    .Y(n_9350));
 HB1xp67_ASAP7_75t_SL drc_bufs221622 (.A(\text_out[11]_3131 ),
    .Y(n_9353));
 HB1xp67_ASAP7_75t_SL drc_bufs221625 (.A(\text_out[10]_3130 ),
    .Y(n_9356));
 HB1xp67_ASAP7_75t_SL drc_bufs221628 (.A(\text_out[9]_3129 ),
    .Y(n_9359));
 HB1xp67_ASAP7_75t_SL drc_bufs221631 (.A(\text_out[8]_3128 ),
    .Y(n_9362));
 HB1xp67_ASAP7_75t_SL drc_bufs221634 (.A(\text_out[7]_3167 ),
    .Y(n_9365));
 HB1xp67_ASAP7_75t_SL drc_bufs221637 (.A(\text_out[62]_3062 ),
    .Y(n_9368));
 HB1xp67_ASAP7_75t_SL drc_bufs221640 (.A(\text_out[5]_3165 ),
    .Y(n_9371));
 HB1xp67_ASAP7_75t_SL drc_bufs221643 (.A(\text_out[4]_3164 ),
    .Y(n_9374));
 HB1xp67_ASAP7_75t_SL drc_bufs221646 (.A(\text_out[3]_3163 ),
    .Y(n_9377));
 HB1xp67_ASAP7_75t_SL drc_bufs221649 (.A(\text_out[126]_3046 ),
    .Y(n_9380));
 HB1xp67_ASAP7_75t_SL drc_bufs221652 (.A(\text_out[1]_3161 ),
    .Y(n_9383));
 HB1xp67_ASAP7_75t_SL drc_bufs221655 (.A(done_3039),
    .Y(n_9386));
 INVxp67_ASAP7_75t_R drc_bufs221659 (.A(n_9393),
    .Y(text_out[0]));
 INVxp67_ASAP7_75t_R drc_bufs221660 (.A(n_9002),
    .Y(n_9393));
 INVxp67_ASAP7_75t_R drc_bufs221662 (.A(n_9398),
    .Y(done));
 INVxp67_ASAP7_75t_R drc_bufs221663 (.A(n_9386),
    .Y(n_9398));
 INVxp67_ASAP7_75t_R drc_bufs221665 (.A(n_9403),
    .Y(text_out[1]));
 INVxp67_ASAP7_75t_R drc_bufs221666 (.A(n_9383),
    .Y(n_9403));
 INVxp67_ASAP7_75t_R drc_bufs221668 (.A(n_9408),
    .Y(text_out[126]));
 INVxp67_ASAP7_75t_R drc_bufs221669 (.A(n_9380),
    .Y(n_9408));
 INVxp67_ASAP7_75t_R drc_bufs221671 (.A(n_9413),
    .Y(text_out[3]));
 INVxp67_ASAP7_75t_R drc_bufs221672 (.A(n_9377),
    .Y(n_9413));
 INVxp67_ASAP7_75t_R drc_bufs221674 (.A(n_9418),
    .Y(text_out[4]));
 INVxp67_ASAP7_75t_R drc_bufs221675 (.A(n_9374),
    .Y(n_9418));
 INVxp67_ASAP7_75t_R drc_bufs221677 (.A(n_9423),
    .Y(text_out[5]));
 INVxp67_ASAP7_75t_R drc_bufs221678 (.A(n_9371),
    .Y(n_9423));
 INVxp67_ASAP7_75t_R drc_bufs221680 (.A(n_9428),
    .Y(text_out[62]));
 INVxp67_ASAP7_75t_R drc_bufs221681 (.A(n_9368),
    .Y(n_9428));
 INVxp67_ASAP7_75t_R drc_bufs221683 (.A(n_9433),
    .Y(text_out[7]));
 INVxp67_ASAP7_75t_R drc_bufs221684 (.A(n_9365),
    .Y(n_9433));
 INVxp67_ASAP7_75t_R drc_bufs221686 (.A(n_9438),
    .Y(text_out[8]));
 INVxp67_ASAP7_75t_R drc_bufs221687 (.A(n_9362),
    .Y(n_9438));
 INVxp67_ASAP7_75t_R drc_bufs221689 (.A(n_9443),
    .Y(text_out[9]));
 INVxp67_ASAP7_75t_R drc_bufs221690 (.A(n_9359),
    .Y(n_9443));
 INVxp67_ASAP7_75t_R drc_bufs221692 (.A(n_9448),
    .Y(text_out[10]));
 INVxp67_ASAP7_75t_R drc_bufs221693 (.A(n_9356),
    .Y(n_9448));
 INVxp67_ASAP7_75t_R drc_bufs221695 (.A(n_9453),
    .Y(text_out[11]));
 INVxp67_ASAP7_75t_R drc_bufs221696 (.A(n_9353),
    .Y(n_9453));
 INVxp67_ASAP7_75t_R drc_bufs221698 (.A(n_9458),
    .Y(text_out[12]));
 INVxp67_ASAP7_75t_R drc_bufs221699 (.A(n_9350),
    .Y(n_9458));
 INVxp67_ASAP7_75t_R drc_bufs221701 (.A(n_9463),
    .Y(text_out[13]));
 INVxp67_ASAP7_75t_R drc_bufs221702 (.A(n_9347),
    .Y(n_9463));
 INVxp67_ASAP7_75t_R drc_bufs221704 (.A(n_9468),
    .Y(text_out[30]));
 INVxp67_ASAP7_75t_R drc_bufs221705 (.A(n_9344),
    .Y(n_9468));
 INVxp67_ASAP7_75t_R drc_bufs221707 (.A(n_9473),
    .Y(text_out[15]));
 INVxp67_ASAP7_75t_R drc_bufs221708 (.A(n_9341),
    .Y(n_9473));
 INVxp67_ASAP7_75t_R drc_bufs221710 (.A(n_9478),
    .Y(text_out[16]));
 INVxp67_ASAP7_75t_R drc_bufs221711 (.A(n_9338),
    .Y(n_9478));
 INVxp67_ASAP7_75t_R drc_bufs221713 (.A(n_9483),
    .Y(text_out[17]));
 INVxp67_ASAP7_75t_R drc_bufs221714 (.A(n_9335),
    .Y(n_9483));
 INVxp67_ASAP7_75t_R drc_bufs221716 (.A(n_9488),
    .Y(text_out[18]));
 INVxp67_ASAP7_75t_R drc_bufs221717 (.A(n_9332),
    .Y(n_9488));
 INVxp67_ASAP7_75t_R drc_bufs221719 (.A(n_9493),
    .Y(text_out[19]));
 INVxp67_ASAP7_75t_R drc_bufs221720 (.A(n_9329),
    .Y(n_9493));
 INVxp67_ASAP7_75t_R drc_bufs221722 (.A(n_9498),
    .Y(text_out[20]));
 INVxp67_ASAP7_75t_R drc_bufs221723 (.A(n_9326),
    .Y(n_9498));
 INVxp67_ASAP7_75t_R drc_bufs221725 (.A(n_9503),
    .Y(text_out[21]));
 INVxp67_ASAP7_75t_R drc_bufs221726 (.A(n_9323),
    .Y(n_9503));
 INVxp67_ASAP7_75t_R drc_bufs221728 (.A(n_9508),
    .Y(text_out[22]));
 INVxp67_ASAP7_75t_R drc_bufs221729 (.A(n_9320),
    .Y(n_9508));
 INVxp67_ASAP7_75t_R drc_bufs221731 (.A(n_9513),
    .Y(text_out[23]));
 INVxp67_ASAP7_75t_R drc_bufs221732 (.A(n_9317),
    .Y(n_9513));
 INVxp67_ASAP7_75t_R drc_bufs221734 (.A(n_9518),
    .Y(text_out[24]));
 INVxp67_ASAP7_75t_R drc_bufs221735 (.A(n_9314),
    .Y(n_9518));
 INVxp67_ASAP7_75t_R drc_bufs221737 (.A(n_9523),
    .Y(text_out[25]));
 INVxp67_ASAP7_75t_R drc_bufs221738 (.A(n_9311),
    .Y(n_9523));
 INVxp67_ASAP7_75t_R drc_bufs221740 (.A(n_9528),
    .Y(text_out[26]));
 INVxp67_ASAP7_75t_R drc_bufs221741 (.A(n_9308),
    .Y(n_9528));
 INVxp67_ASAP7_75t_R drc_bufs221743 (.A(n_9533),
    .Y(text_out[27]));
 INVxp67_ASAP7_75t_R drc_bufs221744 (.A(n_9305),
    .Y(n_9533));
 INVxp67_ASAP7_75t_R drc_bufs221746 (.A(n_9538),
    .Y(text_out[28]));
 INVxp67_ASAP7_75t_R drc_bufs221747 (.A(n_9302),
    .Y(n_9538));
 INVxp67_ASAP7_75t_R drc_bufs221749 (.A(n_9543),
    .Y(text_out[29]));
 INVxp67_ASAP7_75t_R drc_bufs221750 (.A(n_9299),
    .Y(n_9543));
 INVxp67_ASAP7_75t_R drc_bufs221752 (.A(n_9548),
    .Y(text_out[14]));
 INVxp67_ASAP7_75t_R drc_bufs221753 (.A(n_9296),
    .Y(n_9548));
 INVxp67_ASAP7_75t_R drc_bufs221755 (.A(n_9553),
    .Y(text_out[31]));
 INVxp67_ASAP7_75t_R drc_bufs221756 (.A(n_9293),
    .Y(n_9553));
 INVxp67_ASAP7_75t_R drc_bufs221758 (.A(n_9558),
    .Y(text_out[32]));
 INVxp67_ASAP7_75t_R drc_bufs221759 (.A(n_9290),
    .Y(n_9558));
 INVxp67_ASAP7_75t_R drc_bufs221761 (.A(n_9563),
    .Y(text_out[33]));
 INVxp67_ASAP7_75t_R drc_bufs221762 (.A(n_9287),
    .Y(n_9563));
 INVxp67_ASAP7_75t_R drc_bufs221764 (.A(n_9568),
    .Y(text_out[34]));
 INVxp67_ASAP7_75t_R drc_bufs221765 (.A(n_9284),
    .Y(n_9568));
 INVxp67_ASAP7_75t_R drc_bufs221767 (.A(n_9573),
    .Y(text_out[35]));
 INVxp67_ASAP7_75t_R drc_bufs221768 (.A(n_9281),
    .Y(n_9573));
 INVxp67_ASAP7_75t_R drc_bufs221770 (.A(n_9578),
    .Y(text_out[36]));
 INVxp67_ASAP7_75t_R drc_bufs221771 (.A(n_9278),
    .Y(n_9578));
 INVxp67_ASAP7_75t_R drc_bufs221773 (.A(n_9583),
    .Y(text_out[37]));
 INVxp67_ASAP7_75t_R drc_bufs221774 (.A(n_9275),
    .Y(n_9583));
 INVxp67_ASAP7_75t_R drc_bufs221776 (.A(n_9588),
    .Y(text_out[38]));
 INVxp67_ASAP7_75t_R drc_bufs221777 (.A(n_9272),
    .Y(n_9588));
 INVxp67_ASAP7_75t_R drc_bufs221779 (.A(n_9593),
    .Y(text_out[39]));
 INVxp67_ASAP7_75t_R drc_bufs221780 (.A(n_9269),
    .Y(n_9593));
 INVxp67_ASAP7_75t_R drc_bufs221782 (.A(n_9598),
    .Y(text_out[40]));
 INVxp67_ASAP7_75t_R drc_bufs221783 (.A(n_9266),
    .Y(n_9598));
 INVxp67_ASAP7_75t_R drc_bufs221785 (.A(n_9603),
    .Y(text_out[41]));
 INVxp67_ASAP7_75t_R drc_bufs221786 (.A(n_9263),
    .Y(n_9603));
 INVxp67_ASAP7_75t_R drc_bufs221788 (.A(n_9608),
    .Y(text_out[42]));
 INVxp67_ASAP7_75t_R drc_bufs221789 (.A(n_9260),
    .Y(n_9608));
 INVxp67_ASAP7_75t_R drc_bufs221791 (.A(n_9613),
    .Y(text_out[43]));
 INVxp67_ASAP7_75t_R drc_bufs221792 (.A(n_9257),
    .Y(n_9613));
 INVxp67_ASAP7_75t_R drc_bufs221794 (.A(n_9618),
    .Y(text_out[44]));
 INVxp67_ASAP7_75t_R drc_bufs221795 (.A(n_9254),
    .Y(n_9618));
 INVxp67_ASAP7_75t_R drc_bufs221797 (.A(n_9623),
    .Y(text_out[45]));
 INVxp67_ASAP7_75t_R drc_bufs221798 (.A(n_9251),
    .Y(n_9623));
 INVxp67_ASAP7_75t_R drc_bufs221800 (.A(n_9628),
    .Y(text_out[46]));
 INVxp67_ASAP7_75t_R drc_bufs221801 (.A(n_9248),
    .Y(n_9628));
 INVxp67_ASAP7_75t_R drc_bufs221803 (.A(n_9633),
    .Y(text_out[47]));
 INVxp67_ASAP7_75t_R drc_bufs221804 (.A(n_9245),
    .Y(n_9633));
 INVxp67_ASAP7_75t_R drc_bufs221806 (.A(n_9638),
    .Y(text_out[48]));
 INVxp67_ASAP7_75t_R drc_bufs221807 (.A(n_9242),
    .Y(n_9638));
 INVxp67_ASAP7_75t_R drc_bufs221809 (.A(n_9643),
    .Y(text_out[49]));
 INVxp67_ASAP7_75t_R drc_bufs221810 (.A(n_9239),
    .Y(n_9643));
 INVxp67_ASAP7_75t_R drc_bufs221812 (.A(n_9648),
    .Y(text_out[50]));
 INVxp67_ASAP7_75t_R drc_bufs221813 (.A(n_9236),
    .Y(n_9648));
 INVxp67_ASAP7_75t_R drc_bufs221815 (.A(n_9653),
    .Y(text_out[51]));
 INVxp67_ASAP7_75t_R drc_bufs221816 (.A(n_9233),
    .Y(n_9653));
 INVxp67_ASAP7_75t_R drc_bufs221818 (.A(n_9658),
    .Y(text_out[52]));
 INVxp67_ASAP7_75t_R drc_bufs221819 (.A(n_9230),
    .Y(n_9658));
 INVxp67_ASAP7_75t_R drc_bufs221821 (.A(n_9663),
    .Y(text_out[53]));
 INVxp67_ASAP7_75t_R drc_bufs221822 (.A(n_9227),
    .Y(n_9663));
 INVxp67_ASAP7_75t_R drc_bufs221824 (.A(n_9668),
    .Y(text_out[54]));
 INVxp67_ASAP7_75t_R drc_bufs221825 (.A(n_9224),
    .Y(n_9668));
 INVxp67_ASAP7_75t_R drc_bufs221827 (.A(n_9673),
    .Y(text_out[55]));
 INVxp67_ASAP7_75t_R drc_bufs221828 (.A(n_9221),
    .Y(n_9673));
 INVxp67_ASAP7_75t_R drc_bufs221830 (.A(n_9678),
    .Y(text_out[56]));
 INVxp67_ASAP7_75t_R drc_bufs221831 (.A(n_9218),
    .Y(n_9678));
 INVxp67_ASAP7_75t_R drc_bufs221833 (.A(n_9683),
    .Y(text_out[57]));
 INVxp67_ASAP7_75t_R drc_bufs221834 (.A(n_9215),
    .Y(n_9683));
 INVxp67_ASAP7_75t_R drc_bufs221836 (.A(n_9688),
    .Y(text_out[58]));
 INVxp67_ASAP7_75t_R drc_bufs221837 (.A(n_9212),
    .Y(n_9688));
 INVxp67_ASAP7_75t_R drc_bufs221839 (.A(n_9693),
    .Y(text_out[59]));
 INVxp67_ASAP7_75t_R drc_bufs221840 (.A(n_9209),
    .Y(n_9693));
 INVxp67_ASAP7_75t_R drc_bufs221842 (.A(n_9698),
    .Y(text_out[60]));
 INVxp67_ASAP7_75t_R drc_bufs221843 (.A(n_9206),
    .Y(n_9698));
 INVxp67_ASAP7_75t_R drc_bufs221845 (.A(n_9703),
    .Y(text_out[61]));
 INVxp67_ASAP7_75t_R drc_bufs221846 (.A(n_9203),
    .Y(n_9703));
 INVxp67_ASAP7_75t_R drc_bufs221848 (.A(n_9708),
    .Y(text_out[6]));
 INVxp67_ASAP7_75t_R drc_bufs221849 (.A(n_9200),
    .Y(n_9708));
 INVxp67_ASAP7_75t_R drc_bufs221851 (.A(n_9713),
    .Y(text_out[63]));
 INVxp67_ASAP7_75t_R drc_bufs221852 (.A(n_9197),
    .Y(n_9713));
 INVxp67_ASAP7_75t_R drc_bufs221854 (.A(n_9718),
    .Y(text_out[64]));
 INVxp67_ASAP7_75t_R drc_bufs221855 (.A(n_9194),
    .Y(n_9718));
 INVxp67_ASAP7_75t_R drc_bufs221857 (.A(n_9723),
    .Y(text_out[65]));
 INVxp67_ASAP7_75t_R drc_bufs221858 (.A(n_9191),
    .Y(n_9723));
 INVxp67_ASAP7_75t_R drc_bufs221860 (.A(n_9728),
    .Y(text_out[66]));
 INVxp67_ASAP7_75t_R drc_bufs221861 (.A(n_9188),
    .Y(n_9728));
 INVxp67_ASAP7_75t_R drc_bufs221863 (.A(n_9733),
    .Y(text_out[67]));
 INVxp67_ASAP7_75t_R drc_bufs221864 (.A(n_9185),
    .Y(n_9733));
 INVxp67_ASAP7_75t_R drc_bufs221866 (.A(n_9738),
    .Y(text_out[68]));
 INVxp67_ASAP7_75t_R drc_bufs221867 (.A(n_9182),
    .Y(n_9738));
 INVxp67_ASAP7_75t_R drc_bufs221869 (.A(n_9743),
    .Y(text_out[69]));
 INVxp67_ASAP7_75t_R drc_bufs221870 (.A(n_9179),
    .Y(n_9743));
 INVxp67_ASAP7_75t_R drc_bufs221872 (.A(n_9748),
    .Y(text_out[70]));
 INVxp67_ASAP7_75t_R drc_bufs221873 (.A(n_9176),
    .Y(n_9748));
 INVxp67_ASAP7_75t_R drc_bufs221875 (.A(n_9753),
    .Y(text_out[71]));
 INVxp67_ASAP7_75t_R drc_bufs221876 (.A(n_9173),
    .Y(n_9753));
 INVxp67_ASAP7_75t_R drc_bufs221878 (.A(n_9758),
    .Y(text_out[72]));
 INVxp67_ASAP7_75t_R drc_bufs221879 (.A(n_9170),
    .Y(n_9758));
 INVxp67_ASAP7_75t_R drc_bufs221881 (.A(n_9763),
    .Y(text_out[73]));
 INVxp67_ASAP7_75t_R drc_bufs221882 (.A(n_9167),
    .Y(n_9763));
 INVxp67_ASAP7_75t_R drc_bufs221884 (.A(n_9768),
    .Y(text_out[74]));
 INVxp67_ASAP7_75t_R drc_bufs221885 (.A(n_9164),
    .Y(n_9768));
 INVxp67_ASAP7_75t_R drc_bufs221887 (.A(n_9773),
    .Y(text_out[75]));
 INVxp67_ASAP7_75t_R drc_bufs221888 (.A(n_9161),
    .Y(n_9773));
 INVxp67_ASAP7_75t_R drc_bufs221890 (.A(n_9778),
    .Y(text_out[76]));
 INVxp67_ASAP7_75t_R drc_bufs221891 (.A(n_9158),
    .Y(n_9778));
 INVxp67_ASAP7_75t_R drc_bufs221893 (.A(n_9783),
    .Y(text_out[77]));
 INVxp67_ASAP7_75t_R drc_bufs221894 (.A(n_9155),
    .Y(n_9783));
 INVxp67_ASAP7_75t_R drc_bufs221896 (.A(n_9788),
    .Y(text_out[78]));
 INVxp67_ASAP7_75t_R drc_bufs221897 (.A(n_9152),
    .Y(n_9788));
 INVxp67_ASAP7_75t_R drc_bufs221899 (.A(n_9793),
    .Y(text_out[79]));
 INVxp67_ASAP7_75t_R drc_bufs221900 (.A(n_9149),
    .Y(n_9793));
 INVxp67_ASAP7_75t_R drc_bufs221902 (.A(n_9798),
    .Y(text_out[80]));
 INVxp67_ASAP7_75t_R drc_bufs221903 (.A(n_9146),
    .Y(n_9798));
 INVxp67_ASAP7_75t_R drc_bufs221905 (.A(n_9803),
    .Y(text_out[81]));
 INVxp67_ASAP7_75t_R drc_bufs221906 (.A(n_9143),
    .Y(n_9803));
 INVxp67_ASAP7_75t_R drc_bufs221908 (.A(n_9808),
    .Y(text_out[82]));
 INVxp67_ASAP7_75t_R drc_bufs221909 (.A(n_9140),
    .Y(n_9808));
 INVxp67_ASAP7_75t_R drc_bufs221911 (.A(n_9813),
    .Y(text_out[83]));
 INVxp67_ASAP7_75t_R drc_bufs221912 (.A(n_9137),
    .Y(n_9813));
 INVxp67_ASAP7_75t_R drc_bufs221914 (.A(n_9818),
    .Y(text_out[84]));
 INVxp67_ASAP7_75t_R drc_bufs221915 (.A(n_9134),
    .Y(n_9818));
 INVxp67_ASAP7_75t_R drc_bufs221917 (.A(n_9823),
    .Y(text_out[85]));
 INVxp67_ASAP7_75t_R drc_bufs221918 (.A(n_9131),
    .Y(n_9823));
 INVxp67_ASAP7_75t_R drc_bufs221920 (.A(n_9828),
    .Y(text_out[86]));
 INVxp67_ASAP7_75t_R drc_bufs221921 (.A(n_9128),
    .Y(n_9828));
 INVxp67_ASAP7_75t_R drc_bufs221923 (.A(n_9833),
    .Y(text_out[87]));
 INVxp67_ASAP7_75t_R drc_bufs221924 (.A(n_9125),
    .Y(n_9833));
 INVxp67_ASAP7_75t_R drc_bufs221926 (.A(n_9838),
    .Y(text_out[88]));
 INVxp67_ASAP7_75t_R drc_bufs221927 (.A(n_9122),
    .Y(n_9838));
 INVxp67_ASAP7_75t_R drc_bufs221929 (.A(n_9843),
    .Y(text_out[89]));
 INVxp67_ASAP7_75t_R drc_bufs221930 (.A(n_9119),
    .Y(n_9843));
 INVxp67_ASAP7_75t_R drc_bufs221932 (.A(n_9848),
    .Y(text_out[90]));
 INVxp67_ASAP7_75t_R drc_bufs221933 (.A(n_9116),
    .Y(n_9848));
 INVxp67_ASAP7_75t_R drc_bufs221935 (.A(n_9853),
    .Y(text_out[91]));
 INVxp67_ASAP7_75t_R drc_bufs221936 (.A(n_9113),
    .Y(n_9853));
 INVxp67_ASAP7_75t_R drc_bufs221938 (.A(n_9858),
    .Y(text_out[92]));
 INVxp67_ASAP7_75t_R drc_bufs221939 (.A(n_9110),
    .Y(n_9858));
 INVxp67_ASAP7_75t_R drc_bufs221941 (.A(n_9863),
    .Y(text_out[93]));
 INVxp67_ASAP7_75t_R drc_bufs221942 (.A(n_9107),
    .Y(n_9863));
 INVxp67_ASAP7_75t_R drc_bufs221944 (.A(n_9868),
    .Y(text_out[94]));
 INVxp67_ASAP7_75t_R drc_bufs221945 (.A(n_9104),
    .Y(n_9868));
 INVxp67_ASAP7_75t_R drc_bufs221947 (.A(n_9873),
    .Y(text_out[95]));
 INVxp67_ASAP7_75t_R drc_bufs221948 (.A(n_9101),
    .Y(n_9873));
 INVxp67_ASAP7_75t_R drc_bufs221950 (.A(n_9878),
    .Y(text_out[96]));
 INVxp67_ASAP7_75t_R drc_bufs221951 (.A(n_9098),
    .Y(n_9878));
 INVxp67_ASAP7_75t_R drc_bufs221953 (.A(n_9883),
    .Y(text_out[97]));
 INVxp67_ASAP7_75t_R drc_bufs221954 (.A(n_9095),
    .Y(n_9883));
 INVxp67_ASAP7_75t_R drc_bufs221956 (.A(n_9888),
    .Y(text_out[98]));
 INVxp67_ASAP7_75t_R drc_bufs221957 (.A(n_9092),
    .Y(n_9888));
 INVxp67_ASAP7_75t_R drc_bufs221959 (.A(n_9893),
    .Y(text_out[99]));
 INVxp67_ASAP7_75t_R drc_bufs221960 (.A(n_9089),
    .Y(n_9893));
 INVxp67_ASAP7_75t_R drc_bufs221962 (.A(n_9898),
    .Y(text_out[100]));
 INVxp67_ASAP7_75t_R drc_bufs221963 (.A(n_9086),
    .Y(n_9898));
 INVxp67_ASAP7_75t_R drc_bufs221965 (.A(n_9903),
    .Y(text_out[101]));
 INVxp67_ASAP7_75t_R drc_bufs221966 (.A(n_9083),
    .Y(n_9903));
 INVxp67_ASAP7_75t_R drc_bufs221968 (.A(n_9908),
    .Y(text_out[102]));
 INVxp67_ASAP7_75t_R drc_bufs221969 (.A(n_9080),
    .Y(n_9908));
 INVxp67_ASAP7_75t_R drc_bufs221971 (.A(n_9913),
    .Y(text_out[103]));
 INVxp67_ASAP7_75t_R drc_bufs221972 (.A(n_9077),
    .Y(n_9913));
 INVxp67_ASAP7_75t_R drc_bufs221974 (.A(n_9918),
    .Y(text_out[104]));
 INVxp67_ASAP7_75t_R drc_bufs221975 (.A(n_9074),
    .Y(n_9918));
 INVxp67_ASAP7_75t_R drc_bufs221977 (.A(n_9923),
    .Y(text_out[105]));
 INVxp67_ASAP7_75t_R drc_bufs221978 (.A(n_9071),
    .Y(n_9923));
 INVxp67_ASAP7_75t_R drc_bufs221980 (.A(n_9928),
    .Y(text_out[106]));
 INVxp67_ASAP7_75t_R drc_bufs221981 (.A(n_9068),
    .Y(n_9928));
 INVxp67_ASAP7_75t_R drc_bufs221983 (.A(n_9933),
    .Y(text_out[107]));
 INVxp67_ASAP7_75t_R drc_bufs221984 (.A(n_9065),
    .Y(n_9933));
 INVxp67_ASAP7_75t_R drc_bufs221986 (.A(n_9938),
    .Y(text_out[108]));
 INVxp67_ASAP7_75t_R drc_bufs221987 (.A(n_9062),
    .Y(n_9938));
 INVxp67_ASAP7_75t_R drc_bufs221989 (.A(n_9943),
    .Y(text_out[109]));
 INVxp67_ASAP7_75t_R drc_bufs221990 (.A(n_9059),
    .Y(n_9943));
 INVxp67_ASAP7_75t_R drc_bufs221992 (.A(n_9948),
    .Y(text_out[110]));
 INVxp67_ASAP7_75t_R drc_bufs221993 (.A(n_9056),
    .Y(n_9948));
 INVxp67_ASAP7_75t_R drc_bufs221995 (.A(n_9953),
    .Y(text_out[111]));
 INVxp67_ASAP7_75t_R drc_bufs221996 (.A(n_9053),
    .Y(n_9953));
 INVxp67_ASAP7_75t_R drc_bufs221998 (.A(n_9958),
    .Y(text_out[112]));
 INVxp67_ASAP7_75t_R drc_bufs221999 (.A(n_9050),
    .Y(n_9958));
 INVxp67_ASAP7_75t_R drc_bufs222001 (.A(n_9963),
    .Y(text_out[113]));
 INVxp67_ASAP7_75t_R drc_bufs222002 (.A(n_9047),
    .Y(n_9963));
 INVxp67_ASAP7_75t_R drc_bufs222004 (.A(n_9968),
    .Y(text_out[114]));
 INVxp67_ASAP7_75t_R drc_bufs222005 (.A(n_9044),
    .Y(n_9968));
 INVxp67_ASAP7_75t_R drc_bufs222007 (.A(n_9973),
    .Y(text_out[115]));
 INVxp67_ASAP7_75t_R drc_bufs222008 (.A(n_9041),
    .Y(n_9973));
 INVxp67_ASAP7_75t_R drc_bufs222010 (.A(n_9978),
    .Y(text_out[116]));
 INVxp67_ASAP7_75t_R drc_bufs222011 (.A(n_9038),
    .Y(n_9978));
 INVxp67_ASAP7_75t_R drc_bufs222013 (.A(n_9983),
    .Y(text_out[117]));
 INVxp67_ASAP7_75t_R drc_bufs222014 (.A(n_9035),
    .Y(n_9983));
 INVxp67_ASAP7_75t_R drc_bufs222016 (.A(n_9988),
    .Y(text_out[118]));
 INVxp67_ASAP7_75t_R drc_bufs222017 (.A(n_9032),
    .Y(n_9988));
 INVxp67_ASAP7_75t_R drc_bufs222019 (.A(n_9993),
    .Y(text_out[119]));
 INVxp67_ASAP7_75t_R drc_bufs222020 (.A(n_9029),
    .Y(n_9993));
 INVxp67_ASAP7_75t_R drc_bufs222022 (.A(n_9998),
    .Y(text_out[120]));
 INVxp67_ASAP7_75t_R drc_bufs222023 (.A(n_9026),
    .Y(n_9998));
 INVxp67_ASAP7_75t_R drc_bufs222025 (.A(n_10003),
    .Y(text_out[121]));
 INVxp67_ASAP7_75t_R drc_bufs222026 (.A(n_9023),
    .Y(n_10003));
 INVxp67_ASAP7_75t_R drc_bufs222028 (.A(n_10008),
    .Y(text_out[122]));
 INVxp67_ASAP7_75t_R drc_bufs222029 (.A(n_9020),
    .Y(n_10008));
 INVxp67_ASAP7_75t_R drc_bufs222031 (.A(n_10013),
    .Y(text_out[123]));
 INVxp67_ASAP7_75t_R drc_bufs222032 (.A(n_9017),
    .Y(n_10013));
 INVxp67_ASAP7_75t_R drc_bufs222034 (.A(n_10018),
    .Y(text_out[124]));
 INVxp67_ASAP7_75t_R drc_bufs222035 (.A(n_9014),
    .Y(n_10018));
 INVxp67_ASAP7_75t_R drc_bufs222037 (.A(n_10023),
    .Y(text_out[125]));
 INVxp67_ASAP7_75t_R drc_bufs222038 (.A(n_9011),
    .Y(n_10023));
 INVxp67_ASAP7_75t_R drc_bufs222040 (.A(n_10028),
    .Y(text_out[2]));
 INVxp67_ASAP7_75t_R drc_bufs222041 (.A(n_9008),
    .Y(n_10028));
 INVxp67_ASAP7_75t_R drc_bufs222043 (.A(n_10033),
    .Y(text_out[127]));
 INVxp67_ASAP7_75t_R drc_bufs222044 (.A(n_9005),
    .Y(n_10033));
 HB1xp67_ASAP7_75t_R drc_bufs222840 (.A(w3[7]),
    .Y(n_11346));
 HB1xp67_ASAP7_75t_L drc_bufs222864 (.A(w3[18]),
    .Y(n_11371));
 HB1xp67_ASAP7_75t_R drc_bufs222923 (.A(w3[11]),
    .Y(n_11435));
 HB1xp67_ASAP7_75t_R drc_bufs222944 (.A(w3[3]),
    .Y(n_11457));
 HB1xp67_ASAP7_75t_R drc_bufs222968 (.A(w3[0]),
    .Y(n_11482));
 HB1xp67_ASAP7_75t_R drc_bufs222992 (.A(w3[5]),
    .Y(n_11507));
 INVxp33_ASAP7_75t_R fopt (.A(n_1452),
    .Y(n_1453));
 INVx1_ASAP7_75t_R fopt11 (.A(n_2060),
    .Y(n_1430));
 INVx1_ASAP7_75t_R fopt14 (.A(n_8625),
    .Y(n_8629));
 INVx1_ASAP7_75t_SL fopt15 (.A(w3[4]),
    .Y(n_8625));
 INVxp33_ASAP7_75t_R fopt2 (.A(n_2416),
    .Y(n_1452));
 INVx2_ASAP7_75t_SL fopt21 (.A(w3[4]),
    .Y(n_8623));
 BUFx2_ASAP7_75t_L fopt220079 (.A(n_2045),
    .Y(n_1450));
 BUFx2_ASAP7_75t_SL fopt220087 (.A(n_2394),
    .Y(n_1449));
 BUFx2_ASAP7_75t_L fopt220103 (.A(n_2058),
    .Y(n_1448));
 HB1xp67_ASAP7_75t_L fopt220108 (.A(n_2058),
    .Y(n_1447));
 BUFx2_ASAP7_75t_L fopt220118 (.A(n_2425),
    .Y(n_1446));
 BUFx3_ASAP7_75t_L fopt220136 (.A(n_2067),
    .Y(n_1444));
 INVxp33_ASAP7_75t_R fopt220161 (.A(n_2053),
    .Y(n_1441));
 BUFx2_ASAP7_75t_R fopt220168 (.A(n_2054),
    .Y(n_1440));
 BUFx2_ASAP7_75t_L fopt220177 (.A(n_2048),
    .Y(n_1439));
 INVxp67_ASAP7_75t_R fopt220182 (.A(n_1437),
    .Y(n_1438));
 INVxp33_ASAP7_75t_R fopt220183 (.A(n_2048),
    .Y(n_1437));
 INVxp67_ASAP7_75t_SL fopt220213 (.A(n_1434),
    .Y(n_1435));
 HB1xp67_ASAP7_75t_SL fopt220216 (.A(n_2042),
    .Y(n_1433));
 HB1xp67_ASAP7_75t_R fopt220238 (.A(n_2060),
    .Y(n_1352));
 INVx2_ASAP7_75t_L fopt220239 (.A(n_1430),
    .Y(n_1431));
 INVx2_ASAP7_75t_L fopt220259 (.A(n_1436),
    .Y(n_1429));
 INVx2_ASAP7_75t_SL fopt220260 (.A(n_2393),
    .Y(n_1436));
 BUFx3_ASAP7_75t_SL fopt220287 (.A(sa03[4]),
    .Y(n_1425));
 INVxp67_ASAP7_75t_L fopt220288 (.A(n_1426),
    .Y(n_1427));
 INVxp67_ASAP7_75t_SL fopt220290 (.A(sa03[4]),
    .Y(n_1426));
 BUFx2_ASAP7_75t_SL fopt220304 (.A(n_2082),
    .Y(n_1424));
 BUFx2_ASAP7_75t_L fopt220320 (.A(n_2075),
    .Y(n_1423));
 BUFx2_ASAP7_75t_L fopt220330 (.A(n_2400),
    .Y(n_1422));
 INVxp67_ASAP7_75t_R fopt220333 (.A(n_1420),
    .Y(n_1421));
 INVxp33_ASAP7_75t_R fopt220334 (.A(n_2400),
    .Y(n_1420));
 BUFx2_ASAP7_75t_L fopt220349 (.A(n_2062),
    .Y(n_1419));
 BUFx2_ASAP7_75t_R fopt220362 (.A(n_2063),
    .Y(n_1418));
 INVx2_ASAP7_75t_L fopt220377 (.A(n_1416),
    .Y(n_1417));
 INVxp33_ASAP7_75t_R fopt220391 (.A(n_1414),
    .Y(n_1415));
 INVxp33_ASAP7_75t_R fopt220392 (.A(n_2427),
    .Y(n_1414));
 BUFx2_ASAP7_75t_R fopt220394 (.A(n_2427),
    .Y(n_1413));
 INVxp67_ASAP7_75t_R fopt220403 (.A(n_2091),
    .Y(n_1411));
 HB1xp67_ASAP7_75t_SL fopt220409 (.A(n_2090),
    .Y(n_1412));
 INVx1_ASAP7_75t_R fopt220423 (.A(n_1409),
    .Y(n_1346));
 INVx1_ASAP7_75t_L fopt220424 (.A(n_1410),
    .Y(n_1409));
 HB1xp67_ASAP7_75t_SL fopt220425 (.A(sa33[6]),
    .Y(n_1410));
 HB1xp67_ASAP7_75t_R fopt220435 (.A(n_1408),
    .Y(n_1407));
 BUFx2_ASAP7_75t_L fopt220436 (.A(n_2411),
    .Y(n_1408));
 BUFx2_ASAP7_75t_L fopt220451 (.A(n_2435),
    .Y(n_1405));
 BUFx2_ASAP7_75t_SL fopt220462 (.A(n_1810),
    .Y(n_1808));
 INVxp67_ASAP7_75t_R fopt220472 (.A(n_1402),
    .Y(n_1403));
 INVxp67_ASAP7_75t_R fopt220473 (.A(n_1404),
    .Y(n_1402));
 BUFx2_ASAP7_75t_SL fopt220477 (.A(n_8211),
    .Y(n_1404));
 HB1xp67_ASAP7_75t_SL fopt220485 (.A(n_2072),
    .Y(n_1401));
 HB1xp67_ASAP7_75t_R fopt220493 (.A(n_2410),
    .Y(n_1400));
 INVxp67_ASAP7_75t_R fopt220505 (.A(n_1443),
    .Y(n_1399));
 INVxp67_ASAP7_75t_R fopt220506 (.A(n_2397),
    .Y(n_1443));
 HB1xp67_ASAP7_75t_L fopt220507 (.A(n_2397),
    .Y(n_1398));
 INVxp67_ASAP7_75t_R fopt220517 (.A(n_1396),
    .Y(n_1397));
 INVxp33_ASAP7_75t_R fopt220518 (.A(n_1933),
    .Y(n_1396));
 INVxp67_ASAP7_75t_R fopt220532 (.A(n_1393),
    .Y(n_1394));
 INVxp33_ASAP7_75t_R fopt220534 (.A(n_1395),
    .Y(n_1393));
 BUFx2_ASAP7_75t_R fopt220535 (.A(sa22[6]),
    .Y(n_1395));
 HB1xp67_ASAP7_75t_L fopt220544 (.A(n_2083),
    .Y(n_1392));
 INVx1_ASAP7_75t_R fopt220558 (.A(n_2078),
    .Y(n_1391));
 HB1xp67_ASAP7_75t_R fopt220571 (.A(n_2043),
    .Y(n_1390));
 INVx2_ASAP7_75t_L fopt220572 (.A(n_2042),
    .Y(n_1434));
 BUFx2_ASAP7_75t_SL fopt220595 (.A(sa11[4]),
    .Y(n_1387));
 INVx1_ASAP7_75t_L fopt220614 (.A(n_2056),
    .Y(n_1416));
 BUFx2_ASAP7_75t_L fopt220623 (.A(sa01[4]),
    .Y(n_1386));
 INVx2_ASAP7_75t_SL fopt220627 (.A(n_1384),
    .Y(n_1385));
 INVxp67_ASAP7_75t_R fopt220638 (.A(n_2435),
    .Y(n_1383));
 HB1xp67_ASAP7_75t_L fopt220654 (.A(n_2428),
    .Y(n_1382));
 BUFx2_ASAP7_75t_L fopt220664 (.A(n_2078),
    .Y(n_1381));
 HB1xp67_ASAP7_75t_L fopt220695 (.A(n_2424),
    .Y(n_1376));
 BUFx3_ASAP7_75t_SL fopt220708 (.A(sa30[4]),
    .Y(n_1375));
 HB1xp67_ASAP7_75t_L fopt220723 (.A(n_2088),
    .Y(n_1373));
 INVxp67_ASAP7_75t_R fopt220805 (.A(n_1337),
    .Y(n_1362));
 INVxp67_ASAP7_75t_SL fopt220808 (.A(n_1362),
    .Y(n_1363));
 BUFx4f_ASAP7_75t_SL fopt220860 (.A(n_2387),
    .Y(n_1633));
 INVxp67_ASAP7_75t_R fopt220876 (.A(n_1355),
    .Y(n_1356));
 BUFx2_ASAP7_75t_L fopt220918 (.A(n_2053),
    .Y(n_1354));
 INVxp67_ASAP7_75t_SL fopt220933 (.A(n_2072),
    .Y(n_1355));
 INVx1_ASAP7_75t_SL fopt220993 (.A(w3[19]),
    .Y(n_8652));
 INVxp67_ASAP7_75t_R fopt221011 (.A(n_8656),
    .Y(n_8668));
 INVx1_ASAP7_75t_SL fopt221014 (.A(w3[19]),
    .Y(n_8656));
 INVxp67_ASAP7_75t_L fopt221020 (.A(n_8245),
    .Y(n_8679));
 INVx2_ASAP7_75t_SL fopt221021 (.A(n_8245),
    .Y(n_8678));
 INVxp67_ASAP7_75t_R fopt221022 (.A(n_8688),
    .Y(n_8687));
 INVx2_ASAP7_75t_SL fopt221023 (.A(n_8245),
    .Y(n_8688));
 INVx2_ASAP7_75t_SL fopt221030 (.A(n_8690),
    .Y(n_8691));
 BUFx2_ASAP7_75t_SL fopt221031 (.A(n_1351),
    .Y(n_8690));
 INVx1_ASAP7_75t_SL fopt221039 (.A(n_8703),
    .Y(n_8702));
 BUFx3_ASAP7_75t_SL fopt221042 (.A(n_1351),
    .Y(n_8703));
 INVxp67_ASAP7_75t_R fopt221043 (.A(n_8720),
    .Y(n_8719));
 INVxp67_ASAP7_75t_L fopt221044 (.A(n_1351),
    .Y(n_8720));
 INVx1_ASAP7_75t_SL fopt221050 (.A(n_8280),
    .Y(n_8723));
 INVxp67_ASAP7_75t_L fopt221055 (.A(n_8733),
    .Y(n_8732));
 HB1xp67_ASAP7_75t_L fopt221056 (.A(n_8221),
    .Y(n_8733));
 INVxp67_ASAP7_75t_L fopt221058 (.A(n_8221),
    .Y(n_8738));
 INVx3_ASAP7_75t_SL fopt221062 (.A(w3[1]),
    .Y(n_8742));
 INVxp67_ASAP7_75t_SL fopt221072 (.A(n_8747),
    .Y(n_8748));
 INVxp67_ASAP7_75t_R fopt221073 (.A(w3[1]),
    .Y(n_8747));
 INVxp33_ASAP7_75t_R fopt221081 (.A(n_8760),
    .Y(n_8766));
 INVx3_ASAP7_75t_SL fopt221082 (.A(n_8253),
    .Y(n_8760));
 INVx1_ASAP7_75t_R fopt221088 (.A(n_8771),
    .Y(n_8770));
 INVx3_ASAP7_75t_SL fopt221089 (.A(n_8307),
    .Y(n_8771));
 INVxp33_ASAP7_75t_R fopt221090 (.A(n_8780),
    .Y(n_8779));
 INVx1_ASAP7_75t_SL fopt221091 (.A(n_8239),
    .Y(n_8780));
 INVx2_ASAP7_75t_SL fopt221095 (.A(n_8783),
    .Y(n_8785));
 BUFx2_ASAP7_75t_SL fopt221096 (.A(n_8239),
    .Y(n_8783));
 INVx1_ASAP7_75t_SL fopt221098 (.A(n_579),
    .Y(n_8789));
 INVx2_ASAP7_75t_SL fopt221106 (.A(n_8299),
    .Y(n_8792));
 INVx1_ASAP7_75t_SL fopt221126 (.A(n_8801),
    .Y(n_8820));
 INVx2_ASAP7_75t_R fopt221139 (.A(n_8833),
    .Y(n_8831));
 INVx3_ASAP7_75t_SL fopt221143 (.A(w3[23]),
    .Y(n_8833));
 INVx1_ASAP7_75t_SL fopt221145 (.A(u0_n_29390),
    .Y(n_8847));
 INVx2_ASAP7_75t_L fopt221161 (.A(n_8851),
    .Y(n_8856));
 INVx2_ASAP7_75t_SL fopt221163 (.A(w3[9]),
    .Y(n_8851));
 INVxp67_ASAP7_75t_SL fopt221169 (.A(n_8879),
    .Y(n_8877));
 INVxp67_ASAP7_75t_L fopt221171 (.A(n_8881),
    .Y(n_8879));
 INVx1_ASAP7_75t_SL fopt221172 (.A(n_8872),
    .Y(n_8881));
 INVx3_ASAP7_75t_SL fopt221173 (.A(n_8301),
    .Y(n_8872));
 INVxp67_ASAP7_75t_SL fopt221178 (.A(n_8884),
    .Y(n_8887));
 INVx1_ASAP7_75t_SL fopt221179 (.A(n_8234),
    .Y(n_8884));
 INVx1_ASAP7_75t_SL fopt221185 (.A(n_8894),
    .Y(n_8896));
 INVx4_ASAP7_75t_SL fopt221188 (.A(n_8894),
    .Y(n_8899));
 INVx1_ASAP7_75t_SL fopt221196 (.A(n_8896),
    .Y(n_8908));
 INVx4_ASAP7_75t_SL fopt221204 (.A(n_8899),
    .Y(n_8912));
 INVx6_ASAP7_75t_SL fopt221206 (.A(sa32[4]),
    .Y(n_8894));
 INVxp67_ASAP7_75t_SL fopt221208 (.A(n_8923),
    .Y(n_8922));
 INVx2_ASAP7_75t_L fopt221212 (.A(n_8335),
    .Y(n_8923));
 INVxp33_ASAP7_75t_R fopt221216 (.A(n_8933),
    .Y(n_8932));
 INVx2_ASAP7_75t_SL fopt221219 (.A(n_8261),
    .Y(n_8933));
 INVx2_ASAP7_75t_L fopt221238 (.A(n_8946),
    .Y(n_8942));
 INVx2_ASAP7_75t_SL fopt221241 (.A(w3[28]),
    .Y(n_8946));
 BUFx3_ASAP7_75t_L fopt222901 (.A(w3[8]),
    .Y(n_11401));
 INVx4_ASAP7_75t_SL fopt24 (.A(w3[14]),
    .Y(n_8801));
 INVx2_ASAP7_75t_SL fopt27 (.A(n_8963),
    .Y(n_8964));
 BUFx3_ASAP7_75t_SL fopt29 (.A(w3[28]),
    .Y(n_8963));
 BUFx2_ASAP7_75t_L fopt8 (.A(n_2416),
    .Y(n_1451));
 BUFx2_ASAP7_75t_L fopt9 (.A(n_2396),
    .Y(n_1442));
 OAI22xp5_ASAP7_75t_SL g109565 (.A1(n_40),
    .A2(n_1325),
    .B1(n_112),
    .B2(n_451),
    .Y(n_1335));
 AOI21xp5_ASAP7_75t_SL g109566 (.A1(n_1313),
    .A2(n_112),
    .B(n_974),
    .Y(n_1334));
 OAI22xp5_ASAP7_75t_SL g109567 (.A1(n_40),
    .A2(n_1305),
    .B1(n_112),
    .B2(n_541),
    .Y(n_1333));
 OAI22xp5_ASAP7_75t_SL g109568 (.A1(n_40),
    .A2(n_1295),
    .B1(n_112),
    .B2(n_556),
    .Y(n_1332));
 OAI222xp33_ASAP7_75t_SL g109569 (.A1(n_1274),
    .A2(n_8290),
    .B1(n_1275),
    .B2(n_156),
    .C1(n_458),
    .C2(n_112),
    .Y(n_1331));
 OAI22xp5_ASAP7_75t_SL g109570 (.A1(n_1287),
    .A2(n_40),
    .B1(n_112),
    .B2(n_549),
    .Y(n_1330));
 OAI22xp5_ASAP7_75t_SL g109642 (.A1(n_40),
    .A2(n_1250),
    .B1(n_112),
    .B2(n_533),
    .Y(n_1329));
 XNOR2xp5_ASAP7_75t_SL g109643 (.A(n_1228),
    .B(n_421),
    .Y(n_1328));
 XOR2xp5_ASAP7_75t_SL g109644 (.A(n_1244),
    .B(n_900),
    .Y(n_1327));
 XOR2xp5_ASAP7_75t_SL g109645 (.A(n_1226),
    .B(n_713),
    .Y(n_1326));
 XOR2xp5_ASAP7_75t_SL g109646 (.A(n_1236),
    .B(n_666),
    .Y(n_1325));
 XOR2xp5_ASAP7_75t_SL g109648 (.A(n_1219),
    .B(n_1124),
    .Y(n_1324));
 XOR2xp5_ASAP7_75t_SL g109649 (.A(n_1157),
    .B(n_910),
    .Y(n_1323));
 XOR2xp5_ASAP7_75t_SL g109650 (.A(n_1232),
    .B(n_389),
    .Y(n_1322));
 XOR2xp5_ASAP7_75t_SL g109651 (.A(n_1230),
    .B(n_87),
    .Y(n_1321));
 XOR2xp5_ASAP7_75t_SL g109652 (.A(n_1224),
    .B(n_420),
    .Y(n_1320));
 XOR2xp5_ASAP7_75t_SL g109653 (.A(n_1239),
    .B(n_411),
    .Y(n_1319));
 XOR2xp5_ASAP7_75t_SL g109654 (.A(n_1165),
    .B(n_1095),
    .Y(n_1318));
 XOR2xp5_ASAP7_75t_SL g109655 (.A(n_26),
    .B(n_900),
    .Y(n_1317));
 XOR2xp5_ASAP7_75t_SL g109656 (.A(n_1092),
    .B(n_1233),
    .Y(n_1316));
 XOR2xp5_ASAP7_75t_SL g109657 (.A(n_1235),
    .B(n_1090),
    .Y(n_1315));
 XOR2xp5_ASAP7_75t_SL g109658 (.A(n_1231),
    .B(n_1020),
    .Y(n_1314));
 XOR2xp5_ASAP7_75t_SL g109659 (.A(n_1225),
    .B(n_700),
    .Y(n_1313));
 XOR2xp5_ASAP7_75t_SL g109660 (.A(n_1223),
    .B(n_1082),
    .Y(n_1312));
 XOR2xp5_ASAP7_75t_SL g109661 (.A(n_1222),
    .B(n_993),
    .Y(n_1311));
 XOR2xp5_ASAP7_75t_SL g109662 (.A(n_1218),
    .B(n_1009),
    .Y(n_1310));
 XOR2xp5_ASAP7_75t_SL g109663 (.A(n_17),
    .B(n_1071),
    .Y(n_1309));
 XOR2xp5_ASAP7_75t_SL g109664 (.A(n_1217),
    .B(n_432),
    .Y(n_1308));
 XOR2xp5_ASAP7_75t_SL g109665 (.A(n_1216),
    .B(n_1067),
    .Y(n_1307));
 XOR2xp5_ASAP7_75t_SL g109666 (.A(n_1215),
    .B(n_1065),
    .Y(n_1306));
 XOR2xp5_ASAP7_75t_SL g109667 (.A(n_1214),
    .B(n_697),
    .Y(n_1305));
 XOR2xp5_ASAP7_75t_SL g109668 (.A(n_1242),
    .B(n_1064),
    .Y(n_1304));
 XOR2xp5_ASAP7_75t_SL g109669 (.A(n_1155),
    .B(n_82),
    .Y(n_1303));
 XOR2xp5_ASAP7_75t_SL g109670 (.A(n_1151),
    .B(n_1008),
    .Y(n_1302));
 XOR2xp5_ASAP7_75t_SL g109671 (.A(n_1153),
    .B(n_18),
    .Y(n_1301));
 XOR2xp5_ASAP7_75t_SL g109672 (.A(n_1154),
    .B(n_1049),
    .Y(n_1300));
 XOR2xp5_ASAP7_75t_SL g109673 (.A(n_1037),
    .B(n_1159),
    .Y(n_1299));
 XOR2xp5_ASAP7_75t_SL g109674 (.A(n_1161),
    .B(n_1006),
    .Y(n_1298));
 XOR2xp5_ASAP7_75t_SL g109675 (.A(n_1162),
    .B(n_1025),
    .Y(n_1297));
 XOR2xp5_ASAP7_75t_SL g109676 (.A(n_1163),
    .B(n_1017),
    .Y(n_1296));
 XOR2xp5_ASAP7_75t_SL g109677 (.A(n_1164),
    .B(n_438),
    .Y(n_1295));
 XOR2xp5_ASAP7_75t_SL g109678 (.A(n_1238),
    .B(n_1002),
    .Y(n_1294));
 XOR2xp5_ASAP7_75t_SL g109679 (.A(n_1240),
    .B(n_1001),
    .Y(n_1293));
 XOR2xp5_ASAP7_75t_SL g109680 (.A(n_1234),
    .B(n_999),
    .Y(n_1292));
 XOR2xp5_ASAP7_75t_SL g109681 (.A(n_1229),
    .B(n_998),
    .Y(n_1291));
 XOR2xp5_ASAP7_75t_SL g109682 (.A(n_1220),
    .B(n_997),
    .Y(n_1290));
 XOR2xp5_ASAP7_75t_SL g109683 (.A(n_1241),
    .B(n_996),
    .Y(n_1289));
 XOR2xp5_ASAP7_75t_SL g109684 (.A(n_1237),
    .B(n_985),
    .Y(n_1288));
 XOR2xp5_ASAP7_75t_SL g109685 (.A(n_1152),
    .B(n_433),
    .Y(n_1287));
 XOR2xp5_ASAP7_75t_SL g109686 (.A(n_1169),
    .B(n_643),
    .Y(n_1286));
 XOR2xp5_ASAP7_75t_SL g109687 (.A(n_1227),
    .B(n_8789),
    .Y(n_1285));
 XOR2xp5_ASAP7_75t_SL g109688 (.A(n_1168),
    .B(n_579),
    .Y(n_1284));
 XOR2xp5_ASAP7_75t_SL g109689 (.A(n_13),
    .B(n_1156),
    .Y(n_1283));
 XOR2xp5_ASAP7_75t_SL g109690 (.A(n_74),
    .B(n_1167),
    .Y(n_1282));
 XOR2xp5_ASAP7_75t_SL g109691 (.A(n_572),
    .B(n_1158),
    .Y(n_1281));
 XOR2xp5_ASAP7_75t_SL g109692 (.A(n_1160),
    .B(n_75),
    .Y(n_1280));
 OAI22xp5_ASAP7_75t_SL g109693 (.A1(n_40),
    .A2(n_1175),
    .B1(n_112),
    .B2(n_503),
    .Y(n_1279));
 XOR2xp5_ASAP7_75t_SL g109694 (.A(n_1166),
    .B(n_663),
    .Y(n_1278));
 XOR2xp5_ASAP7_75t_SL g109695 (.A(n_1243),
    .B(n_401),
    .Y(n_1277));
 XOR2xp5_ASAP7_75t_SL g109696 (.A(n_1150),
    .B(n_21),
    .Y(n_1276));
 AOI22xp5_ASAP7_75t_SL g109699 (.A1(n_565),
    .A2(n_1149),
    .B1(n_566),
    .B2(n_1148),
    .Y(n_1275));
 AOI22xp5_ASAP7_75t_SL g109700 (.A1(n_566),
    .A2(n_1149),
    .B1(n_565),
    .B2(n_1148),
    .Y(n_1274));
 XNOR2xp5_ASAP7_75t_L g109702 (.A(n_1004),
    .B(n_1078),
    .Y(n_1273));
 OA21x2_ASAP7_75t_R g109703 (.A1(dcnt[0]),
    .A2(n_1055),
    .B(n_379),
    .Y(n_1272));
 AOI31xp33_ASAP7_75t_R g109704 (.A1(n_1054),
    .A2(n_921),
    .A3(dcnt[3]),
    .B(n_380),
    .Y(n_1271));
 XOR2xp5_ASAP7_75t_SL g109705 (.A(n_989),
    .B(n_758),
    .Y(n_1270));
 XOR2xp5_ASAP7_75t_SL g109706 (.A(n_1133),
    .B(n_719),
    .Y(n_1269));
 XNOR2xp5_ASAP7_75t_SL g109707 (.A(n_988),
    .B(n_755),
    .Y(n_1268));
 XOR2xp5_ASAP7_75t_SL g109708 (.A(n_975),
    .B(n_1127),
    .Y(n_1267));
 XOR2xp5_ASAP7_75t_SL g109709 (.A(n_1122),
    .B(n_1123),
    .Y(n_1266));
 XOR2xp5_ASAP7_75t_SL g109710 (.A(n_707),
    .B(n_1121),
    .Y(n_1265));
 XNOR2xp5_ASAP7_75t_SL g109711 (.A(n_1119),
    .B(n_615),
    .Y(n_1264));
 XOR2xp5_ASAP7_75t_SL g109712 (.A(n_1005),
    .B(n_752),
    .Y(n_1263));
 XOR2xp5_ASAP7_75t_L g109713 (.A(n_1108),
    .B(n_1110),
    .Y(n_1262));
 XOR2xp5_ASAP7_75t_SL g109714 (.A(n_1107),
    .B(n_976),
    .Y(n_1261));
 XOR2xp5_ASAP7_75t_L g109716 (.A(n_15),
    .B(n_750),
    .Y(n_1260));
 XOR2xp5_ASAP7_75t_L g109717 (.A(n_1102),
    .B(n_982),
    .Y(n_1259));
 XOR2xp5_ASAP7_75t_L g109718 (.A(n_1099),
    .B(n_716),
    .Y(n_1258));
 XOR2xp5_ASAP7_75t_L g109719 (.A(n_1098),
    .B(n_749),
    .Y(n_1257));
 XOR2xp5_ASAP7_75t_SL g109720 (.A(n_1011),
    .B(n_747),
    .Y(n_1256));
 XOR2xp5_ASAP7_75t_L g109721 (.A(n_1093),
    .B(n_666),
    .Y(n_1255));
 XOR2xp5_ASAP7_75t_L g109722 (.A(n_1088),
    .B(n_702),
    .Y(n_1254));
 XOR2xp5_ASAP7_75t_SL g109723 (.A(n_1087),
    .B(n_745),
    .Y(n_1253));
 XOR2xp5_ASAP7_75t_SL g109724 (.A(n_1012),
    .B(n_744),
    .Y(n_1252));
 XNOR2xp5_ASAP7_75t_SL g109725 (.A(n_1091),
    .B(n_906),
    .Y(n_1251));
 XOR2xp5_ASAP7_75t_L g109726 (.A(n_1085),
    .B(n_743),
    .Y(n_1250));
 XOR2xp5_ASAP7_75t_SL g109727 (.A(n_1083),
    .B(n_742),
    .Y(n_1249));
 XNOR2xp5_ASAP7_75t_SL g109728 (.A(n_984),
    .B(n_741),
    .Y(n_1248));
 XOR2xp5_ASAP7_75t_SL g109729 (.A(n_980),
    .B(n_1079),
    .Y(n_1247));
 XOR2xp5_ASAP7_75t_L g109730 (.A(n_1077),
    .B(n_740),
    .Y(n_1246));
 OA21x2_ASAP7_75t_R g109731 (.A1(n_887),
    .A2(n_1055),
    .B(n_379),
    .Y(n_1245));
 XNOR2xp5_ASAP7_75t_SL g109732 (.A(n_1135),
    .B(n_756),
    .Y(n_1244));
 XOR2xp5_ASAP7_75t_SL g109733 (.A(n_25),
    .B(n_891),
    .Y(n_1243));
 XNOR2xp5_ASAP7_75t_SL g109734 (.A(n_911),
    .B(n_1111),
    .Y(n_1242));
 XNOR2xp5_ASAP7_75t_SL g109735 (.A(n_1100),
    .B(n_628),
    .Y(n_1241));
 AOI22xp5_ASAP7_75t_SL g109736 (.A1(n_1146),
    .A2(n_9000),
    .B1(n_1145),
    .B2(n_599),
    .Y(n_1240));
 XNOR2xp5_ASAP7_75t_SL g109737 (.A(n_1101),
    .B(n_8274),
    .Y(n_1239));
 XNOR2xp5_ASAP7_75t_L g109738 (.A(n_14),
    .B(n_388),
    .Y(n_1238));
 XNOR2xp5_ASAP7_75t_SL g109739 (.A(n_1094),
    .B(n_588),
    .Y(n_1237));
 XNOR2xp5_ASAP7_75t_SL g109740 (.A(n_8336),
    .B(n_1118),
    .Y(n_1236));
 XNOR2xp5_ASAP7_75t_SL g109742 (.A(n_994),
    .B(n_605),
    .Y(n_1235));
 XNOR2xp5_ASAP7_75t_SL g109743 (.A(n_1117),
    .B(n_572),
    .Y(n_1234));
 XNOR2xp5_ASAP7_75t_SL g109744 (.A(n_1089),
    .B(n_746),
    .Y(n_1233));
 XNOR2xp5_ASAP7_75t_SL g109745 (.A(n_1116),
    .B(n_169),
    .Y(n_1232));
 XNOR2xp5_ASAP7_75t_SL g109746 (.A(n_701),
    .B(n_1019),
    .Y(n_1231));
 XNOR2xp5_ASAP7_75t_SL g109747 (.A(n_1114),
    .B(n_89),
    .Y(n_1230));
 XNOR2xp5_ASAP7_75t_SL g109748 (.A(n_1112),
    .B(n_75),
    .Y(n_1229));
 XOR2xp5_ASAP7_75t_L g109749 (.A(n_1136),
    .B(n_8336),
    .Y(n_1228));
 XNOR2xp5_ASAP7_75t_SL g109750 (.A(n_1010),
    .B(n_1084),
    .Y(n_1227));
 XNOR2xp5_ASAP7_75t_SL g109751 (.A(n_977),
    .B(n_8328),
    .Y(n_1226));
 XNOR2xp5_ASAP7_75t_SL g109752 (.A(n_981),
    .B(n_8304),
    .Y(n_1225));
 XNOR2xp5_ASAP7_75t_SL g109753 (.A(n_342),
    .B(n_1106),
    .Y(n_1224));
 XNOR2xp5_ASAP7_75t_L g109754 (.A(n_1081),
    .B(n_82),
    .Y(n_1223));
 XNOR2xp5_ASAP7_75t_L g109755 (.A(n_1080),
    .B(n_13),
    .Y(n_1222));
 XNOR2xp5_ASAP7_75t_SL g109756 (.A(n_1125),
    .B(n_754),
    .Y(n_1221));
 XNOR2xp5_ASAP7_75t_SL g109757 (.A(n_1103),
    .B(n_912),
    .Y(n_1220));
 XNOR2xp5_ASAP7_75t_L g109758 (.A(n_889),
    .B(n_1000),
    .Y(n_1219));
 XNOR2xp5_ASAP7_75t_SL g109759 (.A(n_1072),
    .B(n_74),
    .Y(n_1218));
 XNOR2xp5_ASAP7_75t_L g109760 (.A(n_1069),
    .B(n_8330),
    .Y(n_1217));
 XNOR2xp5_ASAP7_75t_L g109762 (.A(n_20),
    .B(n_603),
    .Y(n_1216));
 XNOR2xp5_ASAP7_75t_SL g109763 (.A(n_992),
    .B(n_663),
    .Y(n_1215));
 XOR2xp5_ASAP7_75t_SL g109764 (.A(n_979),
    .B(n_200),
    .Y(n_1214));
 XOR2xp5_ASAP7_75t_SL g109766 (.A(n_1130),
    .B(n_391),
    .Y(n_1213));
 XOR2xp5_ASAP7_75t_L g109767 (.A(n_1022),
    .B(n_641),
    .Y(n_1212));
 XOR2xp5_ASAP7_75t_SL g109768 (.A(n_1034),
    .B(n_615),
    .Y(n_1211));
 XOR2xp5_ASAP7_75t_SL g109769 (.A(n_1038),
    .B(n_410),
    .Y(n_1210));
 XOR2xp5_ASAP7_75t_L g109770 (.A(n_1048),
    .B(n_1051),
    .Y(n_1209));
 XOR2xp5_ASAP7_75t_SL g109771 (.A(n_1062),
    .B(n_429),
    .Y(n_1208));
 XOR2xp5_ASAP7_75t_SL g109772 (.A(n_22),
    .B(n_1014),
    .Y(n_1207));
 XOR2xp5_ASAP7_75t_SL g109773 (.A(n_1113),
    .B(n_1142),
    .Y(n_1206));
 XNOR2xp5_ASAP7_75t_SL g109774 (.A(n_1046),
    .B(n_983),
    .Y(n_1205));
 XOR2xp5_ASAP7_75t_SL g109775 (.A(n_1047),
    .B(n_696),
    .Y(n_1204));
 XNOR2xp5_ASAP7_75t_SL g109776 (.A(n_990),
    .B(n_1042),
    .Y(n_1203));
 XOR2xp5_ASAP7_75t_SL g109777 (.A(n_987),
    .B(n_1044),
    .Y(n_1202));
 XOR2xp5_ASAP7_75t_L g109778 (.A(n_23),
    .B(n_430),
    .Y(n_1201));
 XOR2xp5_ASAP7_75t_SL g109779 (.A(n_1120),
    .B(n_1015),
    .Y(n_1200));
 XOR2xp5_ASAP7_75t_SL g109780 (.A(n_986),
    .B(n_1126),
    .Y(n_1199));
 XOR2xp5_ASAP7_75t_SL g109781 (.A(n_1128),
    .B(n_1129),
    .Y(n_1198));
 XOR2xp5_ASAP7_75t_L g109782 (.A(n_1033),
    .B(n_1032),
    .Y(n_1197));
 XOR2xp5_ASAP7_75t_SL g109783 (.A(n_1030),
    .B(n_978),
    .Y(n_1196));
 XNOR2xp5_ASAP7_75t_SL g109784 (.A(n_1134),
    .B(n_633),
    .Y(n_1195));
 XOR2xp5_ASAP7_75t_SL g109785 (.A(n_1138),
    .B(n_1140),
    .Y(n_1194));
 XOR2xp5_ASAP7_75t_SL g109786 (.A(n_1097),
    .B(n_565),
    .Y(n_1193));
 XNOR2xp5_ASAP7_75t_L g109787 (.A(n_1045),
    .B(n_417),
    .Y(n_1192));
 XOR2xp5_ASAP7_75t_SL g109789 (.A(n_1131),
    .B(n_415),
    .Y(n_1190));
 XOR2xp5_ASAP7_75t_SL g109790 (.A(n_1139),
    .B(n_414),
    .Y(n_1189));
 XNOR2xp5_ASAP7_75t_SL g109791 (.A(n_1029),
    .B(n_387),
    .Y(n_1188));
 XNOR2xp5_ASAP7_75t_L g109792 (.A(n_1074),
    .B(n_9001),
    .Y(n_1187));
 XOR2xp5_ASAP7_75t_SL g109793 (.A(n_1066),
    .B(n_8789),
    .Y(n_1186));
 XOR2xp5_ASAP7_75t_L g109794 (.A(n_1039),
    .B(n_74),
    .Y(n_1185));
 AOI22xp33_ASAP7_75t_L g109795 (.A1(n_10),
    .A2(n_1059),
    .B1(n_577),
    .B2(n_1058),
    .Y(n_1184));
 XNOR2xp5_ASAP7_75t_SL g109796 (.A(n_1041),
    .B(n_572),
    .Y(n_1183));
 XNOR2xp5_ASAP7_75t_SL g109797 (.A(n_1028),
    .B(n_439),
    .Y(n_1182));
 XNOR2xp5_ASAP7_75t_L g109798 (.A(n_995),
    .B(n_736),
    .Y(n_1181));
 XOR2xp5_ASAP7_75t_SL g109799 (.A(n_1076),
    .B(n_413),
    .Y(n_1180));
 XOR2xp5_ASAP7_75t_SL g109800 (.A(n_24),
    .B(n_664),
    .Y(n_1179));
 XOR2xp5_ASAP7_75t_SL g109801 (.A(n_1132),
    .B(n_396),
    .Y(n_1178));
 XOR2xp5_ASAP7_75t_SL g109802 (.A(n_1031),
    .B(n_409),
    .Y(n_1177));
 XOR2xp5_ASAP7_75t_SL g109803 (.A(n_1104),
    .B(n_399),
    .Y(n_1176));
 XOR2xp5_ASAP7_75t_SL g109804 (.A(n_1096),
    .B(n_402),
    .Y(n_1175));
 XOR2xp5_ASAP7_75t_L g109805 (.A(n_1086),
    .B(n_403),
    .Y(n_1174));
 XNOR2xp5_ASAP7_75t_SL g109806 (.A(n_1075),
    .B(n_404),
    .Y(n_1173));
 XOR2xp5_ASAP7_75t_SL g109807 (.A(n_1073),
    .B(n_406),
    .Y(n_1172));
 XOR2xp5_ASAP7_75t_SL g109808 (.A(n_1063),
    .B(n_664),
    .Y(n_1171));
 XOR2xp5_ASAP7_75t_SL g109809 (.A(n_1053),
    .B(n_407),
    .Y(n_1170));
 XNOR2xp5_ASAP7_75t_SL g109810 (.A(n_1109),
    .B(n_629),
    .Y(n_1169));
 XNOR2xp5_ASAP7_75t_SL g109811 (.A(n_1070),
    .B(n_635),
    .Y(n_1168));
 XNOR2xp5_ASAP7_75t_SL g109812 (.A(n_1026),
    .B(n_576),
    .Y(n_1167));
 XNOR2xp5_ASAP7_75t_SL g109813 (.A(n_1137),
    .B(n_90),
    .Y(n_1166));
 XNOR2xp5_ASAP7_75t_SL g109814 (.A(n_1003),
    .B(n_591),
    .Y(n_1165));
 AOI22xp5_ASAP7_75t_SL g109815 (.A1(n_8318),
    .A2(n_1056),
    .B1(n_187),
    .B2(n_1057),
    .Y(n_1164));
 XNOR2xp5_ASAP7_75t_SL g109816 (.A(n_1016),
    .B(n_710),
    .Y(n_1163));
 XOR2xp5_ASAP7_75t_L g109817 (.A(n_1024),
    .B(n_88),
    .Y(n_1162));
 XNOR2xp5_ASAP7_75t_SL g109818 (.A(n_1027),
    .B(n_693),
    .Y(n_1161));
 XNOR2xp5_ASAP7_75t_SL g109819 (.A(n_1021),
    .B(n_1035),
    .Y(n_1160));
 XOR2xp5_ASAP7_75t_SL g109820 (.A(n_87),
    .B(n_1036),
    .Y(n_1159));
 XNOR2xp5_ASAP7_75t_SL g109821 (.A(n_1007),
    .B(n_1040),
    .Y(n_1158));
 XNOR2xp5_ASAP7_75t_SL g109822 (.A(n_1115),
    .B(n_665),
    .Y(n_1157));
 XNOR2xp5_ASAP7_75t_SL g109823 (.A(n_695),
    .B(n_1013),
    .Y(n_1156));
 XNOR2xp5_ASAP7_75t_SL g109824 (.A(n_1043),
    .B(n_895),
    .Y(n_1155));
 XNOR2xp5_ASAP7_75t_SL g109825 (.A(n_991),
    .B(n_629),
    .Y(n_1154));
 XNOR2xp5_ASAP7_75t_SL g109826 (.A(n_1050),
    .B(n_665),
    .Y(n_1153));
 XNOR2xp5_ASAP7_75t_L g109827 (.A(n_1052),
    .B(n_8344),
    .Y(n_1152));
 AOI22xp5_ASAP7_75t_SL g109828 (.A1(n_10),
    .A2(n_1060),
    .B1(n_577),
    .B2(n_1061),
    .Y(n_1151));
 XNOR2xp5_ASAP7_75t_SL g109829 (.A(n_890),
    .B(n_1018),
    .Y(n_1150));
 NOR2xp33_ASAP7_75t_R g109830 (.A(n_40),
    .B(n_1143),
    .Y(n_1149));
 A2O1A1Ixp33_ASAP7_75t_R g109831 (.A1(dcnt[2]),
    .A2(n_384),
    .B(n_920),
    .C(n_1054),
    .Y(n_1147));
 NOR2xp33_ASAP7_75t_R g109832 (.A(n_40),
    .B(n_1144),
    .Y(n_1148));
 INVx1_ASAP7_75t_SL g109833 (.A(n_1145),
    .Y(n_1146));
 INVxp67_ASAP7_75t_L g109834 (.A(n_1143),
    .Y(n_1144));
 HB1xp67_ASAP7_75t_SL g109835 (.A(n_1141),
    .Y(n_1142));
 OAI22xp5_ASAP7_75t_L g109837 (.A1(n_960),
    .A2(n_913),
    .B1(n_959),
    .B2(n_914),
    .Y(n_1140));
 XNOR2xp5_ASAP7_75t_SL g109838 (.A(n_428),
    .B(n_759),
    .Y(n_1139));
 AOI22xp5_ASAP7_75t_SL g109839 (.A1(n_603),
    .A2(n_903),
    .B1(n_604),
    .B2(n_904),
    .Y(n_1138));
 OAI22xp5_ASAP7_75t_SL g109841 (.A1(n_7),
    .A2(n_631),
    .B1(n_928),
    .B2(n_630),
    .Y(n_1137));
 XNOR2xp5_ASAP7_75t_SL g109842 (.A(n_422),
    .B(n_8337),
    .Y(n_1136));
 XOR2xp5_ASAP7_75t_SL g109843 (.A(n_918),
    .B(n_395),
    .Y(n_1135));
 OAI22xp5_ASAP7_75t_L g109844 (.A1(n_685),
    .A2(n_658),
    .B1(n_686),
    .B2(n_657),
    .Y(n_1134));
 OAI22xp5_ASAP7_75t_SL g109845 (.A1(n_373),
    .A2(n_660),
    .B1(w0[12]),
    .B2(n_659),
    .Y(n_1145));
 AOI22xp5_ASAP7_75t_L g109846 (.A1(n_934),
    .A2(n_597),
    .B1(n_933),
    .B2(n_598),
    .Y(n_1133));
 AOI22xp5_ASAP7_75t_SL g109847 (.A1(n_972),
    .A2(n_583),
    .B1(n_973),
    .B2(n_584),
    .Y(n_1132));
 XNOR2xp5_ASAP7_75t_L g109848 (.A(n_9),
    .B(n_73),
    .Y(n_1131));
 AOI22xp5_ASAP7_75t_SL g109849 (.A1(n_970),
    .A2(n_583),
    .B1(n_971),
    .B2(n_584),
    .Y(n_1130));
 XOR2xp5_ASAP7_75t_SL g109850 (.A(n_639),
    .B(n_708),
    .Y(n_1129));
 AOI22xp5_ASAP7_75t_L g109851 (.A1(n_568),
    .A2(n_899),
    .B1(n_9001),
    .B2(n_898),
    .Y(n_1128));
 OAI22xp5_ASAP7_75t_L g109852 (.A1(n_280),
    .A2(n_608),
    .B1(w2[31]),
    .B2(n_607),
    .Y(n_1127));
 OAI22xp5_ASAP7_75t_L g109853 (.A1(n_927),
    .A2(n_569),
    .B1(n_71),
    .B2(n_926),
    .Y(n_1126));
 XNOR2xp5_ASAP7_75t_SL g109854 (.A(n_423),
    .B(n_51),
    .Y(n_1143));
 OAI22xp5_ASAP7_75t_SL g109855 (.A1(n_673),
    .A2(n_916),
    .B1(n_674),
    .B2(n_915),
    .Y(n_1125));
 OAI22xp5_ASAP7_75t_SL g109856 (.A1(n_304),
    .A2(n_901),
    .B1(w1[12]),
    .B2(n_902),
    .Y(n_1124));
 XNOR2xp5_ASAP7_75t_L g109857 (.A(n_712),
    .B(n_230),
    .Y(n_1123));
 AOI22xp5_ASAP7_75t_SL g109858 (.A1(w1[13]),
    .A2(n_581),
    .B1(n_263),
    .B2(n_582),
    .Y(n_1122));
 AOI22xp5_ASAP7_75t_SL g109859 (.A1(n_684),
    .A2(n_619),
    .B1(n_683),
    .B2(n_618),
    .Y(n_1121));
 AOI22xp5_ASAP7_75t_SL g109860 (.A1(n_924),
    .A2(n_577),
    .B1(n_925),
    .B2(n_10),
    .Y(n_1120));
 OAI22xp5_ASAP7_75t_L g109861 (.A1(n_929),
    .A2(n_585),
    .B1(n_930),
    .B2(n_586),
    .Y(n_1119));
 XOR2xp5_ASAP7_75t_SL g109863 (.A(n_706),
    .B(n_8313),
    .Y(n_1118));
 XOR2xp5_ASAP7_75t_SL g109864 (.A(n_892),
    .B(w2[9]),
    .Y(n_1117));
 XOR2xp5_ASAP7_75t_SL g109865 (.A(n_715),
    .B(n_8318),
    .Y(n_1116));
 OAI22xp5_ASAP7_75t_SL g109866 (.A1(n_967),
    .A2(n_907),
    .B1(n_8995),
    .B2(n_908),
    .Y(n_1115));
 XOR2xp5_ASAP7_75t_SL g109867 (.A(n_398),
    .B(n_6),
    .Y(n_1114));
 OAI22xp5_ASAP7_75t_L g109868 (.A1(n_965),
    .A2(n_896),
    .B1(n_964),
    .B2(n_897),
    .Y(n_1113));
 XOR2xp5_ASAP7_75t_SL g109869 (.A(n_656),
    .B(w2[12]),
    .Y(n_1112));
 OAI22xp5_ASAP7_75t_SL g109870 (.A1(n_8220),
    .A2(n_895),
    .B1(n_168),
    .B2(n_894),
    .Y(n_1111));
 XNOR2xp5_ASAP7_75t_L g109871 (.A(n_717),
    .B(n_8329),
    .Y(n_1110));
 XOR2xp5_ASAP7_75t_SL g109872 (.A(n_705),
    .B(n_626),
    .Y(n_1109));
 AOI22xp33_ASAP7_75t_R g109873 (.A1(w2[13]),
    .A2(n_72),
    .B1(n_255),
    .B2(n_73),
    .Y(n_1108));
 AOI22xp5_ASAP7_75t_SL g109874 (.A1(n_267),
    .A2(n_649),
    .B1(w2[14]),
    .B2(n_648),
    .Y(n_1107));
 AOI22xp5_ASAP7_75t_SL g109875 (.A1(n_77),
    .A2(w2[15]),
    .B1(n_254),
    .B2(n_76),
    .Y(n_1106));
 XNOR2xp5_ASAP7_75t_SL g109876 (.A(n_425),
    .B(n_400),
    .Y(n_1105));
 AOI22xp5_ASAP7_75t_SL g109877 (.A1(n_963),
    .A2(n_78),
    .B1(n_962),
    .B2(n_79),
    .Y(n_1104));
 OAI22xp5_ASAP7_75t_L g109878 (.A1(n_8851),
    .A2(n_83),
    .B1(n_8856),
    .B2(n_84),
    .Y(n_1103));
 XNOR2xp5_ASAP7_75t_L g109880 (.A(n_426),
    .B(n_8344),
    .Y(n_1102));
 OAI22xp5_ASAP7_75t_L g109882 (.A1(u0_n_32715),
    .A2(n_78),
    .B1(w3[31]),
    .B2(n_79),
    .Y(n_1101));
 XOR2xp5_ASAP7_75t_SL g109883 (.A(n_601),
    .B(w3[12]),
    .Y(n_1100));
 XNOR2xp5_ASAP7_75t_SL g109884 (.A(n_718),
    .B(n_617),
    .Y(n_1099));
 XNOR2xp5_ASAP7_75t_L g109885 (.A(n_386),
    .B(n_588),
    .Y(n_1098));
 XNOR2xp5_ASAP7_75t_L g109886 (.A(n_392),
    .B(n_748),
    .Y(n_1097));
 OAI22xp5_ASAP7_75t_SL g109887 (.A1(n_687),
    .A2(n_9000),
    .B1(n_688),
    .B2(n_599),
    .Y(n_1096));
 OAI22xp5_ASAP7_75t_SL g109888 (.A1(n_301),
    .A2(n_652),
    .B1(w0[1]),
    .B2(n_653),
    .Y(n_1095));
 XOR2xp5_ASAP7_75t_SL g109889 (.A(n_427),
    .B(n_8337),
    .Y(n_1094));
 XNOR2xp5_ASAP7_75t_L g109890 (.A(n_703),
    .B(n_390),
    .Y(n_1093));
 AOI22xp5_ASAP7_75t_L g109891 (.A1(n_58),
    .A2(n_896),
    .B1(n_57),
    .B2(n_897),
    .Y(n_1092));
 OAI22xp5_ASAP7_75t_SL g109892 (.A1(n_937),
    .A2(n_597),
    .B1(n_938),
    .B2(n_598),
    .Y(n_1091));
 OAI22xp5_ASAP7_75t_SL g109893 (.A1(n_245),
    .A2(n_650),
    .B1(w0[4]),
    .B2(n_651),
    .Y(n_1090));
 OAI22xp5_ASAP7_75t_L g109894 (.A1(n_8227),
    .A2(n_919),
    .B1(n_210),
    .B2(n_918),
    .Y(n_1089));
 AOI22xp5_ASAP7_75t_L g109895 (.A1(n_940),
    .A2(n_654),
    .B1(n_939),
    .B2(n_655),
    .Y(n_1088));
 AOI22xp5_ASAP7_75t_SL g109896 (.A1(n_680),
    .A2(n_905),
    .B1(n_679),
    .B2(n_906),
    .Y(n_1087));
 AOI22xp33_ASAP7_75t_R g109897 (.A1(n_8996),
    .A2(n_573),
    .B1(n_958),
    .B2(n_574),
    .Y(n_1086));
 XNOR2xp5_ASAP7_75t_SL g109898 (.A(n_726),
    .B(n_727),
    .Y(n_1085));
 OAI22xp5_ASAP7_75t_SL g109899 (.A1(n_282),
    .A2(n_638),
    .B1(w1[1]),
    .B2(n_639),
    .Y(n_1084));
 OAI22xp5_ASAP7_75t_SL g109900 (.A1(n_612),
    .A2(n_261),
    .B1(w0[31]),
    .B2(n_611),
    .Y(n_1083));
 OAI22xp33_ASAP7_75t_R g109901 (.A1(n_8220),
    .A2(n_86),
    .B1(n_168),
    .B2(n_85),
    .Y(n_1082));
 OAI22xp5_ASAP7_75t_SL g109902 (.A1(n_319),
    .A2(n_916),
    .B1(w1[3]),
    .B2(n_915),
    .Y(n_1081));
 OAI22xp5_ASAP7_75t_SL g109903 (.A1(n_266),
    .A2(n_637),
    .B1(w1[4]),
    .B2(n_636),
    .Y(n_1080));
 XNOR2xp5_ASAP7_75t_L g109904 (.A(n_699),
    .B(n_8254),
    .Y(n_1079));
 XNOR2xp5_ASAP7_75t_L g109905 (.A(n_739),
    .B(n_165),
    .Y(n_1078));
 XNOR2xp5_ASAP7_75t_L g109906 (.A(n_412),
    .B(n_698),
    .Y(n_1077));
 AOI22xp5_ASAP7_75t_L g109907 (.A1(n_586),
    .A2(n_8997),
    .B1(n_585),
    .B2(n_950),
    .Y(n_1076));
 OAI22xp5_ASAP7_75t_SL g109908 (.A1(n_953),
    .A2(n_585),
    .B1(n_954),
    .B2(n_586),
    .Y(n_1075));
 XNOR2xp5_ASAP7_75t_L g109909 (.A(n_385),
    .B(n_738),
    .Y(n_1074));
 AOI22xp5_ASAP7_75t_L g109910 (.A1(n_951),
    .A2(n_576),
    .B1(n_952),
    .B2(n_575),
    .Y(n_1073));
 XOR2xp5_ASAP7_75t_L g109911 (.A(n_8),
    .B(w2[1]),
    .Y(n_1072));
 OAI22xp5_ASAP7_75t_L g109912 (.A1(n_217),
    .A2(n_9001),
    .B1(n_8328),
    .B2(n_568),
    .Y(n_1071));
 OAI22xp5_ASAP7_75t_SL g109913 (.A1(n_1),
    .A2(n_573),
    .B1(n_923),
    .B2(n_574),
    .Y(n_1070));
 XOR2xp5_ASAP7_75t_SL g109914 (.A(n_704),
    .B(n_8318),
    .Y(n_1069));
 XOR2xp5_ASAP7_75t_SL g109915 (.A(n_5),
    .B(n_8304),
    .Y(n_1068));
 OAI22xp5_ASAP7_75t_L g109916 (.A1(n_8733),
    .A2(n_904),
    .B1(n_8732),
    .B2(n_903),
    .Y(n_1067));
 XNOR2xp5_ASAP7_75t_SL g109918 (.A(n_397),
    .B(n_720),
    .Y(n_1066));
 OAI22xp5_ASAP7_75t_SL g109919 (.A1(n_299),
    .A2(n_624),
    .B1(w2[4]),
    .B2(n_625),
    .Y(n_1065));
 XNOR2xp5_ASAP7_75t_L g109920 (.A(n_737),
    .B(n_8228),
    .Y(n_1064));
 XNOR2xp5_ASAP7_75t_L g109921 (.A(n_394),
    .B(n_757),
    .Y(n_1063));
 AOI22xp5_ASAP7_75t_SL g109922 (.A1(n_690),
    .A2(n_899),
    .B1(n_689),
    .B2(n_898),
    .Y(n_1062));
 XNOR2xp5_ASAP7_75t_SL g109923 (.A(n_424),
    .B(n_723),
    .Y(n_1141));
 INVx1_ASAP7_75t_L g109924 (.A(n_1060),
    .Y(n_1061));
 INVxp67_ASAP7_75t_L g109925 (.A(n_1058),
    .Y(n_1059));
 INVx1_ASAP7_75t_SL g109926 (.A(n_1056),
    .Y(n_1057));
 INVxp33_ASAP7_75t_R g109927 (.A(n_1055),
    .Y(n_1054));
 OAI22xp5_ASAP7_75t_SL g109928 (.A1(n_948),
    .A2(n_570),
    .B1(n_947),
    .B2(n_571),
    .Y(n_1053));
 AOI22xp5_ASAP7_75t_L g109930 (.A1(n_8748),
    .A2(n_0),
    .B1(n_8747),
    .B2(n_81),
    .Y(n_1060));
 XOR2xp5_ASAP7_75t_L g109931 (.A(n_721),
    .B(n_8310),
    .Y(n_1052));
 XNOR2xp5_ASAP7_75t_SL g109933 (.A(n_751),
    .B(n_8254),
    .Y(n_1051));
 OAI22xp5_ASAP7_75t_SL g109934 (.A1(n_8222),
    .A2(n_907),
    .B1(n_152),
    .B2(n_908),
    .Y(n_1050));
 OAI22xp5_ASAP7_75t_L g109935 (.A1(n_8625),
    .A2(n_613),
    .B1(n_8629),
    .B2(n_614),
    .Y(n_1049));
 OAI22xp5_ASAP7_75t_SL g109936 (.A1(n_209),
    .A2(n_13),
    .B1(n_8238),
    .B2(n_578),
    .Y(n_1048));
 AOI22xp5_ASAP7_75t_SL g109937 (.A1(n_941),
    .A2(n_641),
    .B1(n_942),
    .B2(n_640),
    .Y(n_1047));
 XNOR2xp5_ASAP7_75t_L g109938 (.A(n_735),
    .B(n_165),
    .Y(n_1046));
 XNOR2xp5_ASAP7_75t_SL g109939 (.A(n_434),
    .B(n_753),
    .Y(n_1045));
 XNOR2xp5_ASAP7_75t_L g109940 (.A(n_709),
    .B(n_8270),
    .Y(n_1044));
 OAI22xp5_ASAP7_75t_SL g109941 (.A1(n_946),
    .A2(n_86),
    .B1(n_3),
    .B2(n_85),
    .Y(n_1043));
 XOR2xp5_ASAP7_75t_R g109942 (.A(n_734),
    .B(n_8253),
    .Y(n_1042));
 XNOR2xp5_ASAP7_75t_SL g109943 (.A(n_711),
    .B(n_733),
    .Y(n_1041));
 XOR2xp5_ASAP7_75t_R g109944 (.A(n_8999),
    .B(n_8331),
    .Y(n_1040));
 XNOR2xp5_ASAP7_75t_SL g109945 (.A(n_435),
    .B(n_714),
    .Y(n_1039));
 AOI22xp5_ASAP7_75t_SL g109946 (.A1(n_692),
    .A2(n_902),
    .B1(n_691),
    .B2(n_901),
    .Y(n_1038));
 AOI22xp5_ASAP7_75t_L g109947 (.A1(n_8732),
    .A2(n_913),
    .B1(n_8733),
    .B2(n_914),
    .Y(n_1037));
 XNOR2xp5_ASAP7_75t_L g109948 (.A(n_4),
    .B(n_8229),
    .Y(n_1036));
 XOR2xp5_ASAP7_75t_SL g109949 (.A(n_11),
    .B(n_8329),
    .Y(n_1035));
 XNOR2xp5_ASAP7_75t_SL g109950 (.A(n_732),
    .B(n_581),
    .Y(n_1034));
 AOI22xp33_ASAP7_75t_L g109951 (.A1(n_59),
    .A2(n_968),
    .B1(n_200),
    .B2(n_969),
    .Y(n_1033));
 XNOR2xp5_ASAP7_75t_L g109952 (.A(n_731),
    .B(n_8329),
    .Y(n_1032));
 XNOR2xp5_ASAP7_75t_SL g109953 (.A(n_2),
    .B(n_436),
    .Y(n_1031));
 OAI22xp5_ASAP7_75t_L g109955 (.A1(n_270),
    .A2(n_610),
    .B1(w1[31]),
    .B2(n_609),
    .Y(n_1030));
 AOI22xp5_ASAP7_75t_L g109956 (.A1(n_945),
    .A2(n_83),
    .B1(n_944),
    .B2(n_84),
    .Y(n_1029));
 OAI22xp5_ASAP7_75t_L g109957 (.A1(n_956),
    .A2(n_77),
    .B1(n_955),
    .B2(n_76),
    .Y(n_1028));
 OAI22xp5_ASAP7_75t_SL g109958 (.A1(n_362),
    .A2(n_83),
    .B1(n_8334),
    .B2(n_84),
    .Y(n_1027));
 XNOR2xp5_ASAP7_75t_L g109959 (.A(n_722),
    .B(n_437),
    .Y(n_1058));
 OAI22xp5_ASAP7_75t_SL g109960 (.A1(n_593),
    .A2(n_931),
    .B1(n_932),
    .B2(n_594),
    .Y(n_1026));
 OAI22xp5_ASAP7_75t_L g109961 (.A1(n_8222),
    .A2(n_910),
    .B1(n_152),
    .B2(n_909),
    .Y(n_1025));
 XNOR2xp5_ASAP7_75t_L g109962 (.A(n_8998),
    .B(n_227),
    .Y(n_1024));
 AOI22xp5_ASAP7_75t_SL g109964 (.A1(w2[26]),
    .A2(n_893),
    .B1(n_264),
    .B2(n_892),
    .Y(n_1056));
 XNOR2xp5_ASAP7_75t_SL g109965 (.A(n_728),
    .B(n_419),
    .Y(n_1022));
 OAI22xp5_ASAP7_75t_SL g109966 (.A1(n_191),
    .A2(n_90),
    .B1(n_193),
    .B2(n_917),
    .Y(n_1021));
 OAI22xp5_ASAP7_75t_L g109967 (.A1(n_8792),
    .A2(n_589),
    .B1(n_8299),
    .B2(n_590),
    .Y(n_1020));
 OAI22xp5_ASAP7_75t_L g109968 (.A1(n_150),
    .A2(n_660),
    .B1(n_8323),
    .B2(n_659),
    .Y(n_1019));
 OAI22xp5_ASAP7_75t_SL g109969 (.A1(n_345),
    .A2(n_662),
    .B1(n_8302),
    .B2(n_661),
    .Y(n_1018));
 OAI22xp5_ASAP7_75t_L g109970 (.A1(n_196),
    .A2(n_643),
    .B1(n_8308),
    .B2(n_642),
    .Y(n_1017));
 OAI22xp5_ASAP7_75t_SL g109971 (.A1(n_184),
    .A2(n_601),
    .B1(n_8332),
    .B2(n_602),
    .Y(n_1016));
 OAI22xp5_ASAP7_75t_SL g109972 (.A1(n_645),
    .A2(n_571),
    .B1(n_644),
    .B2(n_570),
    .Y(n_1015));
 OAI22xp5_ASAP7_75t_SL g109973 (.A1(n_623),
    .A2(n_589),
    .B1(n_622),
    .B2(n_590),
    .Y(n_1014));
 XOR2xp5_ASAP7_75t_SL g109974 (.A(n_80),
    .B(n_661),
    .Y(n_1013));
 AOI22xp5_ASAP7_75t_SL g109975 (.A1(n_668),
    .A2(n_584),
    .B1(n_667),
    .B2(n_583),
    .Y(n_1012));
 AOI22xp5_ASAP7_75t_L g109976 (.A1(n_678),
    .A2(n_71),
    .B1(n_677),
    .B2(n_569),
    .Y(n_1011));
 OAI22xp5_ASAP7_75t_SL g109977 (.A1(n_348),
    .A2(n_573),
    .B1(n_8304),
    .B2(n_574),
    .Y(n_1010));
 OAI22xp5_ASAP7_75t_SL g109978 (.A1(n_8771),
    .A2(n_576),
    .B1(n_8770),
    .B2(n_575),
    .Y(n_1009));
 OAI22xp5_ASAP7_75t_SL g109979 (.A1(n_159),
    .A2(n_571),
    .B1(n_8310),
    .B2(n_570),
    .Y(n_1008));
 OAI22xp5_ASAP7_75t_SL g109980 (.A1(n_593),
    .A2(n_8771),
    .B1(n_8770),
    .B2(n_594),
    .Y(n_1007));
 AOI22xp5_ASAP7_75t_L g109981 (.A1(n_8310),
    .A2(n_645),
    .B1(n_159),
    .B2(n_644),
    .Y(n_1006));
 OAI22xp5_ASAP7_75t_L g109982 (.A1(n_676),
    .A2(n_607),
    .B1(n_675),
    .B2(n_608),
    .Y(n_1005));
 XNOR2xp5_ASAP7_75t_SL g109983 (.A(n_405),
    .B(n_8272),
    .Y(n_1004));
 OAI22xp5_ASAP7_75t_SL g109985 (.A1(n_8872),
    .A2(n_569),
    .B1(n_8881),
    .B2(n_71),
    .Y(n_1003));
 OAI22xp5_ASAP7_75t_SL g109986 (.A1(n_340),
    .A2(n_652),
    .B1(n_8337),
    .B2(n_653),
    .Y(n_1002));
 OAI22xp5_ASAP7_75t_SL g109987 (.A1(n_8923),
    .A2(n_650),
    .B1(n_8922),
    .B2(n_651),
    .Y(n_1001));
 AOI22xp5_ASAP7_75t_SL g109988 (.A1(n_8338),
    .A2(n_636),
    .B1(n_134),
    .B2(n_637),
    .Y(n_1000));
 OAI22xp5_ASAP7_75t_R g109989 (.A1(n_137),
    .A2(n_8),
    .B1(n_50),
    .B2(n_634),
    .Y(n_999));
 OAI22xp5_ASAP7_75t_SL g109990 (.A1(n_49),
    .A2(n_624),
    .B1(n_128),
    .B2(n_625),
    .Y(n_998));
 OAI22xp33_ASAP7_75t_R g109991 (.A1(n_125),
    .A2(n_81),
    .B1(n_8344),
    .B2(n_0),
    .Y(n_997));
 OAI22xp5_ASAP7_75t_L g109992 (.A1(n_47),
    .A2(n_613),
    .B1(n_48),
    .B2(n_614),
    .Y(n_996));
 XOR2xp5_ASAP7_75t_SL g109993 (.A(n_393),
    .B(n_606),
    .Y(n_995));
 OAI22xp5_ASAP7_75t_SL g109994 (.A1(n_8792),
    .A2(n_620),
    .B1(n_8299),
    .B2(n_621),
    .Y(n_994));
 OAI22xp33_ASAP7_75t_R g109995 (.A1(n_345),
    .A2(n_616),
    .B1(n_8302),
    .B2(n_80),
    .Y(n_993));
 OAI22xp5_ASAP7_75t_SL g109996 (.A1(n_191),
    .A2(n_631),
    .B1(n_193),
    .B2(n_630),
    .Y(n_992));
 OAI22xp5_ASAP7_75t_SL g109997 (.A1(n_627),
    .A2(n_196),
    .B1(n_8308),
    .B2(n_626),
    .Y(n_991));
 XOR2xp5_ASAP7_75t_SL g109998 (.A(n_418),
    .B(n_165),
    .Y(n_990));
 AOI22xp5_ASAP7_75t_SL g109999 (.A1(n_670),
    .A2(n_612),
    .B1(n_669),
    .B2(n_611),
    .Y(n_989));
 OAI22xp5_ASAP7_75t_SL g110000 (.A1(n_672),
    .A2(n_609),
    .B1(n_671),
    .B2(n_610),
    .Y(n_988));
 OAI22xp5_ASAP7_75t_SL g110001 (.A1(n_8282),
    .A2(n_565),
    .B1(n_163),
    .B2(n_566),
    .Y(n_987));
 AOI22xp5_ASAP7_75t_SL g110002 (.A1(n_591),
    .A2(n_647),
    .B1(n_592),
    .B2(n_646),
    .Y(n_986));
 OAI22xp5_ASAP7_75t_SL g110003 (.A1(n_8879),
    .A2(n_646),
    .B1(n_8877),
    .B2(n_647),
    .Y(n_985));
 OAI22xp5_ASAP7_75t_SL g110004 (.A1(n_682),
    .A2(n_654),
    .B1(n_681),
    .B2(n_655),
    .Y(n_984));
 XNOR2xp5_ASAP7_75t_SL g110005 (.A(n_408),
    .B(n_8254),
    .Y(n_983));
 XNOR2xp5_ASAP7_75t_L g110006 (.A(n_431),
    .B(n_8346),
    .Y(n_982));
 OAI22xp5_ASAP7_75t_SL g110007 (.A1(n_346),
    .A2(n_596),
    .B1(n_8327),
    .B2(n_595),
    .Y(n_981));
 AOI22xp5_ASAP7_75t_R g110008 (.A1(n_345),
    .A2(n_581),
    .B1(n_8302),
    .B2(n_582),
    .Y(n_980));
 AOI22xp5_ASAP7_75t_SL g110009 (.A1(n_191),
    .A2(n_72),
    .B1(n_193),
    .B2(n_73),
    .Y(n_979));
 AOI22xp5_ASAP7_75t_SL g110010 (.A1(n_619),
    .A2(n_8679),
    .B1(n_8245),
    .B2(n_618),
    .Y(n_978));
 OAI22xp5_ASAP7_75t_SL g110011 (.A1(n_46),
    .A2(n_596),
    .B1(n_45),
    .B2(n_595),
    .Y(n_977));
 OAI22xp5_ASAP7_75t_SL g110012 (.A1(n_145),
    .A2(n_633),
    .B1(n_144),
    .B2(n_632),
    .Y(n_976));
 AOI22xp5_ASAP7_75t_SL g110013 (.A1(n_330),
    .A2(n_649),
    .B1(n_8247),
    .B2(n_648),
    .Y(n_975));
 OAI211xp5_ASAP7_75t_R g110014 (.A1(dcnt[3]),
    .A2(n_921),
    .B(n_101),
    .C(rst),
    .Y(n_1055));
 NOR2xp33_ASAP7_75t_R g110079 (.A(n_112),
    .B(n_523),
    .Y(n_974));
 INVxp67_ASAP7_75t_L g110144 (.A(n_972),
    .Y(n_973));
 INVxp67_ASAP7_75t_L g110145 (.A(n_970),
    .Y(n_971));
 INVxp67_ASAP7_75t_R g110146 (.A(n_968),
    .Y(n_969));
 INVxp67_ASAP7_75t_R g110147 (.A(n_8995),
    .Y(n_967));
 INVxp67_ASAP7_75t_R g110148 (.A(n_964),
    .Y(n_965));
 INVxp67_ASAP7_75t_L g110149 (.A(n_962),
    .Y(n_963));
 INVx1_ASAP7_75t_SL g110151 (.A(n_959),
    .Y(n_960));
 INVxp67_ASAP7_75t_R g110152 (.A(n_8996),
    .Y(n_958));
 INVx1_ASAP7_75t_L g110153 (.A(n_955),
    .Y(n_956));
 INVx1_ASAP7_75t_L g110154 (.A(n_953),
    .Y(n_954));
 INVx1_ASAP7_75t_L g110155 (.A(n_951),
    .Y(n_952));
 INVxp67_ASAP7_75t_R g110156 (.A(n_8997),
    .Y(n_950));
 INVx1_ASAP7_75t_L g110157 (.A(n_947),
    .Y(n_948));
 INVxp67_ASAP7_75t_L g110158 (.A(n_3),
    .Y(n_946));
 INVx1_ASAP7_75t_L g110159 (.A(n_944),
    .Y(n_945));
 INVx1_ASAP7_75t_L g110161 (.A(n_941),
    .Y(n_942));
 INVxp67_ASAP7_75t_L g110162 (.A(n_939),
    .Y(n_940));
 INVxp67_ASAP7_75t_R g110163 (.A(n_937),
    .Y(n_938));
 INVxp67_ASAP7_75t_R g110166 (.A(n_933),
    .Y(n_934));
 INVx1_ASAP7_75t_SL g110167 (.A(n_931),
    .Y(n_932));
 INVxp67_ASAP7_75t_R g110168 (.A(n_929),
    .Y(n_930));
 INVxp67_ASAP7_75t_R g110169 (.A(n_7),
    .Y(n_928));
 INVx1_ASAP7_75t_L g110170 (.A(n_926),
    .Y(n_927));
 INVxp67_ASAP7_75t_L g110171 (.A(n_924),
    .Y(n_925));
 INVxp67_ASAP7_75t_R g110173 (.A(n_1),
    .Y(n_923));
 INVxp33_ASAP7_75t_R g110175 (.A(n_920),
    .Y(n_921));
 INVx1_ASAP7_75t_L g110176 (.A(n_918),
    .Y(n_919));
 INVx1_ASAP7_75t_SL g110178 (.A(n_90),
    .Y(n_917));
 INVx1_ASAP7_75t_SL g110181 (.A(n_916),
    .Y(n_915));
 INVx1_ASAP7_75t_L g110182 (.A(n_914),
    .Y(n_913));
 INVx1_ASAP7_75t_L g110187 (.A(n_909),
    .Y(n_910));
 INVx1_ASAP7_75t_SL g110189 (.A(n_908),
    .Y(n_907));
 INVx1_ASAP7_75t_L g110190 (.A(n_905),
    .Y(n_906));
 INVx1_ASAP7_75t_L g110191 (.A(n_904),
    .Y(n_903));
 INVx1_ASAP7_75t_L g110192 (.A(n_902),
    .Y(n_901));
 INVx1_ASAP7_75t_L g110193 (.A(n_899),
    .Y(n_898));
 INVx1_ASAP7_75t_SL g110194 (.A(n_897),
    .Y(n_896));
 INVx1_ASAP7_75t_SL g110195 (.A(n_894),
    .Y(n_895));
 INVx1_ASAP7_75t_SL g110196 (.A(n_892),
    .Y(n_893));
 INVx1_ASAP7_75t_R g110198 (.A(n_889),
    .Y(n_890));
 INVx1_ASAP7_75t_L g110201 (.A(n_85),
    .Y(n_86));
 INVx1_ASAP7_75t_SL g110204 (.A(n_84),
    .Y(n_83));
 AOI22xp33_ASAP7_75t_R g110205 (.A1(n_34),
    .A2(text_in_r[127]),
    .B1(text_in[127]),
    .B2(n_91),
    .Y(n_888));
 AOI21xp33_ASAP7_75t_R g110206 (.A1(dcnt[0]),
    .A2(dcnt[1]),
    .B(n_383),
    .Y(n_887));
 AOI22xp33_ASAP7_75t_R g110207 (.A1(n_35),
    .A2(text_in_r[38]),
    .B1(text_in[38]),
    .B2(n_92),
    .Y(n_886));
 AOI22xp33_ASAP7_75t_R g110208 (.A1(n_33),
    .A2(text_in_r[2]),
    .B1(text_in[2]),
    .B2(n_99),
    .Y(n_885));
 AOI22xp33_ASAP7_75t_R g110209 (.A1(n_97),
    .A2(text_in_r[126]),
    .B1(text_in[126]),
    .B2(n_92),
    .Y(n_884));
 AOI22xp33_ASAP7_75t_R g110210 (.A1(n_27),
    .A2(text_in_r[60]),
    .B1(text_in[60]),
    .B2(n_39),
    .Y(n_883));
 AOI22xp33_ASAP7_75t_R g110211 (.A1(n_27),
    .A2(text_in_r[29]),
    .B1(text_in[29]),
    .B2(n_94),
    .Y(n_882));
 AOI22xp33_ASAP7_75t_R g110212 (.A1(n_36),
    .A2(text_in_r[76]),
    .B1(text_in[76]),
    .B2(n_99),
    .Y(n_881));
 AOI22xp33_ASAP7_75t_R g110213 (.A1(n_97),
    .A2(text_in_r[98]),
    .B1(text_in[98]),
    .B2(n_92),
    .Y(n_880));
 AOI22xp33_ASAP7_75t_R g110214 (.A1(n_28),
    .A2(text_in_r[80]),
    .B1(text_in[80]),
    .B2(n_93),
    .Y(n_879));
 AOI22xp33_ASAP7_75t_R g110215 (.A1(n_96),
    .A2(text_in_r[28]),
    .B1(text_in[28]),
    .B2(n_100),
    .Y(n_878));
 AOI22xp33_ASAP7_75t_R g110216 (.A1(n_27),
    .A2(text_in_r[65]),
    .B1(text_in[65]),
    .B2(ld),
    .Y(n_877));
 AOI22xp33_ASAP7_75t_R g110217 (.A1(n_27),
    .A2(text_in_r[88]),
    .B1(text_in[88]),
    .B2(n_94),
    .Y(n_876));
 AOI22xp33_ASAP7_75t_R g110218 (.A1(n_97),
    .A2(text_in_r[24]),
    .B1(text_in[24]),
    .B2(n_92),
    .Y(n_875));
 AOI22xp33_ASAP7_75t_R g110219 (.A1(n_34),
    .A2(text_in_r[6]),
    .B1(text_in[6]),
    .B2(n_91),
    .Y(n_874));
 AOI22xp33_ASAP7_75t_R g110220 (.A1(n_33),
    .A2(text_in_r[122]),
    .B1(text_in[122]),
    .B2(n_100),
    .Y(n_873));
 AOI22xp33_ASAP7_75t_R g110221 (.A1(n_97),
    .A2(text_in_r[0]),
    .B1(text_in[0]),
    .B2(ld),
    .Y(n_872));
 AOI22xp33_ASAP7_75t_R g110222 (.A1(n_27),
    .A2(text_in_r[1]),
    .B1(text_in[1]),
    .B2(n_92),
    .Y(n_871));
 AOI22xp33_ASAP7_75t_R g110223 (.A1(n_34),
    .A2(text_in_r[3]),
    .B1(text_in[3]),
    .B2(n_39),
    .Y(n_870));
 AOI22xp33_ASAP7_75t_R g110224 (.A1(n_29),
    .A2(text_in_r[4]),
    .B1(text_in[4]),
    .B2(n_100),
    .Y(n_869));
 AOI22xp33_ASAP7_75t_R g110225 (.A1(n_33),
    .A2(text_in_r[5]),
    .B1(text_in[5]),
    .B2(n_91),
    .Y(n_868));
 AOI22xp33_ASAP7_75t_R g110226 (.A1(n_31),
    .A2(text_in_r[7]),
    .B1(text_in[7]),
    .B2(n_92),
    .Y(n_867));
 AOI22xp33_ASAP7_75t_R g110227 (.A1(n_32),
    .A2(text_in_r[8]),
    .B1(text_in[8]),
    .B2(n_100),
    .Y(n_866));
 AOI22xp33_ASAP7_75t_R g110228 (.A1(n_36),
    .A2(text_in_r[42]),
    .B1(text_in[42]),
    .B2(n_92),
    .Y(n_865));
 AOI22xp33_ASAP7_75t_R g110229 (.A1(n_35),
    .A2(text_in_r[9]),
    .B1(text_in[9]),
    .B2(n_91),
    .Y(n_864));
 AOI22xp33_ASAP7_75t_R g110230 (.A1(n_36),
    .A2(text_in_r[10]),
    .B1(text_in[10]),
    .B2(n_92),
    .Y(n_863));
 AOI22xp33_ASAP7_75t_R g110231 (.A1(n_101),
    .A2(text_in_r[11]),
    .B1(text_in[11]),
    .B2(n_94),
    .Y(n_862));
 AOI22xp33_ASAP7_75t_R g110232 (.A1(n_32),
    .A2(text_in_r[12]),
    .B1(text_in[12]),
    .B2(n_91),
    .Y(n_861));
 AOI22xp33_ASAP7_75t_R g110233 (.A1(n_101),
    .A2(text_in_r[13]),
    .B1(text_in[13]),
    .B2(n_100),
    .Y(n_860));
 AOI22xp33_ASAP7_75t_R g110234 (.A1(n_34),
    .A2(text_in_r[14]),
    .B1(text_in[14]),
    .B2(n_91),
    .Y(n_859));
 AOI22xp33_ASAP7_75t_R g110235 (.A1(n_33),
    .A2(text_in_r[15]),
    .B1(text_in[15]),
    .B2(n_91),
    .Y(n_858));
 AOI22xp33_ASAP7_75t_R g110236 (.A1(n_101),
    .A2(text_in_r[16]),
    .B1(text_in[16]),
    .B2(n_100),
    .Y(n_857));
 AOI22xp33_ASAP7_75t_R g110237 (.A1(n_101),
    .A2(text_in_r[17]),
    .B1(text_in[17]),
    .B2(n_100),
    .Y(n_856));
 AOI22xp33_ASAP7_75t_R g110238 (.A1(n_31),
    .A2(text_in_r[18]),
    .B1(text_in[18]),
    .B2(n_100),
    .Y(n_855));
 AOI22xp33_ASAP7_75t_R g110239 (.A1(n_32),
    .A2(text_in_r[19]),
    .B1(text_in[19]),
    .B2(n_92),
    .Y(n_854));
 AOI22xp33_ASAP7_75t_R g110240 (.A1(n_27),
    .A2(text_in_r[20]),
    .B1(text_in[20]),
    .B2(n_93),
    .Y(n_853));
 AOI22xp33_ASAP7_75t_R g110241 (.A1(n_101),
    .A2(text_in_r[21]),
    .B1(text_in[21]),
    .B2(n_39),
    .Y(n_852));
 AOI22xp33_ASAP7_75t_R g110242 (.A1(n_101),
    .A2(text_in_r[22]),
    .B1(text_in[22]),
    .B2(n_93),
    .Y(n_851));
 AOI22xp33_ASAP7_75t_R g110243 (.A1(n_96),
    .A2(text_in_r[23]),
    .B1(text_in[23]),
    .B2(n_93),
    .Y(n_850));
 AOI22xp33_ASAP7_75t_R g110244 (.A1(n_101),
    .A2(text_in_r[25]),
    .B1(text_in[25]),
    .B2(n_93),
    .Y(n_849));
 AOI22xp33_ASAP7_75t_R g110245 (.A1(n_28),
    .A2(text_in_r[26]),
    .B1(text_in[26]),
    .B2(n_98),
    .Y(n_848));
 AOI22xp33_ASAP7_75t_R g110246 (.A1(n_28),
    .A2(text_in_r[27]),
    .B1(text_in[27]),
    .B2(n_91),
    .Y(n_847));
 AOI22xp33_ASAP7_75t_R g110247 (.A1(n_96),
    .A2(text_in_r[116]),
    .B1(text_in[116]),
    .B2(n_91),
    .Y(n_846));
 AOI22xp33_ASAP7_75t_R g110248 (.A1(n_36),
    .A2(text_in_r[30]),
    .B1(text_in[30]),
    .B2(n_94),
    .Y(n_845));
 AOI22xp33_ASAP7_75t_R g110249 (.A1(n_97),
    .A2(text_in_r[31]),
    .B1(text_in[31]),
    .B2(n_92),
    .Y(n_844));
 AOI22xp33_ASAP7_75t_R g110250 (.A1(n_27),
    .A2(text_in_r[32]),
    .B1(text_in[32]),
    .B2(n_93),
    .Y(n_843));
 AOI22xp33_ASAP7_75t_R g110251 (.A1(n_28),
    .A2(text_in_r[33]),
    .B1(text_in[33]),
    .B2(n_93),
    .Y(n_842));
 AOI22xp33_ASAP7_75t_R g110252 (.A1(n_96),
    .A2(text_in_r[34]),
    .B1(text_in[34]),
    .B2(n_99),
    .Y(n_841));
 AOI22xp33_ASAP7_75t_R g110253 (.A1(n_30),
    .A2(text_in_r[35]),
    .B1(text_in[35]),
    .B2(n_100),
    .Y(n_840));
 AOI22xp33_ASAP7_75t_R g110254 (.A1(n_29),
    .A2(text_in_r[36]),
    .B1(text_in[36]),
    .B2(ld),
    .Y(n_839));
 AOI22xp33_ASAP7_75t_R g110255 (.A1(n_27),
    .A2(text_in_r[37]),
    .B1(text_in[37]),
    .B2(n_99),
    .Y(n_838));
 AOI22xp33_ASAP7_75t_R g110256 (.A1(n_97),
    .A2(text_in_r[39]),
    .B1(text_in[39]),
    .B2(n_91),
    .Y(n_837));
 AOI22xp33_ASAP7_75t_R g110257 (.A1(n_35),
    .A2(text_in_r[40]),
    .B1(text_in[40]),
    .B2(n_39),
    .Y(n_836));
 AOI22xp33_ASAP7_75t_R g110258 (.A1(n_96),
    .A2(text_in_r[41]),
    .B1(text_in[41]),
    .B2(n_91),
    .Y(n_835));
 AOI22xp33_ASAP7_75t_R g110259 (.A1(n_28),
    .A2(text_in_r[43]),
    .B1(text_in[43]),
    .B2(ld),
    .Y(n_834));
 AOI22xp33_ASAP7_75t_R g110260 (.A1(n_34),
    .A2(text_in_r[45]),
    .B1(text_in[45]),
    .B2(n_100),
    .Y(n_833));
 AOI22xp33_ASAP7_75t_R g110261 (.A1(n_33),
    .A2(text_in_r[46]),
    .B1(text_in[46]),
    .B2(n_94),
    .Y(n_832));
 AOI22xp33_ASAP7_75t_R g110262 (.A1(n_34),
    .A2(text_in_r[47]),
    .B1(text_in[47]),
    .B2(n_99),
    .Y(n_831));
 AOI22xp33_ASAP7_75t_R g110263 (.A1(n_33),
    .A2(text_in_r[48]),
    .B1(text_in[48]),
    .B2(n_99),
    .Y(n_830));
 AOI22xp33_ASAP7_75t_R g110264 (.A1(n_101),
    .A2(text_in_r[49]),
    .B1(text_in[49]),
    .B2(n_94),
    .Y(n_829));
 AOI22xp33_ASAP7_75t_R g110265 (.A1(n_27),
    .A2(text_in_r[50]),
    .B1(text_in[50]),
    .B2(n_93),
    .Y(n_828));
 AOI22xp33_ASAP7_75t_R g110266 (.A1(n_97),
    .A2(text_in_r[51]),
    .B1(text_in[51]),
    .B2(n_94),
    .Y(n_827));
 AOI22xp33_ASAP7_75t_R g110267 (.A1(n_30),
    .A2(text_in_r[52]),
    .B1(text_in[52]),
    .B2(n_98),
    .Y(n_826));
 AOI22xp33_ASAP7_75t_R g110268 (.A1(n_29),
    .A2(text_in_r[53]),
    .B1(text_in[53]),
    .B2(n_93),
    .Y(n_825));
 AOI22xp33_ASAP7_75t_R g110269 (.A1(n_30),
    .A2(text_in_r[54]),
    .B1(text_in[54]),
    .B2(n_94),
    .Y(n_824));
 AOI22xp33_ASAP7_75t_R g110270 (.A1(n_29),
    .A2(text_in_r[55]),
    .B1(text_in[55]),
    .B2(n_98),
    .Y(n_823));
 AOI22xp33_ASAP7_75t_R g110271 (.A1(n_97),
    .A2(text_in_r[56]),
    .B1(text_in[56]),
    .B2(n_99),
    .Y(n_822));
 AOI22xp33_ASAP7_75t_R g110272 (.A1(n_31),
    .A2(text_in_r[57]),
    .B1(text_in[57]),
    .B2(n_94),
    .Y(n_821));
 AOI22xp33_ASAP7_75t_R g110273 (.A1(n_32),
    .A2(text_in_r[58]),
    .B1(text_in[58]),
    .B2(n_39),
    .Y(n_820));
 AOI22xp33_ASAP7_75t_R g110274 (.A1(n_30),
    .A2(text_in_r[59]),
    .B1(text_in[59]),
    .B2(ld),
    .Y(n_819));
 AOI22xp33_ASAP7_75t_R g110275 (.A1(n_29),
    .A2(text_in_r[61]),
    .B1(text_in[61]),
    .B2(n_39),
    .Y(n_818));
 AOI22xp33_ASAP7_75t_R g110276 (.A1(n_35),
    .A2(text_in_r[62]),
    .B1(text_in[62]),
    .B2(n_92),
    .Y(n_817));
 AOI22xp33_ASAP7_75t_R g110277 (.A1(n_36),
    .A2(text_in_r[63]),
    .B1(text_in[63]),
    .B2(n_93),
    .Y(n_816));
 AOI22xp33_ASAP7_75t_R g110278 (.A1(n_35),
    .A2(text_in_r[64]),
    .B1(text_in[64]),
    .B2(n_100),
    .Y(n_815));
 AOI22xp33_ASAP7_75t_R g110279 (.A1(n_29),
    .A2(text_in_r[66]),
    .B1(text_in[66]),
    .B2(n_93),
    .Y(n_814));
 AOI22xp33_ASAP7_75t_R g110280 (.A1(n_34),
    .A2(text_in_r[67]),
    .B1(text_in[67]),
    .B2(n_100),
    .Y(n_813));
 AOI22xp33_ASAP7_75t_R g110281 (.A1(n_33),
    .A2(text_in_r[68]),
    .B1(text_in[68]),
    .B2(n_39),
    .Y(n_812));
 AOI22xp33_ASAP7_75t_R g110282 (.A1(n_35),
    .A2(text_in_r[69]),
    .B1(text_in[69]),
    .B2(n_92),
    .Y(n_811));
 AOI22xp33_ASAP7_75t_R g110283 (.A1(n_36),
    .A2(text_in_r[70]),
    .B1(text_in[70]),
    .B2(n_92),
    .Y(n_810));
 AOI22xp33_ASAP7_75t_R g110284 (.A1(n_34),
    .A2(text_in_r[71]),
    .B1(text_in[71]),
    .B2(ld),
    .Y(n_809));
 AOI22xp33_ASAP7_75t_R g110285 (.A1(n_33),
    .A2(text_in_r[72]),
    .B1(text_in[72]),
    .B2(n_99),
    .Y(n_808));
 AOI22xp33_ASAP7_75t_R g110286 (.A1(n_31),
    .A2(text_in_r[73]),
    .B1(text_in[73]),
    .B2(n_99),
    .Y(n_807));
 AOI22xp33_ASAP7_75t_R g110287 (.A1(n_31),
    .A2(text_in_r[74]),
    .B1(text_in[74]),
    .B2(n_94),
    .Y(n_806));
 AOI22xp33_ASAP7_75t_R g110288 (.A1(n_32),
    .A2(text_in_r[75]),
    .B1(text_in[75]),
    .B2(n_93),
    .Y(n_805));
 AOI22xp33_ASAP7_75t_R g110289 (.A1(n_30),
    .A2(text_in_r[77]),
    .B1(text_in[77]),
    .B2(n_99),
    .Y(n_804));
 AOI22xp33_ASAP7_75t_R g110290 (.A1(n_29),
    .A2(text_in_r[78]),
    .B1(text_in[78]),
    .B2(n_94),
    .Y(n_803));
 AOI22xp33_ASAP7_75t_R g110291 (.A1(n_35),
    .A2(text_in_r[79]),
    .B1(text_in[79]),
    .B2(n_91),
    .Y(n_802));
 AOI22xp33_ASAP7_75t_R g110292 (.A1(n_36),
    .A2(text_in_r[81]),
    .B1(text_in[81]),
    .B2(n_92),
    .Y(n_801));
 AOI22xp33_ASAP7_75t_R g110293 (.A1(n_35),
    .A2(text_in_r[82]),
    .B1(text_in[82]),
    .B2(n_92),
    .Y(n_800));
 AOI22xp33_ASAP7_75t_R g110294 (.A1(n_31),
    .A2(text_in_r[83]),
    .B1(text_in[83]),
    .B2(n_100),
    .Y(n_799));
 AOI22xp33_ASAP7_75t_R g110295 (.A1(n_32),
    .A2(text_in_r[84]),
    .B1(text_in[84]),
    .B2(n_39),
    .Y(n_798));
 AOI22xp33_ASAP7_75t_R g110296 (.A1(n_30),
    .A2(text_in_r[85]),
    .B1(text_in[85]),
    .B2(n_39),
    .Y(n_797));
 AOI22xp33_ASAP7_75t_R g110297 (.A1(n_29),
    .A2(text_in_r[86]),
    .B1(text_in[86]),
    .B2(n_94),
    .Y(n_796));
 AOI22xp33_ASAP7_75t_R g110298 (.A1(n_34),
    .A2(text_in_r[87]),
    .B1(text_in[87]),
    .B2(n_94),
    .Y(n_795));
 AOI22xp33_ASAP7_75t_R g110299 (.A1(n_33),
    .A2(text_in_r[89]),
    .B1(text_in[89]),
    .B2(n_94),
    .Y(n_794));
 AOI22xp33_ASAP7_75t_R g110300 (.A1(n_30),
    .A2(text_in_r[90]),
    .B1(text_in[90]),
    .B2(n_93),
    .Y(n_793));
 AOI22xp33_ASAP7_75t_R g110301 (.A1(n_27),
    .A2(text_in_r[44]),
    .B1(text_in[44]),
    .B2(n_94),
    .Y(n_792));
 AOI22xp33_ASAP7_75t_R g110302 (.A1(n_97),
    .A2(text_in_r[91]),
    .B1(text_in[91]),
    .B2(n_99),
    .Y(n_791));
 AOI22xp33_ASAP7_75t_R g110303 (.A1(n_97),
    .A2(text_in_r[92]),
    .B1(text_in[92]),
    .B2(n_98),
    .Y(n_790));
 AOI22xp33_ASAP7_75t_R g110304 (.A1(n_27),
    .A2(text_in_r[93]),
    .B1(text_in[93]),
    .B2(n_93),
    .Y(n_789));
 AOI22xp33_ASAP7_75t_R g110305 (.A1(n_96),
    .A2(text_in_r[94]),
    .B1(text_in[94]),
    .B2(ld),
    .Y(n_788));
 AOI22xp33_ASAP7_75t_R g110306 (.A1(n_28),
    .A2(text_in_r[95]),
    .B1(text_in[95]),
    .B2(n_98),
    .Y(n_787));
 AOI22xp33_ASAP7_75t_R g110307 (.A1(n_31),
    .A2(text_in_r[96]),
    .B1(text_in[96]),
    .B2(n_98),
    .Y(n_786));
 AOI22xp33_ASAP7_75t_R g110308 (.A1(n_32),
    .A2(text_in_r[97]),
    .B1(text_in[97]),
    .B2(n_39),
    .Y(n_785));
 AOI22xp33_ASAP7_75t_R g110309 (.A1(n_27),
    .A2(text_in_r[99]),
    .B1(text_in[99]),
    .B2(n_99),
    .Y(n_784));
 AOI22xp33_ASAP7_75t_R g110310 (.A1(n_97),
    .A2(text_in_r[100]),
    .B1(text_in[100]),
    .B2(n_100),
    .Y(n_783));
 AOI22xp33_ASAP7_75t_R g110311 (.A1(n_28),
    .A2(text_in_r[101]),
    .B1(text_in[101]),
    .B2(n_39),
    .Y(n_782));
 AOI22xp33_ASAP7_75t_R g110312 (.A1(n_96),
    .A2(text_in_r[102]),
    .B1(text_in[102]),
    .B2(n_91),
    .Y(n_781));
 AOI22xp33_ASAP7_75t_R g110313 (.A1(n_96),
    .A2(text_in_r[103]),
    .B1(text_in[103]),
    .B2(n_98),
    .Y(n_780));
 AOI22xp33_ASAP7_75t_R g110314 (.A1(n_28),
    .A2(text_in_r[104]),
    .B1(text_in[104]),
    .B2(n_93),
    .Y(n_779));
 AOI22xp33_ASAP7_75t_R g110315 (.A1(n_97),
    .A2(text_in_r[105]),
    .B1(text_in[105]),
    .B2(n_99),
    .Y(n_778));
 AOI22xp33_ASAP7_75t_R g110316 (.A1(n_28),
    .A2(text_in_r[106]),
    .B1(text_in[106]),
    .B2(n_39),
    .Y(n_777));
 AOI22xp33_ASAP7_75t_R g110317 (.A1(n_96),
    .A2(text_in_r[107]),
    .B1(text_in[107]),
    .B2(n_99),
    .Y(n_776));
 AOI22xp33_ASAP7_75t_R g110318 (.A1(n_31),
    .A2(text_in_r[108]),
    .B1(text_in[108]),
    .B2(n_98),
    .Y(n_775));
 AOI22xp33_ASAP7_75t_R g110319 (.A1(n_32),
    .A2(text_in_r[109]),
    .B1(text_in[109]),
    .B2(n_39),
    .Y(n_774));
 AOI22xp33_ASAP7_75t_R g110320 (.A1(n_35),
    .A2(text_in_r[110]),
    .B1(text_in[110]),
    .B2(n_39),
    .Y(n_773));
 AOI22xp33_ASAP7_75t_R g110321 (.A1(n_36),
    .A2(text_in_r[111]),
    .B1(text_in[111]),
    .B2(ld),
    .Y(n_772));
 AOI22xp33_ASAP7_75t_R g110322 (.A1(n_30),
    .A2(text_in_r[112]),
    .B1(text_in[112]),
    .B2(n_92),
    .Y(n_771));
 AOI22xp33_ASAP7_75t_R g110323 (.A1(n_28),
    .A2(text_in_r[113]),
    .B1(text_in[113]),
    .B2(n_99),
    .Y(n_770));
 AOI22xp33_ASAP7_75t_R g110324 (.A1(n_96),
    .A2(text_in_r[114]),
    .B1(text_in[114]),
    .B2(n_91),
    .Y(n_769));
 AOI22xp33_ASAP7_75t_R g110325 (.A1(n_31),
    .A2(text_in_r[115]),
    .B1(text_in[115]),
    .B2(n_91),
    .Y(n_768));
 AOI22xp33_ASAP7_75t_R g110326 (.A1(n_32),
    .A2(text_in_r[117]),
    .B1(text_in[117]),
    .B2(n_94),
    .Y(n_767));
 AOI22xp33_ASAP7_75t_R g110327 (.A1(n_96),
    .A2(text_in_r[118]),
    .B1(text_in[118]),
    .B2(n_91),
    .Y(n_766));
 AOI22xp33_ASAP7_75t_R g110328 (.A1(n_28),
    .A2(text_in_r[119]),
    .B1(text_in[119]),
    .B2(n_39),
    .Y(n_765));
 AOI22xp33_ASAP7_75t_R g110329 (.A1(n_36),
    .A2(text_in_r[121]),
    .B1(text_in[121]),
    .B2(n_39),
    .Y(n_764));
 AOI22xp33_ASAP7_75t_R g110330 (.A1(n_30),
    .A2(text_in_r[123]),
    .B1(text_in[123]),
    .B2(n_93),
    .Y(n_763));
 AOI22xp33_ASAP7_75t_R g110331 (.A1(n_29),
    .A2(text_in_r[124]),
    .B1(text_in[124]),
    .B2(n_100),
    .Y(n_762));
 AOI22xp33_ASAP7_75t_R g110332 (.A1(n_96),
    .A2(text_in_r[125]),
    .B1(text_in[125]),
    .B2(n_100),
    .Y(n_761));
 AOI22xp33_ASAP7_75t_R g110333 (.A1(n_28),
    .A2(text_in_r[120]),
    .B1(text_in[120]),
    .B2(n_99),
    .Y(n_760));
 AOI22xp5_ASAP7_75t_R g110334 (.A1(n_8833),
    .A2(n_116),
    .B1(n_114),
    .B2(n_8831),
    .Y(n_759));
 XNOR2xp5_ASAP7_75t_R g110335 (.A(n_8295),
    .B(w0[8]),
    .Y(n_758));
 OAI22xp33_ASAP7_75t_L g110336 (.A1(w2[6]),
    .A2(n_8264),
    .B1(n_259),
    .B2(n_164),
    .Y(n_757));
 OAI22xp33_ASAP7_75t_R g110337 (.A1(w0[11]),
    .A2(n_8231),
    .B1(n_313),
    .B2(n_186),
    .Y(n_756));
 AOI22xp5_ASAP7_75t_L g110338 (.A1(n_256),
    .A2(n_174),
    .B1(w0[24]),
    .B2(n_8287),
    .Y(n_972));
 AOI22xp5_ASAP7_75t_L g110340 (.A1(n_312),
    .A2(n_161),
    .B1(w0[15]),
    .B2(n_8275),
    .Y(n_970));
 XNOR2xp5_ASAP7_75t_R g110341 (.A(n_8296),
    .B(w1[8]),
    .Y(n_755));
 XNOR2xp5_ASAP7_75t_SL g110342 (.A(n_176),
    .B(w1[11]),
    .Y(n_754));
 AOI22xp5_ASAP7_75t_L g110343 (.A1(u0_n_32766),
    .A2(n_190),
    .B1(w3[6]),
    .B2(n_8266),
    .Y(n_753));
 AOI22xp5_ASAP7_75t_L g110344 (.A1(n_302),
    .A2(n_164),
    .B1(w2[21]),
    .B2(n_8264),
    .Y(n_968));
 XOR2xp5_ASAP7_75t_R g110346 (.A(n_69),
    .B(w2[8]),
    .Y(n_752));
 AOI22xp5_ASAP7_75t_SL g110349 (.A1(n_296),
    .A2(n_186),
    .B1(w0[27]),
    .B2(n_8231),
    .Y(n_964));
 OAI22xp5_ASAP7_75t_L g110350 (.A1(w1[21]),
    .A2(n_8262),
    .B1(n_252),
    .B2(n_143),
    .Y(n_751));
 XNOR2xp5_ASAP7_75t_SL g110351 (.A(n_51),
    .B(n_11401),
    .Y(n_962));
 OAI21xp33_ASAP7_75t_R g110352 (.A1(w3[30]),
    .A2(n_8274),
    .B(n_378),
    .Y(n_750));
 AOI22xp33_ASAP7_75t_SL g110353 (.A1(n_8884),
    .A2(u0_n_32749),
    .B1(n_11435),
    .B2(n_8234),
    .Y(n_961));
 XNOR2xp5_ASAP7_75t_R g110354 (.A(n_8295),
    .B(w0[16]),
    .Y(n_749));
 AOI22xp5_ASAP7_75t_L g110355 (.A1(u0_n_32714),
    .A2(n_138),
    .B1(w3[15]),
    .B2(n_8278),
    .Y(n_748));
 OAI22xp33_ASAP7_75t_R g110356 (.A1(w0[0]),
    .A2(n_8259),
    .B1(n_320),
    .B2(n_119),
    .Y(n_747));
 AOI22xp33_ASAP7_75t_R g110357 (.A1(n_247),
    .A2(n_186),
    .B1(w0[19]),
    .B2(n_8231),
    .Y(n_746));
 AOI22xp5_ASAP7_75t_L g110358 (.A1(n_300),
    .A2(n_179),
    .B1(w2[27]),
    .B2(n_178),
    .Y(n_959));
 XNOR2xp5_ASAP7_75t_R g110359 (.A(n_8260),
    .B(w0[6]),
    .Y(n_745));
 OAI21xp33_ASAP7_75t_R g110360 (.A1(w0[7]),
    .A2(n_8279),
    .B(n_381),
    .Y(n_744));
 XOR2xp5_ASAP7_75t_R g110362 (.A(n_8260),
    .B(w0[21]),
    .Y(n_743));
 AOI22xp33_ASAP7_75t_L g110363 (.A1(n_122),
    .A2(n_375),
    .B1(n_8243),
    .B2(n_8218),
    .Y(n_742));
 OAI21xp33_ASAP7_75t_R g110364 (.A1(w0[22]),
    .A2(n_8279),
    .B(n_377),
    .Y(n_741));
 XOR2xp5_ASAP7_75t_SL g110365 (.A(n_54),
    .B(w2[24]),
    .Y(n_955));
 OAI22xp5_ASAP7_75t_SL g110366 (.A1(w1[24]),
    .A2(n_37),
    .B1(n_291),
    .B2(n_167),
    .Y(n_953));
 OAI22xp33_ASAP7_75t_R g110367 (.A1(w0[23]),
    .A2(n_8259),
    .B1(n_278),
    .B2(n_119),
    .Y(n_740));
 AOI22xp5_ASAP7_75t_SL g110368 (.A1(n_368),
    .A2(n_42),
    .B1(w2[0]),
    .B2(n_44),
    .Y(n_951));
 OAI22xp5_ASAP7_75t_L g110369 (.A1(w1[6]),
    .A2(n_8262),
    .B1(n_271),
    .B2(n_143),
    .Y(n_739));
 XOR2xp5_ASAP7_75t_R g110371 (.A(n_8296),
    .B(w1[16]),
    .Y(n_738));
 XOR2xp5_ASAP7_75t_SL g110372 (.A(w1[19]),
    .B(n_176),
    .Y(n_737));
 OAI22xp5_ASAP7_75t_L g110373 (.A1(w2[7]),
    .A2(n_144),
    .B1(n_369),
    .B2(n_145),
    .Y(n_736));
 AOI22xp5_ASAP7_75t_L g110374 (.A1(n_321),
    .A2(n_116),
    .B1(w3[0]),
    .B2(n_114),
    .Y(n_947));
 OAI22xp5_ASAP7_75t_L g110375 (.A1(w1[22]),
    .A2(n_8280),
    .B1(n_316),
    .B2(n_8723),
    .Y(n_735));
 OAI22xp33_ASAP7_75t_R g110377 (.A1(w1[23]),
    .A2(n_8261),
    .B1(n_272),
    .B2(n_8933),
    .Y(n_734));
 AOI22xp5_ASAP7_75t_R g110378 (.A1(n_265),
    .A2(n_70),
    .B1(w2[16]),
    .B2(n_69),
    .Y(n_733));
 OAI22xp5_ASAP7_75t_SL g110379 (.A1(w3[16]),
    .A2(n_51),
    .B1(n_290),
    .B2(n_149),
    .Y(n_944));
 OAI22xp5_ASAP7_75t_SL g110380 (.A1(w1[30]),
    .A2(n_8272),
    .B1(u0_n_32676),
    .B2(n_199),
    .Y(n_732));
 AOI22xp33_ASAP7_75t_R g110381 (.A1(n_239),
    .A2(n_241),
    .B1(n_8317),
    .B2(n_8240),
    .Y(n_731));
 AOI22xp5_ASAP7_75t_L g110383 (.A1(n_322),
    .A2(n_42),
    .B1(w2[23]),
    .B2(n_44),
    .Y(n_943));
 OAI22xp5_ASAP7_75t_SL g110385 (.A1(w3[21]),
    .A2(n_8266),
    .B1(n_190),
    .B2(u0_n_32731),
    .Y(n_729));
 OAI22xp5_ASAP7_75t_L g110386 (.A1(w3[22]),
    .A2(n_8282),
    .B1(u0_n_33008),
    .B2(n_163),
    .Y(n_728));
 AOI22xp5_ASAP7_75t_L g110387 (.A1(n_361),
    .A2(n_150),
    .B1(n_8252),
    .B2(n_8323),
    .Y(n_727));
 OAI22xp5_ASAP7_75t_L g110388 (.A1(n_8236),
    .A2(n_8311),
    .B1(n_173),
    .B2(n_355),
    .Y(n_726));
 OAI22xp5_ASAP7_75t_L g110389 (.A1(n_8242),
    .A2(n_8320),
    .B1(n_349),
    .B2(n_350),
    .Y(n_725));
 OAI22xp5_ASAP7_75t_R g110390 (.A1(n_8258),
    .A2(n_8332),
    .B1(n_242),
    .B2(n_184),
    .Y(n_724));
 AOI22xp5_ASAP7_75t_SL g110391 (.A1(n_235),
    .A2(n_147),
    .B1(n_8300),
    .B2(n_8235),
    .Y(n_723));
 AOI22xp5_ASAP7_75t_L g110392 (.A1(w3[18]),
    .A2(n_166),
    .B1(u0_n_32741),
    .B2(n_8346),
    .Y(n_722));
 AOI22xp5_ASAP7_75t_L g110393 (.A1(n_349),
    .A2(n_196),
    .B1(n_8242),
    .B2(n_8308),
    .Y(n_941));
 OAI22xp5_ASAP7_75t_L g110394 (.A1(n_8236),
    .A2(n_8299),
    .B1(n_173),
    .B2(n_8792),
    .Y(n_939));
 OAI22xp5_ASAP7_75t_L g110395 (.A1(u0_n_32695),
    .A2(n_8309),
    .B1(w3[2]),
    .B2(n_182),
    .Y(n_721));
 XOR2xp5_ASAP7_75t_SL g110396 (.A(n_52),
    .B(w1[18]),
    .Y(n_720));
 AOI22xp5_ASAP7_75t_L g110397 (.A1(n_194),
    .A2(w0[30]),
    .B1(n_306),
    .B2(n_8279),
    .Y(n_937));
 OAI22xp5_ASAP7_75t_L g110398 (.A1(n_311),
    .A2(n_57),
    .B1(w0[3]),
    .B2(n_58),
    .Y(n_936));
 OAI22xp33_ASAP7_75t_R g110399 (.A1(n_8260),
    .A2(n_8922),
    .B1(n_148),
    .B2(n_8923),
    .Y(n_719));
 OAI22xp5_ASAP7_75t_L g110400 (.A1(u0_n_32685),
    .A2(n_8332),
    .B1(w3[13]),
    .B2(n_184),
    .Y(n_718));
 AOI22xp5_ASAP7_75t_L g110401 (.A1(n_164),
    .A2(n_49),
    .B1(n_8264),
    .B2(n_129),
    .Y(n_717));
 AOI22xp33_ASAP7_75t_R g110402 (.A1(n_190),
    .A2(n_47),
    .B1(n_8266),
    .B2(n_48),
    .Y(n_716));
 OAI22xp5_ASAP7_75t_L g110403 (.A1(n_303),
    .A2(n_8342),
    .B1(w2[10]),
    .B2(n_195),
    .Y(n_715));
 OAI22xp33_ASAP7_75t_R g110404 (.A1(u0_n_32687),
    .A2(n_8321),
    .B1(w3[26]),
    .B2(n_154),
    .Y(n_935));
 OAI22xp33_ASAP7_75t_R g110405 (.A1(n_289),
    .A2(n_8342),
    .B1(w2[18]),
    .B2(n_195),
    .Y(n_714));
 XOR2xp5_ASAP7_75t_R g110406 (.A(n_52),
    .B(w1[10]),
    .Y(n_713));
 OAI22xp33_ASAP7_75t_L g110407 (.A1(n_8262),
    .A2(n_8338),
    .B1(n_143),
    .B2(n_134),
    .Y(n_712));
 OAI22xp5_ASAP7_75t_L g110408 (.A1(n_365),
    .A2(n_8323),
    .B1(w0[13]),
    .B2(n_150),
    .Y(n_933));
 OAI22xp5_ASAP7_75t_R g110409 (.A1(n_8285),
    .A2(n_330),
    .B1(n_229),
    .B2(n_8247),
    .Y(n_711));
 OAI22xp5_ASAP7_75t_L g110410 (.A1(u0_n_33138),
    .A2(n_48),
    .B1(w3[20]),
    .B2(n_47),
    .Y(n_710));
 AOI22xp5_ASAP7_75t_L g110411 (.A1(w2[25]),
    .A2(n_136),
    .B1(n_258),
    .B2(n_8343),
    .Y(n_931));
 OAI22xp33_ASAP7_75t_R g110412 (.A1(n_328),
    .A2(n_8261),
    .B1(w1[15]),
    .B2(n_8933),
    .Y(n_929));
 OAI22xp5_ASAP7_75t_L g110413 (.A1(n_314),
    .A2(n_336),
    .B1(n_11346),
    .B2(n_337),
    .Y(n_709));
 XNOR2xp5_ASAP7_75t_L g110415 (.A(n_45),
    .B(w1[9]),
    .Y(n_708));
 OAI22xp5_ASAP7_75t_SL g110416 (.A1(n_309),
    .A2(n_8337),
    .B1(w0[25]),
    .B2(n_340),
    .Y(n_926));
 XOR2xp5_ASAP7_75t_R g110417 (.A(n_8254),
    .B(w1[14]),
    .Y(n_707));
 OAI22xp5_ASAP7_75t_SL g110418 (.A1(n_281),
    .A2(n_8344),
    .B1(w3[25]),
    .B2(n_125),
    .Y(n_924));
 OAI22xp5_ASAP7_75t_SL g110419 (.A1(n_253),
    .A2(n_8301),
    .B1(w0[26]),
    .B2(n_8872),
    .Y(n_706));
 AOI22xp5_ASAP7_75t_SL g110420 (.A1(n_8942),
    .A2(n_47),
    .B1(n_8946),
    .B2(n_8345),
    .Y(n_705));
 OAI22xp5_ASAP7_75t_SL g110422 (.A1(n_326),
    .A2(n_8343),
    .B1(w2[2]),
    .B2(n_136),
    .Y(n_704));
 AOI22xp5_ASAP7_75t_L g110423 (.A1(n_340),
    .A2(w0[2]),
    .B1(n_279),
    .B2(n_8337),
    .Y(n_703));
 OAI22xp33_ASAP7_75t_R g110424 (.A1(n_268),
    .A2(n_8335),
    .B1(w0[5]),
    .B2(n_8923),
    .Y(n_702));
 OAI22xp5_ASAP7_75t_L g110425 (.A1(n_260),
    .A2(n_8335),
    .B1(w0[20]),
    .B2(n_8923),
    .Y(n_701));
 AOI22xp33_ASAP7_75t_R g110426 (.A1(w1[2]),
    .A2(n_46),
    .B1(n_243),
    .B2(n_45),
    .Y(n_700));
 AOI22xp33_ASAP7_75t_R g110427 (.A1(n_134),
    .A2(w1[5]),
    .B1(n_298),
    .B2(n_8338),
    .Y(n_699));
 AOI22xp33_ASAP7_75t_R g110428 (.A1(n_8271),
    .A2(n_147),
    .B1(n_8235),
    .B2(n_364),
    .Y(n_698));
 OAI22xp33_ASAP7_75t_R g110431 (.A1(n_305),
    .A2(n_128),
    .B1(w2[5]),
    .B2(n_49),
    .Y(n_697));
 AOI22xp5_ASAP7_75t_L g110432 (.A1(w1[20]),
    .A2(n_134),
    .B1(n_269),
    .B2(n_8338),
    .Y(n_922));
 OAI22xp33_ASAP7_75t_R g110433 (.A1(u0_n_32691),
    .A2(n_48),
    .B1(w3[5]),
    .B2(n_47),
    .Y(n_696));
 OAI22xp5_ASAP7_75t_R g110434 (.A1(n_293),
    .A2(n_8338),
    .B1(w1[28]),
    .B2(n_134),
    .Y(n_695));
 AOI22xp5_ASAP7_75t_R g110437 (.A1(w3[17]),
    .A2(n_125),
    .B1(u0_n_32735),
    .B2(n_8344),
    .Y(n_693));
 NOR2xp33_ASAP7_75t_R g110438 (.A(dcnt[2]),
    .B(n_384),
    .Y(n_920));
 AOI22xp5_ASAP7_75t_SL g110439 (.A1(n_325),
    .A2(n_332),
    .B1(n_8324),
    .B2(n_7537),
    .Y(n_918));
 OAI22xp5_ASAP7_75t_SL g110440 (.A1(n_8225),
    .A2(n_330),
    .B1(n_218),
    .B2(n_8247),
    .Y(n_90));
 OAI22xp5_ASAP7_75t_SL g110441 (.A1(n_8342),
    .A2(n_8263),
    .B1(n_195),
    .B2(n_120),
    .Y(n_89));
 XNOR2x1_ASAP7_75t_L g110442 (.B(n_8339),
    .Y(n_916),
    .A(n_8261));
 AO22x1_ASAP7_75t_SL g110443 (.A1(n_330),
    .A2(n_187),
    .B1(n_8247),
    .B2(n_8318),
    .Y(n_914));
 OAI22xp5_ASAP7_75t_SL g110444 (.A1(n_8310),
    .A2(n_292),
    .B1(n_159),
    .B2(n_8322),
    .Y(n_912));
 XNOR2xp5_ASAP7_75t_SL g110445 (.A(n_68),
    .B(n_7447),
    .Y(n_88));
 AOI22xp5_ASAP7_75t_SL g110446 (.A1(n_346),
    .A2(n_8760),
    .B1(n_8253),
    .B2(n_8327),
    .Y(n_911));
 AOI22xp5_ASAP7_75t_L g110447 (.A1(n_154),
    .A2(n_338),
    .B1(n_8321),
    .B2(n_8249),
    .Y(n_909));
 OAI22xp5_ASAP7_75t_L g110448 (.A1(n_8255),
    .A2(n_8330),
    .B1(n_189),
    .B2(n_127),
    .Y(n_87));
 AOI22xp5_ASAP7_75t_SL g110449 (.A1(n_126),
    .A2(n_181),
    .B1(n_8241),
    .B2(n_8309),
    .Y(n_908));
 AO22x1_ASAP7_75t_SL g110450 (.A1(n_8271),
    .A2(n_161),
    .B1(n_364),
    .B2(n_8275),
    .Y(n_905));
 AO22x1_ASAP7_75t_SL g110451 (.A1(n_8785),
    .A2(n_53),
    .B1(n_8783),
    .B2(n_169),
    .Y(n_904));
 AOI22xp5_ASAP7_75t_SL g110452 (.A1(n_371),
    .A2(n_8302),
    .B1(n_8314),
    .B2(n_345),
    .Y(n_902));
 OAI22xp5_ASAP7_75t_SL g110453 (.A1(n_8336),
    .A2(n_8259),
    .B1(n_233),
    .B2(n_119),
    .Y(n_900));
 AO22x1_ASAP7_75t_SL g110454 (.A1(n_283),
    .A2(n_8304),
    .B1(n_8316),
    .B2(n_348),
    .Y(n_899));
 OAI22xp5_ASAP7_75t_SL g110455 (.A1(n_8312),
    .A2(n_8243),
    .B1(n_211),
    .B2(n_122),
    .Y(n_897));
 AOI22xp5_ASAP7_75t_SL g110456 (.A1(n_8678),
    .A2(n_232),
    .B1(n_8315),
    .B2(n_8245),
    .Y(n_894));
 OAI22x1_ASAP7_75t_SL g110457 (.A1(n_8319),
    .A2(n_8771),
    .B1(n_363),
    .B2(n_8307),
    .Y(n_892));
 AO22x1_ASAP7_75t_SL g110458 (.A1(n_166),
    .A2(n_113),
    .B1(n_8346),
    .B2(n_117),
    .Y(n_891));
 OA22x2_ASAP7_75t_L g110459 (.A1(n_8253),
    .A2(n_202),
    .B1(n_8228),
    .B2(n_8760),
    .Y(n_889));
 AOI22xp5_ASAP7_75t_SL g110460 (.A1(n_237),
    .A2(n_130),
    .B1(n_8303),
    .B2(n_131),
    .Y(n_85));
 OA21x2_ASAP7_75t_SL g110461 (.A1(n_360),
    .A2(n_7447),
    .B(n_376),
    .Y(n_84));
 INVxp67_ASAP7_75t_L g110462 (.A(n_691),
    .Y(n_692));
 INVxp67_ASAP7_75t_R g110463 (.A(n_689),
    .Y(n_690));
 INVxp67_ASAP7_75t_R g110464 (.A(n_687),
    .Y(n_688));
 INVxp67_ASAP7_75t_R g110465 (.A(n_685),
    .Y(n_686));
 INVxp67_ASAP7_75t_L g110466 (.A(n_683),
    .Y(n_684));
 INVxp67_ASAP7_75t_L g110467 (.A(n_681),
    .Y(n_682));
 INVx1_ASAP7_75t_L g110468 (.A(n_679),
    .Y(n_680));
 INVxp67_ASAP7_75t_L g110469 (.A(n_677),
    .Y(n_678));
 INVxp67_ASAP7_75t_R g110470 (.A(n_675),
    .Y(n_676));
 INVx1_ASAP7_75t_L g110471 (.A(n_673),
    .Y(n_674));
 INVx1_ASAP7_75t_SL g110472 (.A(n_671),
    .Y(n_672));
 INVxp67_ASAP7_75t_L g110473 (.A(n_669),
    .Y(n_670));
 INVxp67_ASAP7_75t_L g110474 (.A(n_667),
    .Y(n_668));
 INVx1_ASAP7_75t_L g110475 (.A(n_661),
    .Y(n_662));
 INVx2_ASAP7_75t_L g110476 (.A(n_660),
    .Y(n_659));
 INVxp67_ASAP7_75t_L g110477 (.A(n_657),
    .Y(n_658));
 INVxp67_ASAP7_75t_L g110478 (.A(n_656),
    .Y(n_657));
 INVx1_ASAP7_75t_SL g110479 (.A(n_655),
    .Y(n_654));
 INVx1_ASAP7_75t_L g110480 (.A(n_653),
    .Y(n_652));
 INVx1_ASAP7_75t_L g110481 (.A(n_651),
    .Y(n_650));
 INVx1_ASAP7_75t_SL g110482 (.A(n_648),
    .Y(n_649));
 INVx1_ASAP7_75t_L g110483 (.A(n_647),
    .Y(n_646));
 INVx1_ASAP7_75t_L g110485 (.A(n_644),
    .Y(n_645));
 INVxp67_ASAP7_75t_L g110486 (.A(n_643),
    .Y(n_642));
 INVx1_ASAP7_75t_L g110487 (.A(n_640),
    .Y(n_641));
 INVxp67_ASAP7_75t_SL g110488 (.A(n_638),
    .Y(n_639));
 INVx1_ASAP7_75t_SL g110490 (.A(n_637),
    .Y(n_636));
 INVxp33_ASAP7_75t_R g110493 (.A(n_8),
    .Y(n_634));
 INVx1_ASAP7_75t_L g110494 (.A(n_632),
    .Y(n_633));
 INVx1_ASAP7_75t_SL g110495 (.A(n_631),
    .Y(n_630));
 INVx1_ASAP7_75t_L g110497 (.A(n_626),
    .Y(n_627));
 INVx1_ASAP7_75t_SL g110498 (.A(n_625),
    .Y(n_624));
 INVxp67_ASAP7_75t_L g110499 (.A(n_622),
    .Y(n_623));
 HB1xp67_ASAP7_75t_SL g110500 (.A(n_620),
    .Y(n_622));
 INVx1_ASAP7_75t_L g110501 (.A(n_620),
    .Y(n_621));
 INVx1_ASAP7_75t_SL g110503 (.A(n_0),
    .Y(n_81));
 INVx2_ASAP7_75t_SL g110505 (.A(n_618),
    .Y(n_619));
 INVxp67_ASAP7_75t_R g110508 (.A(n_80),
    .Y(n_616));
 INVx1_ASAP7_75t_L g110509 (.A(n_614),
    .Y(n_613));
 INVx1_ASAP7_75t_SL g110512 (.A(n_78),
    .Y(n_79));
 INVx1_ASAP7_75t_SL g110513 (.A(n_611),
    .Y(n_612));
 INVx1_ASAP7_75t_L g110514 (.A(n_610),
    .Y(n_609));
 INVx1_ASAP7_75t_SL g110515 (.A(n_608),
    .Y(n_607));
 INVx1_ASAP7_75t_SL g110520 (.A(n_76),
    .Y(n_77));
 INVx1_ASAP7_75t_SL g110521 (.A(n_603),
    .Y(n_604));
 INVxp67_ASAP7_75t_L g110522 (.A(n_601),
    .Y(n_602));
 INVx1_ASAP7_75t_SL g110524 (.A(n_9000),
    .Y(n_599));
 INVx1_ASAP7_75t_SL g110525 (.A(n_598),
    .Y(n_597));
 INVx1_ASAP7_75t_SL g110526 (.A(n_596),
    .Y(n_595));
 INVx2_ASAP7_75t_L g110527 (.A(n_594),
    .Y(n_593));
 INVx1_ASAP7_75t_L g110528 (.A(n_591),
    .Y(n_592));
 INVx1_ASAP7_75t_L g110529 (.A(n_590),
    .Y(n_589));
 INVxp67_ASAP7_75t_SL g110531 (.A(n_587),
    .Y(n_588));
 INVx1_ASAP7_75t_L g110532 (.A(n_585),
    .Y(n_586));
 INVx1_ASAP7_75t_SL g110533 (.A(n_584),
    .Y(n_583));
 INVx1_ASAP7_75t_SL g110535 (.A(n_581),
    .Y(n_582));
 INVx1_ASAP7_75t_SL g110538 (.A(n_13),
    .Y(n_578));
 INVx1_ASAP7_75t_SL g110539 (.A(n_10),
    .Y(n_577));
 INVx1_ASAP7_75t_L g110541 (.A(n_72),
    .Y(n_73));
 INVx1_ASAP7_75t_SL g110543 (.A(n_576),
    .Y(n_575));
 INVx2_ASAP7_75t_L g110544 (.A(n_574),
    .Y(n_573));
 INVx1_ASAP7_75t_L g110545 (.A(n_571),
    .Y(n_570));
 INVx1_ASAP7_75t_SL g110547 (.A(n_71),
    .Y(n_569));
 INVx1_ASAP7_75t_L g110549 (.A(n_9001),
    .Y(n_568));
 INVx1_ASAP7_75t_L g110550 (.A(n_565),
    .Y(n_566));
 XNOR2xp5_ASAP7_75t_R g110553 (.A(w0[15]),
    .B(text_in_r[111]),
    .Y(n_564));
 XOR2xp5_ASAP7_75t_R g110554 (.A(n_265),
    .B(text_in_r[48]),
    .Y(n_563));
 XNOR2xp5_ASAP7_75t_R g110555 (.A(text_in_r[7]),
    .B(w3[7]),
    .Y(n_562));
 XNOR2xp5_ASAP7_75t_R g110556 (.A(text_in_r[22]),
    .B(w3[22]),
    .Y(n_561));
 XNOR2xp5_ASAP7_75t_R g110557 (.A(w1[23]),
    .B(text_in_r[87]),
    .Y(n_560));
 XNOR2xp5_ASAP7_75t_R g110558 (.A(w3[5]),
    .B(text_in_r[5]),
    .Y(n_559));
 XOR2xp5_ASAP7_75t_R g110559 (.A(n_316),
    .B(text_in_r[86]),
    .Y(n_558));
 XNOR2xp5_ASAP7_75t_R g110560 (.A(w3[21]),
    .B(text_in_r[21]),
    .Y(n_557));
 XOR2xp5_ASAP7_75t_R g110561 (.A(n_264),
    .B(text_in_r[58]),
    .Y(n_556));
 XNOR2xp5_ASAP7_75t_R g110562 (.A(text_in_r[20]),
    .B(w3[20]),
    .Y(n_555));
 XNOR2xp5_ASAP7_75t_R g110563 (.A(text_in_r[3]),
    .B(w3[3]),
    .Y(n_554));
 XNOR2xp5_ASAP7_75t_R g110564 (.A(text_in_r[19]),
    .B(n_8668),
    .Y(n_553));
 XNOR2xp5_ASAP7_75t_R g110565 (.A(w1[21]),
    .B(text_in_r[85]),
    .Y(n_552));
 XOR2xp5_ASAP7_75t_R g110566 (.A(u0_n_32741),
    .B(text_in_r[18]),
    .Y(n_551));
 XNOR2xp5_ASAP7_75t_R g110567 (.A(w1[27]),
    .B(text_in_r[91]),
    .Y(n_550));
 XOR2xp5_ASAP7_75t_R g110568 (.A(u0_n_32695),
    .B(text_in_r[2]),
    .Y(n_549));
 XNOR2xp5_ASAP7_75t_R g110569 (.A(text_in_r[1]),
    .B(n_8748),
    .Y(n_548));
 XNOR2xp5_ASAP7_75t_R g110570 (.A(w3[0]),
    .B(text_in_r[0]),
    .Y(n_547));
 XNOR2xp5_ASAP7_75t_R g110571 (.A(w2[7]),
    .B(text_in_r[39]),
    .Y(n_546));
 XNOR2xp5_ASAP7_75t_R g110572 (.A(w1[20]),
    .B(text_in_r[84]),
    .Y(n_545));
 XNOR2xp5_ASAP7_75t_R g110573 (.A(w1[26]),
    .B(text_in_r[90]),
    .Y(n_544));
 XNOR2xp5_ASAP7_75t_R g110574 (.A(w2[6]),
    .B(text_in_r[38]),
    .Y(n_543));
 XNOR2xp5_ASAP7_75t_R g110575 (.A(w1[19]),
    .B(text_in_r[83]),
    .Y(n_542));
 XOR2xp5_ASAP7_75t_R g110576 (.A(n_305),
    .B(text_in_r[37]),
    .Y(n_541));
 XNOR2xp5_ASAP7_75t_R g110577 (.A(w2[4]),
    .B(text_in_r[36]),
    .Y(n_540));
 XNOR2xp5_ASAP7_75t_R g110578 (.A(w2[0]),
    .B(text_in_r[32]),
    .Y(n_539));
 XNOR2xp5_ASAP7_75t_R g110579 (.A(w2[3]),
    .B(text_in_r[35]),
    .Y(n_538));
 XNOR2xp5_ASAP7_75t_R g110580 (.A(w2[2]),
    .B(text_in_r[34]),
    .Y(n_537));
 XNOR2xp5_ASAP7_75t_R g110581 (.A(w1[17]),
    .B(text_in_r[81]),
    .Y(n_536));
 XNOR2xp5_ASAP7_75t_R g110582 (.A(w2[1]),
    .B(text_in_r[33]),
    .Y(n_535));
 XNOR2xp5_ASAP7_75t_R g110583 (.A(w1[25]),
    .B(text_in_r[89]),
    .Y(n_534));
 XNOR2xp5_ASAP7_75t_R g110584 (.A(w0[21]),
    .B(text_in_r[117]),
    .Y(n_533));
 XNOR2xp5_ASAP7_75t_R g110585 (.A(w1[16]),
    .B(text_in_r[80]),
    .Y(n_532));
 XNOR2xp5_ASAP7_75t_R g110586 (.A(w1[7]),
    .B(text_in_r[71]),
    .Y(n_531));
 XOR2xp5_ASAP7_75t_R g110587 (.A(n_271),
    .B(text_in_r[70]),
    .Y(n_530));
 XNOR2xp5_ASAP7_75t_R g110588 (.A(text_in_r[4]),
    .B(n_8629),
    .Y(n_529));
 XNOR2xp5_ASAP7_75t_R g110589 (.A(w0[23]),
    .B(text_in_r[119]),
    .Y(n_528));
 XNOR2xp5_ASAP7_75t_R g110590 (.A(w1[5]),
    .B(text_in_r[69]),
    .Y(n_527));
 XNOR2xp5_ASAP7_75t_R g110591 (.A(w1[24]),
    .B(text_in_r[88]),
    .Y(n_526));
 XNOR2xp5_ASAP7_75t_R g110592 (.A(w1[3]),
    .B(text_in_r[67]),
    .Y(n_525));
 XNOR2xp5_ASAP7_75t_R g110593 (.A(w0[22]),
    .B(text_in_r[118]),
    .Y(n_524));
 XNOR2xp5_ASAP7_75t_R g110594 (.A(w1[2]),
    .B(text_in_r[66]),
    .Y(n_523));
 XNOR2xp5_ASAP7_75t_R g110595 (.A(w1[1]),
    .B(text_in_r[65]),
    .Y(n_522));
 XNOR2xp5_ASAP7_75t_R g110596 (.A(w1[0]),
    .B(text_in_r[64]),
    .Y(n_521));
 XNOR2xp5_ASAP7_75t_R g110597 (.A(w0[31]),
    .B(text_in_r[127]),
    .Y(n_520));
 XNOR2xp5_ASAP7_75t_R g110598 (.A(w0[7]),
    .B(text_in_r[103]),
    .Y(n_519));
 XNOR2xp5_ASAP7_75t_R g110599 (.A(w2[17]),
    .B(text_in_r[49]),
    .Y(n_518));
 XNOR2xp5_ASAP7_75t_R g110600 (.A(w0[6]),
    .B(text_in_r[102]),
    .Y(n_517));
 XNOR2xp5_ASAP7_75t_R g110601 (.A(w0[20]),
    .B(text_in_r[116]),
    .Y(n_516));
 XNOR2xp5_ASAP7_75t_R g110602 (.A(w0[5]),
    .B(text_in_r[101]),
    .Y(n_515));
 XNOR2xp5_ASAP7_75t_R g110603 (.A(w0[4]),
    .B(text_in_r[100]),
    .Y(n_514));
 XNOR2xp5_ASAP7_75t_R g110604 (.A(w2[21]),
    .B(text_in_r[53]),
    .Y(n_513));
 XNOR2xp5_ASAP7_75t_R g110605 (.A(w0[30]),
    .B(text_in_r[126]),
    .Y(n_512));
 XNOR2xp5_ASAP7_75t_R g110606 (.A(w0[19]),
    .B(text_in_r[115]),
    .Y(n_511));
 XNOR2xp5_ASAP7_75t_R g110607 (.A(w0[17]),
    .B(text_in_r[113]),
    .Y(n_510));
 XNOR2xp5_ASAP7_75t_R g110608 (.A(w1[4]),
    .B(text_in_r[68]),
    .Y(n_509));
 XNOR2xp5_ASAP7_75t_R g110609 (.A(w0[1]),
    .B(text_in_r[97]),
    .Y(n_508));
 XNOR2xp5_ASAP7_75t_R g110610 (.A(text_in_r[17]),
    .B(w3[17]),
    .Y(n_507));
 XNOR2xp5_ASAP7_75t_R g110611 (.A(w0[0]),
    .B(text_in_r[96]),
    .Y(n_506));
 XNOR2xp5_ASAP7_75t_R g110612 (.A(text_in_r[15]),
    .B(w3[15]),
    .Y(n_505));
 XNOR2xp5_ASAP7_75t_R g110613 (.A(w0[16]),
    .B(text_in_r[112]),
    .Y(n_504));
 XNOR2xp5_ASAP7_75t_R g110614 (.A(w0[29]),
    .B(text_in_r[125]),
    .Y(n_503));
 XNOR2xp5_ASAP7_75t_R g110615 (.A(w3[13]),
    .B(text_in_r[13]),
    .Y(n_502));
 XNOR2xp5_ASAP7_75t_R g110616 (.A(w2[23]),
    .B(text_in_r[55]),
    .Y(n_501));
 XNOR2xp5_ASAP7_75t_R g110617 (.A(w1[31]),
    .B(text_in_r[95]),
    .Y(n_500));
 XNOR2xp5_ASAP7_75t_R g110618 (.A(w2[18]),
    .B(text_in_r[50]),
    .Y(n_499));
 XNOR2xp5_ASAP7_75t_R g110619 (.A(w1[30]),
    .B(text_in_r[94]),
    .Y(n_498));
 XNOR2xp5_ASAP7_75t_R g110620 (.A(text_in_r[12]),
    .B(w3[12]),
    .Y(n_497));
 XNOR2xp5_ASAP7_75t_R g110621 (.A(w2[20]),
    .B(text_in_r[52]),
    .Y(n_496));
 XNOR2xp5_ASAP7_75t_R g110622 (.A(text_in_r[31]),
    .B(w3[31]),
    .Y(n_495));
 XNOR2xp5_ASAP7_75t_R g110623 (.A(w2[19]),
    .B(text_in_r[51]),
    .Y(n_494));
 XNOR2xp5_ASAP7_75t_R g110624 (.A(w1[29]),
    .B(text_in_r[93]),
    .Y(n_493));
 XNOR2xp5_ASAP7_75t_R g110625 (.A(w0[2]),
    .B(text_in_r[98]),
    .Y(n_492));
 XNOR2xp5_ASAP7_75t_R g110626 (.A(w3[11]),
    .B(text_in_r[11]),
    .Y(n_491));
 XNOR2xp5_ASAP7_75t_R g110627 (.A(w3[10]),
    .B(text_in_r[10]),
    .Y(n_490));
 XNOR2xp5_ASAP7_75t_R g110628 (.A(w3[30]),
    .B(text_in_r[30]),
    .Y(n_489));
 XNOR2xp5_ASAP7_75t_R g110629 (.A(w1[18]),
    .B(text_in_r[82]),
    .Y(n_488));
 XNOR2xp5_ASAP7_75t_R g110630 (.A(w0[28]),
    .B(text_in_r[124]),
    .Y(n_487));
 XNOR2xp5_ASAP7_75t_R g110631 (.A(text_in_r[9]),
    .B(n_8856),
    .Y(n_486));
 XNOR2xp5_ASAP7_75t_R g110632 (.A(n_11401),
    .B(text_in_r[8]),
    .Y(n_485));
 XNOR2xp5_ASAP7_75t_R g110633 (.A(w3[29]),
    .B(text_in_r[29]),
    .Y(n_484));
 XNOR2xp5_ASAP7_75t_R g110634 (.A(w2[15]),
    .B(text_in_r[47]),
    .Y(n_483));
 XNOR2xp5_ASAP7_75t_R g110635 (.A(w2[14]),
    .B(text_in_r[46]),
    .Y(n_482));
 XNOR2xp5_ASAP7_75t_R g110636 (.A(w2[13]),
    .B(text_in_r[45]),
    .Y(n_481));
 XNOR2xp5_ASAP7_75t_R g110637 (.A(text_in_r[23]),
    .B(n_8831),
    .Y(n_480));
 XNOR2xp5_ASAP7_75t_R g110638 (.A(w0[8]),
    .B(text_in_r[104]),
    .Y(n_479));
 XNOR2xp5_ASAP7_75t_R g110639 (.A(w2[28]),
    .B(text_in_r[60]),
    .Y(n_478));
 XNOR2xp5_ASAP7_75t_R g110640 (.A(w0[9]),
    .B(text_in_r[105]),
    .Y(n_477));
 XNOR2xp5_ASAP7_75t_R g110641 (.A(w0[10]),
    .B(text_in_r[106]),
    .Y(n_476));
 XNOR2xp5_ASAP7_75t_R g110642 (.A(w0[3]),
    .B(text_in_r[99]),
    .Y(n_475));
 XNOR2xp5_ASAP7_75t_R g110643 (.A(w0[11]),
    .B(text_in_r[107]),
    .Y(n_474));
 XNOR2xp5_ASAP7_75t_R g110644 (.A(w2[29]),
    .B(text_in_r[61]),
    .Y(n_473));
 XNOR2xp5_ASAP7_75t_R g110645 (.A(w0[12]),
    .B(text_in_r[108]),
    .Y(n_472));
 XNOR2xp5_ASAP7_75t_R g110646 (.A(w0[13]),
    .B(text_in_r[109]),
    .Y(n_471));
 XNOR2xp5_ASAP7_75t_R g110647 (.A(w0[24]),
    .B(text_in_r[120]),
    .Y(n_470));
 XNOR2xp5_ASAP7_75t_R g110648 (.A(w2[30]),
    .B(text_in_r[62]),
    .Y(n_469));
 XNOR2xp5_ASAP7_75t_R g110649 (.A(w2[27]),
    .B(text_in_r[59]),
    .Y(n_468));
 XNOR2xp5_ASAP7_75t_R g110650 (.A(w2[24]),
    .B(text_in_r[56]),
    .Y(n_467));
 XNOR2xp5_ASAP7_75t_R g110651 (.A(w1[8]),
    .B(text_in_r[72]),
    .Y(n_466));
 XOR2xp5_ASAP7_75t_R g110652 (.A(u0_n_32766),
    .B(text_in_r[6]),
    .Y(n_465));
 XNOR2xp5_ASAP7_75t_R g110653 (.A(w2[31]),
    .B(text_in_r[63]),
    .Y(n_464));
 XNOR2xp5_ASAP7_75t_R g110654 (.A(w1[9]),
    .B(text_in_r[73]),
    .Y(n_463));
 XNOR2xp5_ASAP7_75t_R g110655 (.A(w0[25]),
    .B(text_in_r[121]),
    .Y(n_462));
 XNOR2xp5_ASAP7_75t_R g110656 (.A(w1[10]),
    .B(text_in_r[74]),
    .Y(n_461));
 XNOR2xp5_ASAP7_75t_R g110657 (.A(w1[11]),
    .B(text_in_r[75]),
    .Y(n_460));
 XNOR2xp5_ASAP7_75t_R g110658 (.A(w2[22]),
    .B(text_in_r[54]),
    .Y(n_459));
 XNOR2xp5_ASAP7_75t_R g110659 (.A(w3[24]),
    .B(text_in_r[24]),
    .Y(n_458));
 XOR2xp5_ASAP7_75t_R g110660 (.A(n_290),
    .B(text_in_r[16]),
    .Y(n_457));
 XNOR2xp5_ASAP7_75t_R g110661 (.A(w1[12]),
    .B(text_in_r[76]),
    .Y(n_456));
 XNOR2xp5_ASAP7_75t_R g110662 (.A(w2[25]),
    .B(text_in_r[57]),
    .Y(n_455));
 XNOR2xp5_ASAP7_75t_R g110663 (.A(text_in_r[25]),
    .B(w3[25]),
    .Y(n_454));
 XNOR2xp5_ASAP7_75t_R g110664 (.A(w1[13]),
    .B(text_in_r[77]),
    .Y(n_453));
 XNOR2xp5_ASAP7_75t_R g110665 (.A(w1[14]),
    .B(text_in_r[78]),
    .Y(n_452));
 XOR2xp5_ASAP7_75t_R g110666 (.A(n_253),
    .B(text_in_r[122]),
    .Y(n_451));
 XNOR2xp5_ASAP7_75t_R g110667 (.A(w1[15]),
    .B(text_in_r[79]),
    .Y(n_450));
 XNOR2xp5_ASAP7_75t_R g110668 (.A(w1[28]),
    .B(text_in_r[92]),
    .Y(n_449));
 XNOR2xp5_ASAP7_75t_R g110669 (.A(w3[26]),
    .B(text_in_r[26]),
    .Y(n_448));
 XNOR2xp5_ASAP7_75t_R g110670 (.A(w2[8]),
    .B(text_in_r[40]),
    .Y(n_447));
 XNOR2xp5_ASAP7_75t_R g110671 (.A(w2[9]),
    .B(text_in_r[41]),
    .Y(n_446));
 XNOR2xp5_ASAP7_75t_R g110672 (.A(w2[10]),
    .B(text_in_r[42]),
    .Y(n_445));
 XNOR2xp5_ASAP7_75t_R g110673 (.A(w3[27]),
    .B(text_in_r[27]),
    .Y(n_444));
 XNOR2xp5_ASAP7_75t_R g110674 (.A(w2[11]),
    .B(text_in_r[43]),
    .Y(n_443));
 XNOR2xp5_ASAP7_75t_R g110675 (.A(w0[27]),
    .B(text_in_r[123]),
    .Y(n_442));
 XNOR2xp5_ASAP7_75t_R g110676 (.A(w2[12]),
    .B(text_in_r[44]),
    .Y(n_441));
 XNOR2xp5_ASAP7_75t_R g110677 (.A(text_in_r[28]),
    .B(n_8942),
    .Y(n_440));
 OAI22xp33_ASAP7_75t_R g110678 (.A1(n_69),
    .A2(n_60),
    .B1(n_224),
    .B2(n_70),
    .Y(n_439));
 OAI22xp33_ASAP7_75t_R g110679 (.A1(n_8342),
    .A2(n_189),
    .B1(n_8330),
    .B2(n_195),
    .Y(n_438));
 OAI22xp5_ASAP7_75t_L g110680 (.A1(n_183),
    .A2(n_68),
    .B1(n_67),
    .B2(n_180),
    .Y(n_437));
 OAI22xp5_ASAP7_75t_L g110681 (.A1(n_8256),
    .A2(n_341),
    .B1(n_59),
    .B2(n_8277),
    .Y(n_436));
 OAI22xp5_ASAP7_75t_SL g110682 (.A1(n_189),
    .A2(n_169),
    .B1(n_53),
    .B2(n_8330),
    .Y(n_435));
 AOI22xp5_ASAP7_75t_R g110683 (.A1(n_8242),
    .A2(n_158),
    .B1(n_349),
    .B2(n_8270),
    .Y(n_434));
 OAI22xp33_ASAP7_75t_R g110684 (.A1(n_67),
    .A2(n_154),
    .B1(n_68),
    .B2(n_8321),
    .Y(n_433));
 OAI22xp33_ASAP7_75t_R g110685 (.A1(n_8770),
    .A2(n_53),
    .B1(n_169),
    .B2(n_8771),
    .Y(n_432));
 AOI22xp5_ASAP7_75t_L g110686 (.A1(n_8321),
    .A2(n_180),
    .B1(n_183),
    .B2(n_154),
    .Y(n_431));
 OAI22xp33_ASAP7_75t_R g110687 (.A1(n_68),
    .A2(n_8346),
    .B1(n_67),
    .B2(n_166),
    .Y(n_430));
 OAI22xp33_ASAP7_75t_R g110688 (.A1(n_52),
    .A2(n_346),
    .B1(n_157),
    .B2(n_8327),
    .Y(n_429));
 AOI22xp5_ASAP7_75t_R g110689 (.A1(n_336),
    .A2(n_138),
    .B1(n_337),
    .B2(n_8278),
    .Y(n_428));
 OAI22xp5_ASAP7_75t_L g110690 (.A1(n_294),
    .A2(n_8246),
    .B1(n_204),
    .B2(w1[29]),
    .Y(n_691));
 OAI22xp33_ASAP7_75t_R g110691 (.A1(u0_n_32675),
    .A2(n_8315),
    .B1(w1[26]),
    .B2(n_232),
    .Y(n_689));
 OAI22xp5_ASAP7_75t_SL g110692 (.A1(n_367),
    .A2(n_8325),
    .B1(w0[17]),
    .B2(n_203),
    .Y(n_427));
 OAI22xp33_ASAP7_75t_SL g110693 (.A1(n_310),
    .A2(n_8244),
    .B1(w0[29]),
    .B2(n_238),
    .Y(n_687));
 OAI22xp33_ASAP7_75t_L g110694 (.A1(u0_n_32683),
    .A2(n_8334),
    .B1(w3[10]),
    .B2(n_362),
    .Y(n_426));
 AOI22xp5_ASAP7_75t_R g110695 (.A1(w3[29]),
    .A2(n_221),
    .B1(u0_n_32689),
    .B2(n_8250),
    .Y(n_425));
 AOI22xp5_ASAP7_75t_L g110696 (.A1(n_357),
    .A2(n_210),
    .B1(n_356),
    .B2(n_8227),
    .Y(n_424));
 AOI22xp5_ASAP7_75t_L g110697 (.A1(w3[24]),
    .A2(n_360),
    .B1(u0_n_32743),
    .B2(n_8294),
    .Y(n_423));
 OAI22xp5_ASAP7_75t_L g110698 (.A1(n_295),
    .A2(n_8248),
    .B1(w2[29]),
    .B2(n_236),
    .Y(n_685));
 OAI22xp5_ASAP7_75t_L g110699 (.A1(n_370),
    .A2(n_8325),
    .B1(w0[10]),
    .B2(n_203),
    .Y(n_422));
 AOI22xp33_ASAP7_75t_R g110700 (.A1(n_235),
    .A2(n_213),
    .B1(n_8300),
    .B2(n_211),
    .Y(n_421));
 OAI22xp5_ASAP7_75t_SL g110701 (.A1(n_44),
    .A2(n_145),
    .B1(n_43),
    .B2(n_144),
    .Y(n_420));
 OAI22xp5_ASAP7_75t_L g110702 (.A1(n_8270),
    .A2(n_138),
    .B1(n_158),
    .B2(n_8278),
    .Y(n_419));
 AOI22xp5_ASAP7_75t_SL g110703 (.A1(n_130),
    .A2(n_8272),
    .B1(n_199),
    .B2(n_131),
    .Y(n_418));
 AOI22xp33_ASAP7_75t_L g110704 (.A1(n_8274),
    .A2(n_138),
    .B1(n_153),
    .B2(n_8278),
    .Y(n_417));
 OAI22xp5_ASAP7_75t_L g110705 (.A1(n_8282),
    .A2(n_138),
    .B1(n_8278),
    .B2(n_163),
    .Y(n_416));
 OAI22xp5_ASAP7_75t_L g110706 (.A1(n_8262),
    .A2(n_8723),
    .B1(n_8280),
    .B2(n_143),
    .Y(n_683));
 OAI22xp5_ASAP7_75t_SL g110707 (.A1(n_342),
    .A2(n_145),
    .B1(n_344),
    .B2(n_144),
    .Y(n_415));
 OAI22xp33_ASAP7_75t_R g110708 (.A1(n_126),
    .A2(n_8274),
    .B1(n_8241),
    .B2(n_153),
    .Y(n_414));
 OAI22xp33_ASAP7_75t_R g110709 (.A1(n_172),
    .A2(n_8766),
    .B1(n_8268),
    .B2(n_8760),
    .Y(n_413));
 AOI22xp5_ASAP7_75t_L g110710 (.A1(n_63),
    .A2(n_8275),
    .B1(n_334),
    .B2(n_161),
    .Y(n_412));
 AOI22xp33_ASAP7_75t_R g110711 (.A1(n_8249),
    .A2(n_158),
    .B1(n_338),
    .B2(n_8270),
    .Y(n_411));
 OAI22xp5_ASAP7_75t_R g110712 (.A1(n_135),
    .A2(n_8262),
    .B1(n_8254),
    .B2(n_143),
    .Y(n_410));
 OAI22xp33_ASAP7_75t_R g110713 (.A1(n_8248),
    .A2(n_151),
    .B1(n_236),
    .B2(n_8269),
    .Y(n_409));
 AOI22xp5_ASAP7_75t_SL g110714 (.A1(n_204),
    .A2(n_8268),
    .B1(n_8246),
    .B2(n_172),
    .Y(n_408));
 AOI22xp33_ASAP7_75t_R g110715 (.A1(n_8290),
    .A2(n_360),
    .B1(n_8294),
    .B2(n_156),
    .Y(n_407));
 OAI22xp33_ASAP7_75t_R g110716 (.A1(n_55),
    .A2(n_224),
    .B1(n_54),
    .B2(n_60),
    .Y(n_406));
 AOI22xp5_ASAP7_75t_SL g110717 (.A1(n_209),
    .A2(n_8268),
    .B1(n_8238),
    .B2(n_172),
    .Y(n_405));
 OAI22xp33_ASAP7_75t_R g110718 (.A1(n_8296),
    .A2(n_206),
    .B1(n_177),
    .B2(n_207),
    .Y(n_404));
 OAI22xp5_ASAP7_75t_R g110719 (.A1(n_8267),
    .A2(n_161),
    .B1(n_228),
    .B2(n_8275),
    .Y(n_681));
 OAI22xp5_ASAP7_75t_R g110720 (.A1(n_207),
    .A2(n_167),
    .B1(n_37),
    .B2(n_206),
    .Y(n_403));
 OAI22xp5_ASAP7_75t_R g110721 (.A1(n_8236),
    .A2(n_228),
    .B1(n_173),
    .B2(n_8267),
    .Y(n_679));
 AOI22xp5_ASAP7_75t_L g110722 (.A1(n_8291),
    .A2(n_174),
    .B1(n_225),
    .B2(n_8287),
    .Y(n_677));
 AOI22xp33_ASAP7_75t_L g110723 (.A1(n_361),
    .A2(n_8260),
    .B1(n_148),
    .B2(n_8252),
    .Y(n_402));
 OAI22xp33_ASAP7_75t_R g110724 (.A1(n_152),
    .A2(n_8226),
    .B1(n_8222),
    .B2(n_208),
    .Y(n_401));
 OAI22xp5_ASAP7_75t_SL g110725 (.A1(n_190),
    .A2(n_8258),
    .B1(n_8266),
    .B2(n_242),
    .Y(n_400));
 OAI22xp33_ASAP7_75t_R g110726 (.A1(n_8286),
    .A2(n_156),
    .B1(n_8290),
    .B2(n_222),
    .Y(n_399));
 AOI22xp5_ASAP7_75t_L g110727 (.A1(n_8221),
    .A2(n_218),
    .B1(n_8225),
    .B2(n_8738),
    .Y(n_398));
 OAI22xp5_ASAP7_75t_L g110728 (.A1(n_8303),
    .A2(n_346),
    .B1(n_237),
    .B2(n_8327),
    .Y(n_397));
 AOI22xp33_ASAP7_75t_SL g110729 (.A1(n_54),
    .A2(n_229),
    .B1(n_55),
    .B2(n_8285),
    .Y(n_675));
 AOI22xp5_ASAP7_75t_SL g110730 (.A1(n_8224),
    .A2(n_168),
    .B1(n_8220),
    .B2(n_234),
    .Y(n_673));
 AOI22xp5_ASAP7_75t_SL g110731 (.A1(n_61),
    .A2(n_37),
    .B1(n_231),
    .B2(n_167),
    .Y(n_671));
 OAI22xp33_ASAP7_75t_R g110732 (.A1(n_8291),
    .A2(n_175),
    .B1(n_225),
    .B2(n_8295),
    .Y(n_396));
 AOI22xp5_ASAP7_75t_L g110733 (.A1(n_8219),
    .A2(n_356),
    .B1(n_357),
    .B2(n_58),
    .Y(n_395));
 OAI22xp33_ASAP7_75t_L g110734 (.A1(n_8240),
    .A2(n_151),
    .B1(n_241),
    .B2(n_8269),
    .Y(n_394));
 OAI22xp5_ASAP7_75t_L g110735 (.A1(n_215),
    .A2(n_174),
    .B1(n_214),
    .B2(n_8287),
    .Y(n_669));
 AOI22xp33_ASAP7_75t_L g110736 (.A1(n_8247),
    .A2(n_151),
    .B1(n_330),
    .B2(n_8269),
    .Y(n_393));
 AOI22xp5_ASAP7_75t_SL g110737 (.A1(n_116),
    .A2(n_8282),
    .B1(n_114),
    .B2(n_163),
    .Y(n_392));
 OAI22xp33_ASAP7_75t_R g110738 (.A1(n_194),
    .A2(n_8259),
    .B1(n_8279),
    .B2(n_119),
    .Y(n_391));
 AOI22xp5_ASAP7_75t_L g110739 (.A1(n_8300),
    .A2(n_8872),
    .B1(n_235),
    .B2(n_8881),
    .Y(n_390));
 OAI22xp5_ASAP7_75t_R g110740 (.A1(n_50),
    .A2(n_223),
    .B1(n_8331),
    .B2(n_137),
    .Y(n_389));
 OAI22xp5_ASAP7_75t_R g110741 (.A1(n_8313),
    .A2(n_8872),
    .B1(n_8301),
    .B2(n_240),
    .Y(n_388));
 AOI22xp33_ASAP7_75t_R g110742 (.A1(n_222),
    .A2(n_8249),
    .B1(n_8286),
    .B2(n_338),
    .Y(n_387));
 OAI22xp33_ASAP7_75t_R g110743 (.A1(n_215),
    .A2(n_122),
    .B1(n_214),
    .B2(n_8243),
    .Y(n_386));
 OAI22xp33_ASAP7_75t_L g110744 (.A1(n_231),
    .A2(n_8688),
    .B1(n_61),
    .B2(n_8245),
    .Y(n_385));
 AOI22xp5_ASAP7_75t_L g110745 (.A1(n_63),
    .A2(n_8267),
    .B1(n_334),
    .B2(n_228),
    .Y(n_667));
 OAI22xp5_ASAP7_75t_SL g110746 (.A1(n_62),
    .A2(n_211),
    .B1(n_324),
    .B2(n_213),
    .Y(n_666));
 OAI22xp5_ASAP7_75t_R g110747 (.A1(n_8230),
    .A2(n_208),
    .B1(n_8226),
    .B2(n_227),
    .Y(n_665));
 OAI22xp5_ASAP7_75t_SL g110748 (.A1(n_344),
    .A2(n_353),
    .B1(n_342),
    .B2(n_351),
    .Y(n_664));
 OAI22xp5_ASAP7_75t_L g110749 (.A1(n_239),
    .A2(n_8329),
    .B1(n_8317),
    .B2(n_347),
    .Y(n_663));
 AOI22x1_ASAP7_75t_SL g110750 (.A1(n_8688),
    .A2(n_8224),
    .B1(n_234),
    .B2(n_8245),
    .Y(n_661));
 AO22x2_ASAP7_75t_SL g110751 (.A1(n_7537),
    .A2(n_210),
    .B1(n_8227),
    .B2(n_332),
    .Y(n_660));
 OAI22xp5_ASAP7_75t_SL g110752 (.A1(n_8305),
    .A2(n_239),
    .B1(n_8317),
    .B2(n_191),
    .Y(n_656));
 AOI22xp5_ASAP7_75t_SL g110753 (.A1(n_8252),
    .A2(n_238),
    .B1(n_361),
    .B2(n_8244),
    .Y(n_655));
 AOI22xp5_ASAP7_75t_SL g110754 (.A1(n_175),
    .A2(n_8259),
    .B1(n_8295),
    .B2(n_119),
    .Y(n_653));
 AOI22xp5_ASAP7_75t_SL g110755 (.A1(n_186),
    .A2(n_8259),
    .B1(n_8231),
    .B2(n_119),
    .Y(n_651));
 AO22x1_ASAP7_75t_SL g110756 (.A1(n_8273),
    .A2(n_151),
    .B1(n_8269),
    .B2(n_351),
    .Y(n_648));
 OA22x2_ASAP7_75t_SL g110757 (.A1(n_8287),
    .A2(n_122),
    .B1(n_174),
    .B2(n_8243),
    .Y(n_647));
 OAI22xp5_ASAP7_75t_R g110758 (.A1(n_8224),
    .A2(n_202),
    .B1(n_234),
    .B2(n_8228),
    .Y(n_82));
 OAI22xp5_ASAP7_75t_SL g110759 (.A1(n_8290),
    .A2(n_338),
    .B1(n_156),
    .B2(n_8249),
    .Y(n_644));
 AO22x1_ASAP7_75t_SL g110760 (.A1(n_8249),
    .A2(n_208),
    .B1(n_8226),
    .B2(n_338),
    .Y(n_643));
 AOI22xp5_ASAP7_75t_SL g110761 (.A1(n_8258),
    .A2(n_221),
    .B1(n_8250),
    .B2(n_242),
    .Y(n_640));
 OAI22x1_ASAP7_75t_SL g110762 (.A1(n_177),
    .A2(n_8261),
    .B1(n_8296),
    .B2(n_8933),
    .Y(n_638));
 XOR2xp5_ASAP7_75t_SL g110763 (.A(n_8261),
    .B(n_8232),
    .Y(n_637));
 AOI22xp5_ASAP7_75t_SL g110764 (.A1(n_37),
    .A2(n_8679),
    .B1(n_167),
    .B2(n_8687),
    .Y(n_635));
 AOI22xp5_ASAP7_75t_SL g110766 (.A1(n_8256),
    .A2(n_164),
    .B1(n_8264),
    .B2(n_59),
    .Y(n_632));
 XOR2xp5_ASAP7_75t_SL g110767 (.A(n_8239),
    .B(n_8221),
    .Y(n_631));
 OAI22xp5_ASAP7_75t_L g110768 (.A1(n_350),
    .A2(n_8332),
    .B1(n_8320),
    .B2(n_184),
    .Y(n_629));
 OAI22xp5_ASAP7_75t_L g110769 (.A1(n_8320),
    .A2(n_196),
    .B1(n_8308),
    .B2(n_350),
    .Y(n_628));
 AOI22xp5_ASAP7_75t_SL g110770 (.A1(n_152),
    .A2(n_8241),
    .B1(n_126),
    .B2(n_8222),
    .Y(n_626));
 AOI22x1_ASAP7_75t_SL g110771 (.A1(n_179),
    .A2(n_44),
    .B1(n_178),
    .B2(n_42),
    .Y(n_625));
 OAI22xp5_ASAP7_75t_SL g110772 (.A1(n_58),
    .A2(n_8235),
    .B1(n_147),
    .B2(n_8219),
    .Y(n_620));
 OAI22x1_ASAP7_75t_SL g110774 (.A1(n_172),
    .A2(n_8272),
    .B1(n_199),
    .B2(n_8268),
    .Y(n_618));
 OA22x2_ASAP7_75t_L g110775 (.A1(n_8242),
    .A2(n_221),
    .B1(n_8250),
    .B2(n_349),
    .Y(n_617));
 AOI22xp5_ASAP7_75t_SL g110776 (.A1(n_8220),
    .A2(n_130),
    .B1(n_168),
    .B2(n_131),
    .Y(n_80));
 AOI22xp5_ASAP7_75t_L g110777 (.A1(n_8276),
    .A2(n_8723),
    .B1(n_8280),
    .B2(n_165),
    .Y(n_615));
 AOI22xp5_ASAP7_75t_SL g110778 (.A1(n_8887),
    .A2(n_113),
    .B1(n_8884),
    .B2(n_117),
    .Y(n_614));
 OAI22xp5_ASAP7_75t_SL g110779 (.A1(n_8265),
    .A2(n_335),
    .B1(n_113),
    .B2(n_7447),
    .Y(n_78));
 AOI22xp5_ASAP7_75t_SL g110780 (.A1(n_63),
    .A2(n_8259),
    .B1(n_334),
    .B2(n_119),
    .Y(n_611));
 OAI22xp5_ASAP7_75t_L g110781 (.A1(n_8261),
    .A2(n_8760),
    .B1(n_8933),
    .B2(n_8253),
    .Y(n_610));
 AO22x1_ASAP7_75t_SL g110782 (.A1(n_127),
    .A2(n_121),
    .B1(n_8255),
    .B2(n_43),
    .Y(n_608));
 AOI22xp5_ASAP7_75t_SL g110783 (.A1(n_8255),
    .A2(n_8785),
    .B1(n_127),
    .B2(n_8779),
    .Y(n_606));
 OAI22xp5_ASAP7_75t_SL g110784 (.A1(n_8323),
    .A2(n_355),
    .B1(n_150),
    .B2(n_8311),
    .Y(n_605));
 OAI22xp5_ASAP7_75t_SL g110785 (.A1(n_330),
    .A2(n_8239),
    .B1(n_8247),
    .B2(n_8780),
    .Y(n_76));
 OAI22xp5_ASAP7_75t_SL g110786 (.A1(n_219),
    .A2(n_226),
    .B1(n_220),
    .B2(n_8229),
    .Y(n_603));
 OAI22xp5_ASAP7_75t_SL g110787 (.A1(n_8230),
    .A2(n_335),
    .B1(n_227),
    .B2(n_7447),
    .Y(n_601));
 OAI22xp5_ASAP7_75t_L g110788 (.A1(n_8229),
    .A2(n_127),
    .B1(n_8255),
    .B2(n_226),
    .Y(n_75));
 AOI22xp5_ASAP7_75t_SL g110790 (.A1(n_8236),
    .A2(n_238),
    .B1(n_173),
    .B2(n_8244),
    .Y(n_598));
 OAI22xp5_ASAP7_75t_SL g110791 (.A1(n_232),
    .A2(n_8303),
    .B1(n_8315),
    .B2(n_237),
    .Y(n_596));
 XOR2x2_ASAP7_75t_SL g110792 (.A(n_8247),
    .B(n_55),
    .Y(n_594));
 AO22x1_ASAP7_75t_SL g110793 (.A1(n_8325),
    .A2(n_240),
    .B1(n_8313),
    .B2(n_203),
    .Y(n_591));
 AOI22xp5_ASAP7_75t_L g110794 (.A1(n_356),
    .A2(n_8243),
    .B1(n_357),
    .B2(n_122),
    .Y(n_590));
 AOI22xp5_ASAP7_75t_SL g110795 (.A1(n_8291),
    .A2(n_332),
    .B1(n_225),
    .B2(n_7537),
    .Y(n_587));
 AOI22xp5_ASAP7_75t_SL g110796 (.A1(n_8245),
    .A2(n_130),
    .B1(n_131),
    .B2(n_8678),
    .Y(n_585));
 AOI22xp5_ASAP7_75t_SL g110797 (.A1(n_147),
    .A2(n_8243),
    .B1(n_8235),
    .B2(n_122),
    .Y(n_584));
 OAI22xp5_ASAP7_75t_SL g110798 (.A1(n_363),
    .A2(n_8331),
    .B1(n_8319),
    .B2(n_223),
    .Y(n_74));
 AOI22x1_ASAP7_75t_SL g110799 (.A1(n_204),
    .A2(n_8238),
    .B1(n_8246),
    .B2(n_209),
    .Y(n_581));
 AOI22xp5_ASAP7_75t_L g110800 (.A1(n_283),
    .A2(n_8328),
    .B1(n_285),
    .B2(n_217),
    .Y(n_579));
 XNOR2x2_ASAP7_75t_SL g110803 (.A(n_8248),
    .B(n_8240),
    .Y(n_72));
 AO22x1_ASAP7_75t_SL g110804 (.A1(n_229),
    .A2(n_8783),
    .B1(n_8285),
    .B2(n_8780),
    .Y(n_576));
 XOR2x2_ASAP7_75t_SL g110805 (.A(n_131),
    .B(n_61),
    .Y(n_574));
 OAI22xp5_ASAP7_75t_SL g110806 (.A1(n_60),
    .A2(n_8255),
    .B1(n_8293),
    .B2(n_127),
    .Y(n_572));
 AO22x1_ASAP7_75t_SL g110807 (.A1(n_222),
    .A2(n_8241),
    .B1(n_8286),
    .B2(n_126),
    .Y(n_571));
 AOI22x1_ASAP7_75t_SL g110808 (.A1(n_214),
    .A2(n_8235),
    .B1(n_147),
    .B2(n_8283),
    .Y(n_71));
 AO22x2_ASAP7_75t_SL g110810 (.A1(n_8249),
    .A2(n_126),
    .B1(n_8241),
    .B2(n_338),
    .Y(n_565));
 INVxp33_ASAP7_75t_R g110811 (.A(n_383),
    .Y(n_384));
 NAND2xp33_ASAP7_75t_R g110813 (.A(w0[7]),
    .B(n_8279),
    .Y(n_381));
 NOR2xp33_ASAP7_75t_R g110814 (.A(dcnt[1]),
    .B(dcnt[0]),
    .Y(n_383));
 INVxp33_ASAP7_75t_R g110815 (.A(n_379),
    .Y(n_380));
 NAND2xp33_ASAP7_75t_R g110816 (.A(w3[30]),
    .B(n_8274),
    .Y(n_378));
 NAND2xp33_ASAP7_75t_R g110817 (.A(w0[22]),
    .B(n_8279),
    .Y(n_377));
 NAND2xp5_ASAP7_75t_SL g110818 (.A(n_7447),
    .B(n_360),
    .Y(n_376));
 NAND2xp33_ASAP7_75t_R g110819 (.A(ld),
    .B(rst),
    .Y(n_379));
 INVxp67_ASAP7_75t_R g110820 (.A(n_8218),
    .Y(n_375));
 INVxp33_ASAP7_75t_R g110827 (.A(w0[12]),
    .Y(n_373));
 INVxp67_ASAP7_75t_R g110829 (.A(n_8314),
    .Y(n_371));
 INVxp33_ASAP7_75t_R g110833 (.A(w0[10]),
    .Y(n_370));
 INVxp33_ASAP7_75t_R g110834 (.A(w2[7]),
    .Y(n_369));
 INVxp33_ASAP7_75t_R g110835 (.A(w2[0]),
    .Y(n_368));
 INVxp33_ASAP7_75t_R g110836 (.A(w0[17]),
    .Y(n_367));
 INVxp33_ASAP7_75t_R g110838 (.A(w0[13]),
    .Y(n_365));
 INVx1_ASAP7_75t_SL g110842 (.A(n_8319),
    .Y(n_363));
 INVxp67_ASAP7_75t_SL g110844 (.A(n_8334),
    .Y(n_362));
 INVx2_ASAP7_75t_SL g110846 (.A(n_8252),
    .Y(n_361));
 INVx1_ASAP7_75t_SL g110847 (.A(n_8294),
    .Y(n_360));
 INVx2_ASAP7_75t_SL g110851 (.A(n_357),
    .Y(n_356));
 INVx1_ASAP7_75t_R g110852 (.A(n_8311),
    .Y(n_355));
 INVxp33_ASAP7_75t_R g110854 (.A(n_351),
    .Y(n_353));
 INVx1_ASAP7_75t_L g110858 (.A(n_8320),
    .Y(n_350));
 INVxp67_ASAP7_75t_L g110863 (.A(n_69),
    .Y(n_70));
 INVx1_ASAP7_75t_SL g110865 (.A(n_8242),
    .Y(n_349));
 INVx1_ASAP7_75t_SL g110866 (.A(n_8304),
    .Y(n_348));
 INVxp67_ASAP7_75t_R g110870 (.A(n_68),
    .Y(n_67));
 INVx2_ASAP7_75t_L g110871 (.A(n_8333),
    .Y(n_68));
 INVxp67_ASAP7_75t_SL g110872 (.A(n_8329),
    .Y(n_347));
 INVx1_ASAP7_75t_SL g110873 (.A(n_8327),
    .Y(n_346));
 INVx2_ASAP7_75t_SL g110874 (.A(n_8302),
    .Y(n_345));
 INVx1_ASAP7_75t_L g110875 (.A(n_342),
    .Y(n_344));
 BUFx2_ASAP7_75t_L g110876 (.A(n_8277),
    .Y(n_342));
 INVx1_ASAP7_75t_SL g110879 (.A(n_8337),
    .Y(n_340));
 INVx3_ASAP7_75t_SL g110888 (.A(n_8249),
    .Y(n_338));
 INVx1_ASAP7_75t_L g110889 (.A(n_337),
    .Y(n_336));
 INVxp67_ASAP7_75t_R g110890 (.A(n_7447),
    .Y(n_337));
 INVx1_ASAP7_75t_L g110891 (.A(n_7447),
    .Y(n_335));
 HB1xp67_ASAP7_75t_L g110892 (.A(n_7537),
    .Y(n_334));
 INVx1_ASAP7_75t_L g110896 (.A(n_331),
    .Y(n_63));
 HB1xp67_ASAP7_75t_SL g110897 (.A(n_7537),
    .Y(n_331));
 INVx2_ASAP7_75t_SL g110898 (.A(n_8247),
    .Y(n_330));
 INVxp33_ASAP7_75t_R g110900 (.A(w1[15]),
    .Y(n_328));
 INVxp33_ASAP7_75t_R g110902 (.A(w2[2]),
    .Y(n_326));
 INVx1_ASAP7_75t_R g110903 (.A(n_8324),
    .Y(n_325));
 INVxp33_ASAP7_75t_R g110908 (.A(w2[23]),
    .Y(n_322));
 INVxp33_ASAP7_75t_R g110909 (.A(n_11482),
    .Y(n_321));
 INVxp33_ASAP7_75t_R g110911 (.A(w0[0]),
    .Y(n_320));
 INVxp33_ASAP7_75t_R g110912 (.A(w1[3]),
    .Y(n_319));
 INVxp33_ASAP7_75t_R g110916 (.A(w1[22]),
    .Y(n_316));
 INVxp33_ASAP7_75t_R g110918 (.A(n_11346),
    .Y(n_314));
 INVxp33_ASAP7_75t_R g110919 (.A(w0[11]),
    .Y(n_313));
 INVxp33_ASAP7_75t_R g110920 (.A(w0[15]),
    .Y(n_312));
 INVxp33_ASAP7_75t_R g110921 (.A(w0[3]),
    .Y(n_311));
 INVxp33_ASAP7_75t_R g110922 (.A(w0[29]),
    .Y(n_310));
 INVxp33_ASAP7_75t_R g110923 (.A(w0[25]),
    .Y(n_309));
 INVxp33_ASAP7_75t_R g110925 (.A(w1[30]),
    .Y(u0_n_32676));
 INVxp33_ASAP7_75t_R g110926 (.A(w0[30]),
    .Y(n_306));
 INVxp33_ASAP7_75t_R g110927 (.A(w2[5]),
    .Y(n_305));
 INVxp33_ASAP7_75t_R g110929 (.A(w1[12]),
    .Y(n_304));
 INVxp33_ASAP7_75t_R g110930 (.A(w2[10]),
    .Y(n_303));
 INVxp33_ASAP7_75t_R g110931 (.A(w2[21]),
    .Y(n_302));
 INVxp33_ASAP7_75t_R g110932 (.A(w0[1]),
    .Y(n_301));
 INVxp33_ASAP7_75t_R g110934 (.A(w2[27]),
    .Y(n_300));
 INVxp33_ASAP7_75t_R g110935 (.A(w2[4]),
    .Y(n_299));
 INVxp33_ASAP7_75t_R g110936 (.A(w1[5]),
    .Y(n_298));
 INVxp33_ASAP7_75t_R g110938 (.A(w0[27]),
    .Y(n_296));
 INVxp33_ASAP7_75t_R g110939 (.A(w2[29]),
    .Y(n_295));
 INVxp33_ASAP7_75t_R g110940 (.A(w1[29]),
    .Y(n_294));
 INVxp33_ASAP7_75t_R g110942 (.A(w1[28]),
    .Y(n_293));
 INVxp67_ASAP7_75t_L g110943 (.A(n_8322),
    .Y(n_292));
 INVxp33_ASAP7_75t_R g110945 (.A(w1[24]),
    .Y(n_291));
 INVxp33_ASAP7_75t_R g110946 (.A(w3[16]),
    .Y(n_290));
 INVxp33_ASAP7_75t_R g110947 (.A(w2[18]),
    .Y(n_289));
 INVxp67_ASAP7_75t_R g110951 (.A(n_283),
    .Y(n_285));
 INVx2_ASAP7_75t_SL g110952 (.A(n_8316),
    .Y(n_283));
 INVxp33_ASAP7_75t_R g110954 (.A(w1[1]),
    .Y(n_282));
 INVxp33_ASAP7_75t_R g110955 (.A(w3[25]),
    .Y(n_281));
 INVxp33_ASAP7_75t_R g110957 (.A(w2[31]),
    .Y(n_280));
 INVxp33_ASAP7_75t_R g110958 (.A(w0[2]),
    .Y(n_279));
 INVxp33_ASAP7_75t_R g110959 (.A(w0[23]),
    .Y(n_278));
 INVxp33_ASAP7_75t_R g110966 (.A(w1[23]),
    .Y(n_272));
 INVxp33_ASAP7_75t_R g110967 (.A(w1[6]),
    .Y(n_271));
 INVxp33_ASAP7_75t_R g110968 (.A(w1[31]),
    .Y(n_270));
 INVxp33_ASAP7_75t_R g110969 (.A(w1[20]),
    .Y(n_269));
 INVxp33_ASAP7_75t_R g110970 (.A(w0[5]),
    .Y(n_268));
 INVxp33_ASAP7_75t_R g110971 (.A(w2[14]),
    .Y(n_267));
 INVxp33_ASAP7_75t_R g110972 (.A(w1[4]),
    .Y(n_266));
 INVxp33_ASAP7_75t_R g110973 (.A(w2[16]),
    .Y(n_265));
 INVxp67_ASAP7_75t_R g110974 (.A(w2[26]),
    .Y(n_264));
 INVxp33_ASAP7_75t_R g110975 (.A(w1[13]),
    .Y(n_263));
 INVxp33_ASAP7_75t_R g110977 (.A(w0[31]),
    .Y(n_261));
 INVxp33_ASAP7_75t_R g110978 (.A(w0[20]),
    .Y(n_260));
 INVxp33_ASAP7_75t_R g110979 (.A(w2[6]),
    .Y(n_259));
 INVxp33_ASAP7_75t_R g110980 (.A(w2[25]),
    .Y(n_258));
 INVxp33_ASAP7_75t_R g110983 (.A(w0[24]),
    .Y(n_256));
 INVxp33_ASAP7_75t_R g110986 (.A(w2[13]),
    .Y(n_255));
 INVxp33_ASAP7_75t_R g110987 (.A(w2[15]),
    .Y(n_254));
 INVxp67_ASAP7_75t_R g110988 (.A(w0[26]),
    .Y(n_253));
 INVxp33_ASAP7_75t_R g110989 (.A(w1[21]),
    .Y(n_252));
 INVxp33_ASAP7_75t_R g110994 (.A(w0[19]),
    .Y(n_247));
 INVxp33_ASAP7_75t_R g110996 (.A(w0[4]),
    .Y(n_245));
 INVxp33_ASAP7_75t_R g110998 (.A(w1[2]),
    .Y(n_243));
 INVx2_ASAP7_75t_SL g110999 (.A(n_8258),
    .Y(n_242));
 INVxp33_ASAP7_75t_R g111000 (.A(n_8240),
    .Y(n_241));
 INVx1_ASAP7_75t_SL g111001 (.A(n_8313),
    .Y(n_240));
 INVx2_ASAP7_75t_L g111002 (.A(n_8317),
    .Y(n_239));
 INVx2_ASAP7_75t_L g111003 (.A(n_8244),
    .Y(n_238));
 INVx1_ASAP7_75t_SL g111004 (.A(n_8303),
    .Y(n_237));
 INVxp33_ASAP7_75t_R g111005 (.A(n_8248),
    .Y(n_236));
 INVx2_ASAP7_75t_SL g111006 (.A(n_8300),
    .Y(n_235));
 INVx3_ASAP7_75t_SL g111007 (.A(n_8224),
    .Y(n_234));
 INVxp67_ASAP7_75t_SL g111008 (.A(n_8336),
    .Y(n_233));
 INVx2_ASAP7_75t_SL g111009 (.A(n_8315),
    .Y(n_232));
 INVxp67_ASAP7_75t_R g111011 (.A(n_61),
    .Y(n_231));
 INVx1_ASAP7_75t_SL g111012 (.A(n_8284),
    .Y(n_61));
 INVxp67_ASAP7_75t_R g111015 (.A(n_8326),
    .Y(n_230));
 INVx2_ASAP7_75t_SL g111016 (.A(n_8285),
    .Y(n_229));
 INVx3_ASAP7_75t_SL g111017 (.A(n_8267),
    .Y(n_228));
 INVx1_ASAP7_75t_L g111018 (.A(n_8230),
    .Y(n_227));
 INVx1_ASAP7_75t_SL g111019 (.A(n_8229),
    .Y(n_226));
 INVx1_ASAP7_75t_L g111020 (.A(n_8291),
    .Y(n_225));
 INVxp67_ASAP7_75t_R g111022 (.A(n_60),
    .Y(n_224));
 INVx1_ASAP7_75t_SL g111023 (.A(n_8293),
    .Y(n_60));
 INVx1_ASAP7_75t_SL g111024 (.A(n_8331),
    .Y(n_223));
 INVx1_ASAP7_75t_SL g111025 (.A(n_8286),
    .Y(n_222));
 INVx1_ASAP7_75t_L g111026 (.A(n_8250),
    .Y(n_221));
 INVx1_ASAP7_75t_L g111027 (.A(n_219),
    .Y(n_220));
 INVx1_ASAP7_75t_L g111028 (.A(n_218),
    .Y(n_219));
 INVx2_ASAP7_75t_SL g111029 (.A(n_8225),
    .Y(n_218));
 INVx1_ASAP7_75t_L g111030 (.A(n_8328),
    .Y(n_217));
 INVx2_ASAP7_75t_SL g111031 (.A(n_8283),
    .Y(n_214));
 INVxp67_ASAP7_75t_R g111032 (.A(n_214),
    .Y(n_215));
 HB1xp67_ASAP7_75t_R g111034 (.A(n_8312),
    .Y(n_213));
 INVx1_ASAP7_75t_SL g111036 (.A(n_8312),
    .Y(n_211));
 INVx1_ASAP7_75t_SL g111037 (.A(n_8227),
    .Y(n_210));
 INVx1_ASAP7_75t_L g111038 (.A(n_8238),
    .Y(n_209));
 INVx1_ASAP7_75t_L g111039 (.A(n_8226),
    .Y(n_208));
 INVxp67_ASAP7_75t_R g111041 (.A(n_207),
    .Y(n_206));
 INVx2_ASAP7_75t_L g111043 (.A(n_8246),
    .Y(n_204));
 INVx2_ASAP7_75t_SL g111044 (.A(n_8325),
    .Y(n_203));
 INVx1_ASAP7_75t_SL g111045 (.A(n_8228),
    .Y(n_202));
 INVxp67_ASAP7_75t_R g111048 (.A(n_59),
    .Y(n_200));
 INVx1_ASAP7_75t_SL g111049 (.A(n_8256),
    .Y(n_59));
 INVx3_ASAP7_75t_SL g111050 (.A(n_8272),
    .Y(n_199));
 INVxp67_ASAP7_75t_R g111054 (.A(n_58),
    .Y(n_57));
 INVx1_ASAP7_75t_SL g111055 (.A(n_8219),
    .Y(n_58));
 INVx1_ASAP7_75t_SL g111061 (.A(n_8308),
    .Y(n_196));
 INVx1_ASAP7_75t_SL g111062 (.A(n_8342),
    .Y(n_195));
 INVx2_ASAP7_75t_SL g111063 (.A(n_8279),
    .Y(n_194));
 HB1xp67_ASAP7_75t_L g111064 (.A(n_8305),
    .Y(n_193));
 INVx2_ASAP7_75t_SL g111065 (.A(n_8305),
    .Y(n_191));
 INVx1_ASAP7_75t_SL g111067 (.A(n_8266),
    .Y(n_190));
 INVx1_ASAP7_75t_R g111068 (.A(n_8330),
    .Y(n_189));
 INVx1_ASAP7_75t_SL g111070 (.A(n_8318),
    .Y(n_187));
 INVx2_ASAP7_75t_SL g111071 (.A(n_8231),
    .Y(n_186));
 INVx1_ASAP7_75t_SL g111072 (.A(n_8332),
    .Y(n_184));
 INVxp67_ASAP7_75t_L g111074 (.A(n_182),
    .Y(n_183));
 INVx1_ASAP7_75t_L g111075 (.A(n_8309),
    .Y(n_182));
 INVx1_ASAP7_75t_L g111076 (.A(n_8309),
    .Y(n_181));
 INVxp67_ASAP7_75t_R g111077 (.A(n_8309),
    .Y(n_180));
 INVxp67_ASAP7_75t_R g111079 (.A(n_178),
    .Y(n_179));
 INVx3_ASAP7_75t_SL g111082 (.A(n_8296),
    .Y(n_177));
 HB1xp67_ASAP7_75t_L g111083 (.A(n_8232),
    .Y(n_176));
 INVx1_ASAP7_75t_SL g111085 (.A(n_8295),
    .Y(n_175));
 INVx2_ASAP7_75t_SL g111086 (.A(n_8287),
    .Y(n_174));
 INVx2_ASAP7_75t_SL g111087 (.A(n_8236),
    .Y(n_173));
 INVx1_ASAP7_75t_L g111091 (.A(n_55),
    .Y(n_54));
 INVx1_ASAP7_75t_SL g111092 (.A(n_8289),
    .Y(n_55));
 INVx2_ASAP7_75t_L g111093 (.A(n_8268),
    .Y(n_172));
 INVx2_ASAP7_75t_SL g111098 (.A(n_169),
    .Y(n_53));
 INVx2_ASAP7_75t_SL g111099 (.A(n_8220),
    .Y(n_168));
 INVx3_ASAP7_75t_SL g111100 (.A(n_37),
    .Y(n_167));
 INVx1_ASAP7_75t_SL g111101 (.A(n_8346),
    .Y(n_166));
 INVx1_ASAP7_75t_SL g111102 (.A(n_8276),
    .Y(n_165));
 INVx1_ASAP7_75t_SL g111103 (.A(n_8264),
    .Y(n_164));
 INVx1_ASAP7_75t_SL g111104 (.A(n_8282),
    .Y(n_163));
 INVx2_ASAP7_75t_SL g111105 (.A(n_8275),
    .Y(n_161));
 INVx2_ASAP7_75t_SL g111108 (.A(n_8310),
    .Y(n_159));
 INVx2_ASAP7_75t_SL g111109 (.A(n_8270),
    .Y(n_158));
 INVxp67_ASAP7_75t_R g111110 (.A(n_52),
    .Y(n_157));
 HB1xp67_ASAP7_75t_SL g111112 (.A(n_8339),
    .Y(n_52));
 INVx1_ASAP7_75t_SL g111113 (.A(n_8290),
    .Y(n_156));
 INVx1_ASAP7_75t_L g111115 (.A(n_8321),
    .Y(n_154));
 INVxp67_ASAP7_75t_SL g111116 (.A(n_8274),
    .Y(n_153));
 INVx2_ASAP7_75t_SL g111117 (.A(n_8222),
    .Y(n_152));
 INVx2_ASAP7_75t_SL g111118 (.A(n_8269),
    .Y(n_151));
 INVx2_ASAP7_75t_L g111119 (.A(n_8323),
    .Y(n_150));
 INVx1_ASAP7_75t_R g111122 (.A(n_149),
    .Y(n_51));
 INVx1_ASAP7_75t_L g111123 (.A(n_8298),
    .Y(n_149));
 INVxp67_ASAP7_75t_SL g111125 (.A(n_8260),
    .Y(n_148));
 INVx2_ASAP7_75t_SL g111126 (.A(n_8235),
    .Y(n_147));
 INVxp67_ASAP7_75t_L g111129 (.A(n_8281),
    .Y(n_145));
 HB1xp67_ASAP7_75t_L g111130 (.A(n_8281),
    .Y(n_144));
 INVx2_ASAP7_75t_SL g111131 (.A(n_8262),
    .Y(n_143));
 INVx1_ASAP7_75t_SL g111136 (.A(n_8278),
    .Y(n_138));
 INVxp67_ASAP7_75t_L g111138 (.A(n_50),
    .Y(n_137));
 HB1xp67_ASAP7_75t_R g111139 (.A(n_8343),
    .Y(n_50));
 INVx1_ASAP7_75t_SL g111140 (.A(n_8343),
    .Y(n_136));
 INVx2_ASAP7_75t_SL g111142 (.A(n_8338),
    .Y(n_134));
 INVx2_ASAP7_75t_SL g111143 (.A(n_131),
    .Y(n_130));
 INVxp67_ASAP7_75t_R g111150 (.A(n_49),
    .Y(n_128));
 INVxp67_ASAP7_75t_L g111151 (.A(n_129),
    .Y(n_49));
 INVx2_ASAP7_75t_L g111152 (.A(n_8255),
    .Y(n_127));
 INVx1_ASAP7_75t_R g111158 (.A(n_47),
    .Y(n_48));
 INVx2_ASAP7_75t_SL g111159 (.A(n_8345),
    .Y(n_47));
 INVx2_ASAP7_75t_L g111160 (.A(n_8241),
    .Y(n_126));
 INVx1_ASAP7_75t_L g111162 (.A(n_45),
    .Y(n_46));
 HB1xp67_ASAP7_75t_SL g111164 (.A(n_8340),
    .Y(n_45));
 INVx1_ASAP7_75t_SL g111167 (.A(n_8344),
    .Y(n_125));
 INVx2_ASAP7_75t_SL g111170 (.A(n_8243),
    .Y(n_122));
 INVx1_ASAP7_75t_L g111174 (.A(n_43),
    .Y(n_44));
 INVx1_ASAP7_75t_L g111175 (.A(n_8263),
    .Y(n_43));
 INVx1_ASAP7_75t_SL g111177 (.A(n_121),
    .Y(n_42));
 BUFx2_ASAP7_75t_SL g111178 (.A(n_8263),
    .Y(n_121));
 INVxp67_ASAP7_75t_R g111179 (.A(n_8263),
    .Y(n_120));
 INVx2_ASAP7_75t_SL g111181 (.A(n_8259),
    .Y(n_119));
 INVx1_ASAP7_75t_L g111183 (.A(n_117),
    .Y(n_116));
 BUFx2_ASAP7_75t_SL g111184 (.A(n_8265),
    .Y(n_117));
 INVxp67_ASAP7_75t_R g111185 (.A(n_113),
    .Y(n_114));
 INVx2_ASAP7_75t_SL g111186 (.A(n_8265),
    .Y(n_113));
 INVxp33_ASAP7_75t_R g111190 (.A(n_112),
    .Y(n_41));
 BUFx2_ASAP7_75t_R g111193 (.A(n_111),
    .Y(n_112));
 INVx1_ASAP7_75t_R g111200 (.A(n_111),
    .Y(n_40));
 HB1xp67_ASAP7_75t_R g111201 (.A(n_111),
    .Y(n_110));
 HB1xp67_ASAP7_75t_R g111202 (.A(n_111),
    .Y(n_109));
 HB1xp67_ASAP7_75t_R g111203 (.A(n_111),
    .Y(n_108));
 HB1xp67_ASAP7_75t_R g111204 (.A(n_111),
    .Y(n_107));
 HB1xp67_ASAP7_75t_R g111205 (.A(n_111),
    .Y(n_106));
 HB1xp67_ASAP7_75t_R g111206 (.A(n_111),
    .Y(n_105));
 HB1xp67_ASAP7_75t_R g111207 (.A(n_111),
    .Y(n_104));
 HB1xp67_ASAP7_75t_R g111208 (.A(n_111),
    .Y(n_103));
 HB1xp67_ASAP7_75t_R g111209 (.A(n_111),
    .Y(n_102));
 INVx2_ASAP7_75t_SL g111212 (.A(ld_r),
    .Y(n_111));
 INVxp33_ASAP7_75t_R g111215 (.A(n_101),
    .Y(n_39));
 INVxp33_ASAP7_75t_R g111219 (.A(n_101),
    .Y(n_100));
 INVxp33_ASAP7_75t_R g111220 (.A(n_101),
    .Y(n_99));
 INVxp33_ASAP7_75t_R g111222 (.A(n_101),
    .Y(n_98));
 INVxp33_ASAP7_75t_R g111224 (.A(n_95),
    .Y(n_97));
 INVxp33_ASAP7_75t_R g111225 (.A(n_95),
    .Y(n_96));
 HB1xp67_ASAP7_75t_R g111226 (.A(n_95),
    .Y(n_94));
 HB1xp67_ASAP7_75t_R g111227 (.A(n_95),
    .Y(n_93));
 HB1xp67_ASAP7_75t_R g111228 (.A(n_95),
    .Y(n_92));
 HB1xp67_ASAP7_75t_R g111229 (.A(n_95),
    .Y(n_91));
 INVxp67_ASAP7_75t_R g111230 (.A(n_101),
    .Y(n_95));
 INVxp67_ASAP7_75t_R g111231 (.A(ld),
    .Y(n_101));
 XNOR2xp5_ASAP7_75t_L g111261 (.A(n_961),
    .B(n_88),
    .Y(n_25));
 XNOR2xp5_ASAP7_75t_SL g111262 (.A(n_943),
    .B(n_606),
    .Y(n_24));
 XNOR2xp5_ASAP7_75t_L g111263 (.A(n_935),
    .B(n_912),
    .Y(n_23));
 XNOR2xp5_ASAP7_75t_SL g111264 (.A(n_12),
    .B(n_605),
    .Y(n_22));
 XOR2xp5_ASAP7_75t_L g111265 (.A(n_230),
    .B(n_922),
    .Y(n_21));
 XOR2xp5_ASAP7_75t_SL g111266 (.A(w2[3]),
    .B(n_89),
    .Y(n_20));
 XNOR2xp5_ASAP7_75t_SL g111267 (.A(n_1221),
    .B(n_911),
    .Y(n_19));
 XOR2xp5_ASAP7_75t_L g111268 (.A(w3[3]),
    .B(n_891),
    .Y(n_18));
 XOR2xp5_ASAP7_75t_SL g111269 (.A(n_1068),
    .B(n_635),
    .Y(n_17));
 XOR2xp5_ASAP7_75t_L g111270 (.A(n_1105),
    .B(n_628),
    .Y(n_16));
 XOR2xp5_ASAP7_75t_L g111271 (.A(n_416),
    .B(n_617),
    .Y(n_15));
 XNOR2xp5_ASAP7_75t_SL g111272 (.A(w0[9]),
    .B(n_587),
    .Y(n_14));
 XOR2x2_ASAP7_75t_SL g111273 (.A(n_8314),
    .B(n_8326),
    .Y(n_13));
 XOR2xp5_ASAP7_75t_R g111274 (.A(n_8335),
    .B(w0[28]),
    .Y(n_12));
 XOR2xp5_ASAP7_75t_L g111275 (.A(n_129),
    .B(w2[20]),
    .Y(n_11));
 XOR2xp5_ASAP7_75t_L g111276 (.A(n_8334),
    .B(n_8322),
    .Y(n_10));
 XNOR2xp5_ASAP7_75t_R g111277 (.A(w2[30]),
    .B(n_8273),
    .Y(n_9));
 XOR2xp5_ASAP7_75t_SL g111278 (.A(n_69),
    .B(n_8263),
    .Y(n_8));
 XNOR2xp5_ASAP7_75t_L g111279 (.A(w2[28]),
    .B(n_129),
    .Y(n_7));
 XOR2xp5_ASAP7_75t_L g111280 (.A(w2[11]),
    .B(n_178),
    .Y(n_6));
 XOR2xp5_ASAP7_75t_L g111281 (.A(w1[17]),
    .B(n_8340),
    .Y(n_5));
 XNOR2xp5_ASAP7_75t_R g111282 (.A(w2[19]),
    .B(n_178),
    .Y(n_4));
 XNOR2xp5_ASAP7_75t_R g111283 (.A(w1[27]),
    .B(n_8232),
    .Y(n_3));
 XNOR2xp5_ASAP7_75t_L g111284 (.A(w2[22]),
    .B(n_8281),
    .Y(n_2));
 XNOR2xp5_ASAP7_75t_L g111285 (.A(w1[25]),
    .B(n_8340),
    .Y(n_1));
 XNOR2xp5_ASAP7_75t_L g111286 (.A(n_8265),
    .B(n_8298),
    .Y(n_0));
 OR2x2_ASAP7_75t_SL g2 (.A(n_1846),
    .B(sa00[3]),
    .Y(n_1342));
 AO221x1_ASAP7_75t_SL g211727__2398 (.A1(n_8158),
    .A2(sa23[5]),
    .B1(n_8074),
    .B2(n_3493),
    .C(n_8165),
    .Y(n_8328));
 AO221x1_ASAP7_75t_SL g211731__5107 (.A1(n_8160),
    .A2(sa23[5]),
    .B1(n_8147),
    .B2(n_2704),
    .C(n_8152),
    .Y(n_8326));
 AO21x1_ASAP7_75t_SL g211732__6260 (.A1(sa23[5]),
    .A2(n_8164),
    .B(n_8167),
    .Y(n_8327));
 NAND3x1_ASAP7_75t_SL g211733__4319 (.A(n_8155),
    .B(n_8156),
    .C(n_8140),
    .Y(n_207));
 NAND2x1_ASAP7_75t_SL g211738__8428 (.A(n_8169),
    .B(n_8162),
    .Y(n_8228));
 AO21x2_ASAP7_75t_SL g211739__5526 (.A1(sa23[5]),
    .A2(n_8159),
    .B(n_8161),
    .Y(n_8253));
 AO21x1_ASAP7_75t_SL g211740__6783 (.A1(sa23[5]),
    .A2(n_8157),
    .B(n_8166),
    .Y(n_8276));
 AOI21xp5_ASAP7_75t_SL g211741__3680 (.A1(n_2009),
    .A2(n_8154),
    .B(n_8117),
    .Y(n_8169));
 INVxp67_ASAP7_75t_SL g211742 (.A(n_8254),
    .Y(n_135));
 A2O1A1Ixp33_ASAP7_75t_SL g211743__1617 (.A1(n_8118),
    .A2(n_8141),
    .B(n_2713),
    .C(n_8145),
    .Y(n_8167));
 AO21x1_ASAP7_75t_SL g211744__2802 (.A1(sa23[5]),
    .A2(n_8150),
    .B(n_8163),
    .Y(n_8254));
 NAND2xp5_ASAP7_75t_L g211745__1705 (.A(n_8146),
    .B(n_8143),
    .Y(n_8166));
 A2O1A1Ixp33_ASAP7_75t_SL g211746__5122 (.A1(n_8107),
    .A2(n_8123),
    .B(sa23[5]),
    .C(n_8111),
    .Y(n_8165));
 NAND4xp25_ASAP7_75t_SL g211747__8246 (.A(n_8135),
    .B(n_8128),
    .C(n_8130),
    .D(n_8120),
    .Y(n_8164));
 OAI321xp33_ASAP7_75t_SL g211748__7098 (.A1(n_8136),
    .A2(n_8108),
    .A3(n_2713),
    .B1(n_3351),
    .B2(n_8063),
    .C(n_8126),
    .Y(n_8163));
 A2O1A1Ixp33_ASAP7_75t_SL g211749__6131 (.A1(n_2155),
    .A2(n_8092),
    .B(n_8124),
    .C(sa23[5]),
    .Y(n_8162));
 OAI21xp5_ASAP7_75t_SL g211750__1881 (.A1(n_8134),
    .A2(n_8137),
    .B(n_8153),
    .Y(n_8161));
 OAI211xp5_ASAP7_75t_SL g211751__5115 (.A1(n_1537),
    .A2(n_8125),
    .B(n_8142),
    .C(n_8139),
    .Y(n_8160));
 OAI221xp5_ASAP7_75t_SL g211752__7482 (.A1(n_8081),
    .A2(n_2156),
    .B1(n_8106),
    .B2(n_2261),
    .C(n_8144),
    .Y(n_8159));
 OAI211xp5_ASAP7_75t_SL g211753__4733 (.A1(n_2647),
    .A2(n_8098),
    .B(n_8148),
    .C(n_8132),
    .Y(n_8158));
 OAI211xp5_ASAP7_75t_SL g211754__6161 (.A1(n_2261),
    .A2(n_8072),
    .B(n_8149),
    .C(n_8129),
    .Y(n_8157));
 AOI21xp5_ASAP7_75t_SL g211755__9315 (.A1(n_8133),
    .A2(n_8119),
    .B(n_8151),
    .Y(n_8156));
 AOI21xp5_ASAP7_75t_SL g211756__9945 (.A1(n_8133),
    .A2(sa23[0]),
    .B(n_8127),
    .Y(n_8155));
 OAI211xp5_ASAP7_75t_SL g211757__2883 (.A1(n_7976),
    .A2(n_8099),
    .B(n_8138),
    .C(n_8110),
    .Y(n_8154));
 AOI22xp33_ASAP7_75t_SL g211758__2346 (.A1(n_7966),
    .A2(n_8116),
    .B1(n_8048),
    .B2(n_8090),
    .Y(n_8153));
 OAI221xp5_ASAP7_75t_SL g211759__1666 (.A1(n_8122),
    .A2(n_3513),
    .B1(n_8067),
    .B2(n_3351),
    .C(n_8053),
    .Y(n_8152));
 AOI221xp5_ASAP7_75t_L g211760__7410 (.A1(n_8075),
    .A2(n_2012),
    .B1(n_8100),
    .B2(sa23[0]),
    .C(n_2713),
    .Y(n_8151));
 OAI321xp33_ASAP7_75t_L g211761__6417 (.A1(n_8087),
    .A2(n_7954),
    .A3(n_7986),
    .B1(n_2597),
    .B2(n_8070),
    .C(n_8131),
    .Y(n_8150));
 AOI22xp33_ASAP7_75t_SL g211762__5477 (.A1(n_2598),
    .A2(n_8113),
    .B1(n_2648),
    .B2(n_8104),
    .Y(n_8149));
 AOI22xp5_ASAP7_75t_SL g211763__2398 (.A1(n_2155),
    .A2(n_8073),
    .B1(n_2598),
    .B2(n_8105),
    .Y(n_8148));
 OAI221xp5_ASAP7_75t_L g211764__5107 (.A1(n_8019),
    .A2(n_1538),
    .B1(n_8068),
    .B2(n_1537),
    .C(n_7959),
    .Y(n_8147));
 AOI221xp5_ASAP7_75t_L g211765__6260 (.A1(n_7989),
    .A2(n_3469),
    .B1(n_8076),
    .B2(n_3350),
    .C(n_8121),
    .Y(n_8146));
 AOI22xp33_ASAP7_75t_SL g211766__4319 (.A1(n_3493),
    .A2(n_8112),
    .B1(n_3350),
    .B2(n_8078),
    .Y(n_8145));
 AOI22xp33_ASAP7_75t_L g211767__8428 (.A1(n_2598),
    .A2(n_8115),
    .B1(n_2648),
    .B2(n_8069),
    .Y(n_8144));
 OAI331xp33_ASAP7_75t_L g211768__5526 (.A1(n_8079),
    .A2(n_8041),
    .A3(n_1537),
    .B1(n_8060),
    .B2(n_7967),
    .B3(n_1538),
    .C1(n_2704),
    .Y(n_8143));
 OAI21xp5_ASAP7_75t_L g211769__6783 (.A1(n_8086),
    .A2(n_7980),
    .B(n_2598),
    .Y(n_8142));
 A2O1A1Ixp33_ASAP7_75t_R g211770__3680 (.A1(n_1832),
    .A2(n_5375),
    .B(n_8091),
    .C(n_2012),
    .Y(n_8141));
 AOI21xp5_ASAP7_75t_L g211771__1617 (.A1(n_7955),
    .A2(n_3350),
    .B(n_8103),
    .Y(n_8140));
 A2O1A1Ixp33_ASAP7_75t_L g211772__2802 (.A1(n_1916),
    .A2(n_7991),
    .B(n_8065),
    .C(n_2155),
    .Y(n_8139));
 O2A1O1Ixp33_ASAP7_75t_SL g211773__1705 (.A1(n_1835),
    .A2(n_5432),
    .B(n_8088),
    .C(n_8114),
    .Y(n_8138));
 OAI21xp33_ASAP7_75t_L g211774__5122 (.A1(n_1537),
    .A2(n_8064),
    .B(n_2704),
    .Y(n_8137));
 O2A1O1Ixp33_ASAP7_75t_L g211775__8246 (.A1(n_2642),
    .A2(n_7970),
    .B(n_8058),
    .C(n_2012),
    .Y(n_8136));
 OAI21xp33_ASAP7_75t_R g211776__7098 (.A1(n_8085),
    .A2(n_8005),
    .B(n_2598),
    .Y(n_8135));
 AOI31xp33_ASAP7_75t_L g211777__6131 (.A1(n_7988),
    .A2(n_8034),
    .A3(n_8050),
    .B(n_1538),
    .Y(n_8134));
 AO21x1_ASAP7_75t_SL g211778__1881 (.A1(n_8061),
    .A2(n_7966),
    .B(n_2261),
    .Y(n_8132));
 AOI21xp33_ASAP7_75t_L g211779__5115 (.A1(n_8083),
    .A2(n_2262),
    .B(n_8094),
    .Y(n_8131));
 AO21x1_ASAP7_75t_SL g211780__7482 (.A1(n_7966),
    .A2(n_8057),
    .B(n_2261),
    .Y(n_8130));
 OAI21xp33_ASAP7_75t_R g211781__4733 (.A1(n_7980),
    .A2(n_8055),
    .B(n_2155),
    .Y(n_8129));
 A2O1A1Ixp33_ASAP7_75t_L g211782__6161 (.A1(n_1836),
    .A2(n_3919),
    .B(n_8082),
    .C(n_2155),
    .Y(n_8128));
 A2O1A1Ixp33_ASAP7_75t_SL g211783__9315 (.A1(n_8032),
    .A2(n_7950),
    .B(n_3622),
    .C(n_8109),
    .Y(n_8127));
 O2A1O1Ixp33_ASAP7_75t_L g211784__9945 (.A1(n_8027),
    .A2(n_8039),
    .B(n_3493),
    .C(n_8040),
    .Y(n_8126));
 AOI22xp5_ASAP7_75t_SL g211785__2883 (.A1(n_8038),
    .A2(n_8097),
    .B1(sa23[0]),
    .B2(n_8066),
    .Y(n_8125));
 AOI211xp5_ASAP7_75t_SL g211786__2346 (.A1(n_8077),
    .A2(sa23[0]),
    .B(n_8071),
    .C(n_1537),
    .Y(n_8124));
 O2A1O1Ixp33_ASAP7_75t_L g211787__1666 (.A1(n_8028),
    .A2(n_7961),
    .B(sa23[0]),
    .C(n_2038),
    .Y(n_8133));
 OAI21xp33_ASAP7_75t_L g211788__7410 (.A1(n_8020),
    .A2(n_7954),
    .B(n_2598),
    .Y(n_8123));
 NOR2xp33_ASAP7_75t_SL g211789__6417 (.A(n_8089),
    .B(n_7976),
    .Y(n_8122));
 AOI31xp33_ASAP7_75t_L g211790__5477 (.A1(n_8021),
    .A2(n_8004),
    .A3(n_7984),
    .B(n_3513),
    .Y(n_8121));
 A2O1A1Ixp33_ASAP7_75t_L g211791__2398 (.A1(n_2194),
    .A2(n_1824),
    .B(n_8026),
    .C(n_2648),
    .Y(n_8120));
 O2A1O1Ixp33_ASAP7_75t_L g211792__5107 (.A1(n_3526),
    .A2(n_4304),
    .B(n_1836),
    .C(n_8101),
    .Y(n_8119));
 OAI221xp5_ASAP7_75t_L g211793__6260 (.A1(n_7990),
    .A2(n_3459),
    .B1(n_4409),
    .B2(n_1837),
    .C(n_8062),
    .Y(n_8118));
 AOI31xp33_ASAP7_75t_L g211794__4319 (.A1(n_8006),
    .A2(n_8049),
    .A3(n_7975),
    .B(n_3622),
    .Y(n_8117));
 AOI211xp5_ASAP7_75t_SL g211795__8428 (.A1(n_8009),
    .A2(n_1687),
    .B(n_8054),
    .C(n_8001),
    .Y(n_8116));
 OAI221xp5_ASAP7_75t_L g211796__5526 (.A1(n_3458),
    .A2(n_1833),
    .B1(n_2605),
    .B2(n_1823),
    .C(n_8096),
    .Y(n_8115));
 AOI211xp5_ASAP7_75t_L g211797__6783 (.A1(n_4416),
    .A2(n_7953),
    .B(n_8044),
    .C(n_8013),
    .Y(n_8114));
 OAI221xp5_ASAP7_75t_L g211798__3680 (.A1(n_8033),
    .A2(n_7985),
    .B1(n_5529),
    .B2(n_7951),
    .C(n_7996),
    .Y(n_8113));
 OAI211xp5_ASAP7_75t_L g211799__1617 (.A1(n_3481),
    .A2(n_1833),
    .B(n_8084),
    .C(n_7957),
    .Y(n_8112));
 OAI211xp5_ASAP7_75t_SL g211800__2802 (.A1(n_1835),
    .A2(n_3871),
    .B(n_8093),
    .C(n_7975),
    .Y(n_8111));
 OAI311xp33_ASAP7_75t_L g211801__1705 (.A1(n_4406),
    .A2(n_3305),
    .A3(n_1833),
    .B1(n_1838),
    .C1(n_8056),
    .Y(n_8110));
 OAI211xp5_ASAP7_75t_L g211802__5122 (.A1(n_1825),
    .A2(n_3615),
    .B(n_8102),
    .C(n_7965),
    .Y(n_8109));
 AOI211xp5_ASAP7_75t_L g211803__8246 (.A1(n_4416),
    .A2(n_1830),
    .B(n_8095),
    .C(n_7997),
    .Y(n_8108));
 OAI21xp33_ASAP7_75t_SL g211804__7098 (.A1(n_2194),
    .A2(n_7965),
    .B(n_8080),
    .Y(n_8107));
 AOI211xp5_ASAP7_75t_L g211805__6131 (.A1(n_4501),
    .A2(n_1830),
    .B(n_7978),
    .C(n_8059),
    .Y(n_8106));
 OAI221xp5_ASAP7_75t_L g211806__1881 (.A1(n_7994),
    .A2(n_2194),
    .B1(n_3016),
    .B2(n_1825),
    .C(n_8015),
    .Y(n_8105));
 OAI222xp33_ASAP7_75t_SL g211807__5115 (.A1(n_8036),
    .A2(n_2138),
    .B1(n_5453),
    .B2(n_1825),
    .C1(n_3090),
    .C2(n_1837),
    .Y(n_8104));
 AOI321xp33_ASAP7_75t_R g211808__7482 (.A1(n_1750),
    .A2(n_3354),
    .A3(n_1834),
    .B1(n_7964),
    .B2(n_2469),
    .C(n_8024),
    .Y(n_8103));
 AND4x1_ASAP7_75t_L g211809__4733 (.A(n_1838),
    .B(n_7981),
    .C(n_2155),
    .D(sa23[5]),
    .Y(n_8102));
 OAI221xp5_ASAP7_75t_SL g211810__6161 (.A1(n_4428),
    .A2(n_1833),
    .B1(n_3240),
    .B2(n_1825),
    .C(n_7995),
    .Y(n_8101));
 OAI211xp5_ASAP7_75t_R g211811__9315 (.A1(n_1831),
    .A2(n_4135),
    .B(n_7962),
    .C(n_1826),
    .Y(n_8100));
 OAI211xp5_ASAP7_75t_SL g211812__9945 (.A1(n_1833),
    .A2(n_4447),
    .B(n_8047),
    .C(n_2648),
    .Y(n_8099));
 AOI221xp5_ASAP7_75t_R g211813__2883 (.A1(n_3902),
    .A2(n_1830),
    .B1(n_3901),
    .B2(n_1822),
    .C(n_8046),
    .Y(n_8098));
 AOI211xp5_ASAP7_75t_L g211814__2346 (.A1(n_4052),
    .A2(n_1836),
    .B(n_7967),
    .C(sa23[0]),
    .Y(n_8097));
 AOI221xp5_ASAP7_75t_L g211815__1666 (.A1(n_3982),
    .A2(n_1821),
    .B1(n_2605),
    .B2(n_7953),
    .C(n_7993),
    .Y(n_8096));
 OAI211xp5_ASAP7_75t_R g211816__7410 (.A1(n_2139),
    .A2(n_7951),
    .B(n_8000),
    .C(n_2012),
    .Y(n_8095));
 AOI221xp5_ASAP7_75t_R g211817__6417 (.A1(n_4409),
    .A2(n_7953),
    .B1(n_1822),
    .B2(sa23[4]),
    .C(n_8010),
    .Y(n_8094));
 AOI211xp5_ASAP7_75t_SL g211818__5477 (.A1(n_3265),
    .A2(n_1822),
    .B(n_8007),
    .C(n_3513),
    .Y(n_8093));
 OAI221xp5_ASAP7_75t_L g211819__2398 (.A1(n_5054),
    .A2(n_1837),
    .B1(n_4501),
    .B2(n_1825),
    .C(n_8037),
    .Y(n_8092));
 OAI21xp33_ASAP7_75t_R g211820__5107 (.A1(n_3388),
    .A2(n_7992),
    .B(n_8045),
    .Y(n_8091));
 AOI211xp5_ASAP7_75t_R g211821__6260 (.A1(n_4335),
    .A2(n_1830),
    .B(n_8002),
    .C(n_3351),
    .Y(n_8090));
 OAI211xp5_ASAP7_75t_R g211822__4319 (.A1(n_1835),
    .A2(n_4423),
    .B(n_8003),
    .C(n_7971),
    .Y(n_8089));
 AOI211xp5_ASAP7_75t_SL g211823__8428 (.A1(n_4664),
    .A2(n_1827),
    .B(n_8042),
    .C(n_7977),
    .Y(n_8088));
 OAI211xp5_ASAP7_75t_R g211824__5526 (.A1(n_1835),
    .A2(n_1779),
    .B(n_8008),
    .C(n_2648),
    .Y(n_8087));
 OAI221xp5_ASAP7_75t_SL g211825__6783 (.A1(n_3120),
    .A2(n_1820),
    .B1(n_2194),
    .B2(n_1826),
    .C(n_7970),
    .Y(n_8086));
 OAI221xp5_ASAP7_75t_R g211826__3680 (.A1(n_4700),
    .A2(n_1835),
    .B1(n_1825),
    .B2(n_1617),
    .C(n_7990),
    .Y(n_8085));
 AOI221xp5_ASAP7_75t_L g211827__1617 (.A1(n_3638),
    .A2(n_7953),
    .B1(n_1822),
    .B2(n_1513),
    .C(n_7993),
    .Y(n_8084));
 OAI211xp5_ASAP7_75t_L g211828__2802 (.A1(n_1831),
    .A2(n_4111),
    .B(n_8023),
    .C(n_7999),
    .Y(n_8083));
 OAI221xp5_ASAP7_75t_L g211829__1705 (.A1(n_1779),
    .A2(n_1826),
    .B1(n_3703),
    .B2(n_1821),
    .C(n_7971),
    .Y(n_8082));
 AOI211xp5_ASAP7_75t_SL g211830__5122 (.A1(n_4664),
    .A2(n_1830),
    .B(n_8017),
    .C(n_7972),
    .Y(n_8081));
 AOI211xp5_ASAP7_75t_L g211831__8246 (.A1(n_3912),
    .A2(n_1824),
    .B(n_8025),
    .C(n_2647),
    .Y(n_8080));
 O2A1O1Ixp33_ASAP7_75t_L g211832__7098 (.A1(n_1687),
    .A2(n_1831),
    .B(n_7969),
    .C(n_2341),
    .Y(n_8079));
 OAI221xp5_ASAP7_75t_L g211833__6131 (.A1(n_5138),
    .A2(n_1829),
    .B1(n_5099),
    .B2(n_1821),
    .C(n_7960),
    .Y(n_8078));
 OAI211xp5_ASAP7_75t_L g211834__1881 (.A1(n_1833),
    .A2(n_5426),
    .B(n_7973),
    .C(n_8035),
    .Y(n_8077));
 A2O1A1Ixp33_ASAP7_75t_L g211835__5115 (.A1(n_2469),
    .A2(n_1779),
    .B(n_1837),
    .C(n_8031),
    .Y(n_8076));
 OAI211xp5_ASAP7_75t_L g211836__7482 (.A1(n_1835),
    .A2(n_3266),
    .B(n_7995),
    .C(n_8051),
    .Y(n_8075));
 OAI221xp5_ASAP7_75t_R g211837__4733 (.A1(n_4428),
    .A2(n_7951),
    .B1(n_4603),
    .B2(n_1825),
    .C(n_8014),
    .Y(n_8074));
 OAI211xp5_ASAP7_75t_SL g211838__6161 (.A1(n_1837),
    .A2(n_4097),
    .B(n_7979),
    .C(n_8011),
    .Y(n_8073));
 AOI221xp5_ASAP7_75t_R g211839__9315 (.A1(n_3355),
    .A2(n_1830),
    .B1(n_1822),
    .B2(n_2642),
    .C(n_8012),
    .Y(n_8072));
 AOI211xp5_ASAP7_75t_SL g211840__9945 (.A1(n_4447),
    .A2(n_1827),
    .B(n_8030),
    .C(sa23[0]),
    .Y(n_8071));
 AOI211xp5_ASAP7_75t_L g211841__2883 (.A1(n_4111),
    .A2(n_1822),
    .B(n_8029),
    .C(n_7956),
    .Y(n_8070));
 OAI221xp5_ASAP7_75t_R g211842__2346 (.A1(n_3016),
    .A2(n_1831),
    .B1(n_3119),
    .B2(n_1825),
    .C(n_8016),
    .Y(n_8069));
 AOI221xp5_ASAP7_75t_SL g211843__1666 (.A1(n_5318),
    .A2(n_7952),
    .B1(n_4517),
    .B2(n_1834),
    .C(n_8022),
    .Y(n_8068));
 AOI221xp5_ASAP7_75t_L g211844__7410 (.A1(n_4700),
    .A2(sa23[3]),
    .B1(n_2209),
    .B2(n_1983),
    .C(n_8043),
    .Y(n_8067));
 OAI222xp33_ASAP7_75t_SL g211845__6417 (.A1(n_1833),
    .A2(n_2604),
    .B1(n_5099),
    .B2(n_1820),
    .C1(n_4423),
    .C2(n_1823),
    .Y(n_8066));
 OAI222xp33_ASAP7_75t_L g211846__5477 (.A1(n_1826),
    .A2(n_2160),
    .B1(n_3015),
    .B2(n_1823),
    .C1(n_2733),
    .C2(n_1820),
    .Y(n_8065));
 AOI221xp5_ASAP7_75t_L g211847__2398 (.A1(n_2528),
    .A2(n_1822),
    .B1(n_4335),
    .B2(n_7947),
    .C(n_7949),
    .Y(n_8064));
 AOI221xp5_ASAP7_75t_SL g211848__5107 (.A1(n_4409),
    .A2(n_1821),
    .B1(n_1827),
    .B2(n_2604),
    .C(n_7987),
    .Y(n_8063));
 AOI221xp5_ASAP7_75t_L g211849__6260 (.A1(n_1824),
    .A2(n_2515),
    .B1(n_3647),
    .B2(n_7953),
    .C(n_2012),
    .Y(n_8062));
 AOI211xp5_ASAP7_75t_L g211850__4319 (.A1(n_1836),
    .A2(n_1916),
    .B(n_8052),
    .C(n_8009),
    .Y(n_8061));
 OAI322xp33_ASAP7_75t_L g211851__8428 (.A1(n_3638),
    .A2(n_1835),
    .A3(n_2470),
    .B1(n_4586),
    .B2(n_1823),
    .C1(n_1831),
    .C2(n_2469),
    .Y(n_8060));
 OAI22xp33_ASAP7_75t_R g211852__5526 (.A1(n_3364),
    .A2(n_7992),
    .B1(n_1837),
    .B2(n_1687),
    .Y(n_8059));
 AOI221xp5_ASAP7_75t_R g211853__6783 (.A1(n_1827),
    .A2(n_2515),
    .B1(n_4518),
    .B2(n_1832),
    .C(n_7948),
    .Y(n_8058));
 AOI322xp5_ASAP7_75t_L g211854__3680 (.A1(n_3354),
    .A2(n_3304),
    .A3(n_1822),
    .B1(n_1834),
    .B2(n_4603),
    .C1(n_5053),
    .C2(n_1832),
    .Y(n_8057));
 AOI221xp5_ASAP7_75t_L g211855__1617 (.A1(n_4096),
    .A2(n_1822),
    .B1(n_1828),
    .B2(n_3623),
    .C(n_2156),
    .Y(n_8056));
 OAI321xp33_ASAP7_75t_R g211856__2802 (.A1(n_1835),
    .A2(n_3323),
    .A3(n_2605),
    .B1(n_7951),
    .B2(n_4336),
    .C(n_7958),
    .Y(n_8055));
 AO21x1_ASAP7_75t_SL g211857__1705 (.A1(n_1832),
    .A2(n_3015),
    .B(n_3513),
    .Y(n_8054));
 NAND2xp5_ASAP7_75t_R g211858__5122 (.A(n_2208),
    .B(n_7989),
    .Y(n_8053));
 NOR2xp33_ASAP7_75t_R g211859__8246 (.A(n_3388),
    .B(n_7994),
    .Y(n_8052));
 NOR2xp33_ASAP7_75t_R g211860__7098 (.A(n_7977),
    .B(n_7993),
    .Y(n_8051));
 OR2x2_ASAP7_75t_R g211861__6131 (.A(n_2160),
    .B(n_7992),
    .Y(n_8050));
 OA21x2_ASAP7_75t_R g211862__1881 (.A1(n_1835),
    .A2(n_3912),
    .B(n_8004),
    .Y(n_8049));
 O2A1O1Ixp33_ASAP7_75t_R g211863__5115 (.A1(n_3355),
    .A2(n_3469),
    .B(n_1834),
    .C(n_7968),
    .Y(n_8048));
 A2O1A1Ixp33_ASAP7_75t_L g211864__7482 (.A1(n_1821),
    .A2(n_3364),
    .B(n_7953),
    .C(n_5497),
    .Y(n_8047));
 O2A1O1Ixp33_ASAP7_75t_R g211865__4733 (.A1(n_1820),
    .A2(n_2514),
    .B(n_1826),
    .C(n_3481),
    .Y(n_8046));
 A2O1A1Ixp33_ASAP7_75t_R g211866__6161 (.A1(n_1821),
    .A2(n_2208),
    .B(n_7953),
    .C(n_1517),
    .Y(n_8045));
 OAI21xp33_ASAP7_75t_R g211867__9315 (.A1(n_3106),
    .A2(n_1823),
    .B(n_2598),
    .Y(n_8044));
 NOR2xp33_ASAP7_75t_R g211868__9945 (.A(n_2515),
    .B(n_7994),
    .Y(n_8043));
 OAI21xp33_ASAP7_75t_R g211869__2883 (.A1(n_1823),
    .A2(n_3912),
    .B(n_2262),
    .Y(n_8042));
 O2A1O1Ixp33_ASAP7_75t_R g211870__2346 (.A1(n_1820),
    .A2(n_2208),
    .B(n_1837),
    .C(n_2289),
    .Y(n_8041));
 OA21x2_ASAP7_75t_L g211871__1666 (.A1(n_2605),
    .A2(n_3305),
    .B(n_7989),
    .Y(n_8040));
 OAI21xp33_ASAP7_75t_R g211872__7410 (.A1(n_2515),
    .A2(n_1826),
    .B(n_1838),
    .Y(n_8039));
 A2O1A1Ixp33_ASAP7_75t_R g211873__6417 (.A1(n_1820),
    .A2(n_2193),
    .B(n_7952),
    .C(n_3983),
    .Y(n_8038));
 A2O1A1Ixp33_ASAP7_75t_R g211874__5477 (.A1(n_1820),
    .A2(n_2139),
    .B(n_1824),
    .C(n_4305),
    .Y(n_8037));
 AOI31xp33_ASAP7_75t_SL g211875__2398 (.A1(n_1779),
    .A2(n_2469),
    .A3(n_1820),
    .B(n_1830),
    .Y(n_8036));
 AOI21xp5_ASAP7_75t_SL g211876__5107 (.A1(n_1827),
    .A2(n_2208),
    .B(n_3323),
    .Y(n_8035));
 AOI21xp33_ASAP7_75t_R g211877__6260 (.A1(n_1827),
    .A2(n_3919),
    .B(n_7998),
    .Y(n_8034));
 O2A1O1Ixp33_ASAP7_75t_R g211878__4319 (.A1(n_2605),
    .A2(n_3303),
    .B(n_1832),
    .C(n_7974),
    .Y(n_8033));
 INVxp67_ASAP7_75t_SL g211879 (.A(n_8018),
    .Y(n_8032));
 AOI22xp33_ASAP7_75t_R g211880__8428 (.A1(n_7953),
    .A2(n_4501),
    .B1(n_1820),
    .B2(n_2335),
    .Y(n_8031));
 A2O1A1Ixp33_ASAP7_75t_L g211881__5526 (.A1(n_2340),
    .A2(n_3919),
    .B(n_1821),
    .C(n_7983),
    .Y(n_8030));
 AO21x1_ASAP7_75t_R g211882__6783 (.A1(n_1830),
    .A2(n_3983),
    .B(n_7974),
    .Y(n_8029));
 OAI22xp33_ASAP7_75t_R g211883__3680 (.A1(n_1820),
    .A2(n_5161),
    .B1(n_1823),
    .B2(n_3363),
    .Y(n_8028));
 A2O1A1Ixp33_ASAP7_75t_R g211884__1617 (.A1(n_2159),
    .A2(n_2527),
    .B(n_1833),
    .C(n_7982),
    .Y(n_8027));
 OAI21xp33_ASAP7_75t_L g211885__2802 (.A1(n_1983),
    .A2(n_3266),
    .B(n_7963),
    .Y(n_8026));
 OAI22xp33_ASAP7_75t_R g211886__1705 (.A1(n_3901),
    .A2(n_1837),
    .B1(n_3647),
    .B2(n_1829),
    .Y(n_8025));
 OAI221xp5_ASAP7_75t_L g211887__5122 (.A1(n_1826),
    .A2(sa23[4]),
    .B1(n_3692),
    .B2(n_1983),
    .C(n_3493),
    .Y(n_8024));
 AOI22xp33_ASAP7_75t_R g211888__8246 (.A1(n_1827),
    .A2(n_3107),
    .B1(n_7952),
    .B2(n_3594),
    .Y(n_8023));
 OAI22xp33_ASAP7_75t_R g211889__7098 (.A1(n_3594),
    .A2(n_1826),
    .B1(n_2193),
    .B2(n_1831),
    .Y(n_8022));
 AOI22xp33_ASAP7_75t_L g211890__6131 (.A1(n_1821),
    .A2(n_4447),
    .B1(n_2290),
    .B2(n_7952),
    .Y(n_8021));
 OAI32xp33_ASAP7_75t_L g211891__1881 (.A1(n_1833),
    .A2(n_3303),
    .A3(n_1617),
    .B1(n_1820),
    .B2(n_5140),
    .Y(n_8020));
 AOI22xp33_ASAP7_75t_R g211892__5115 (.A1(n_5374),
    .A2(n_1824),
    .B1(n_3912),
    .B2(n_1830),
    .Y(n_8019));
 OAI22xp5_ASAP7_75t_R g211893__7482 (.A1(n_1829),
    .A2(n_4428),
    .B1(n_1835),
    .B2(n_3703),
    .Y(n_8018));
 OAI22xp33_ASAP7_75t_R g211894__4733 (.A1(n_4052),
    .A2(n_1826),
    .B1(n_4416),
    .B2(n_1823),
    .Y(n_8017));
 AOI32xp33_ASAP7_75t_R g211895__6161 (.A1(n_7952),
    .A2(n_2159),
    .A3(n_1513),
    .B1(n_1836),
    .B2(n_2209),
    .Y(n_8016));
 AOI22xp5_ASAP7_75t_L g211896__9315 (.A1(n_3624),
    .A2(n_1834),
    .B1(n_2289),
    .B2(n_1824),
    .Y(n_8015));
 AOI22xp33_ASAP7_75t_R g211897__9945 (.A1(n_1836),
    .A2(n_4429),
    .B1(n_1687),
    .B2(n_1830),
    .Y(n_8014));
 OAI22xp33_ASAP7_75t_L g211898__2883 (.A1(n_3480),
    .A2(n_1833),
    .B1(n_3589),
    .B2(n_1835),
    .Y(n_8013));
 OAI22xp33_ASAP7_75t_R g211899__2346 (.A1(n_1837),
    .A2(n_3364),
    .B1(n_1826),
    .B2(n_3436),
    .Y(n_8012));
 AOI22xp33_ASAP7_75t_R g211900__1666 (.A1(n_1830),
    .A2(n_4429),
    .B1(n_3303),
    .B2(n_1822),
    .Y(n_8011));
 OAI221xp5_ASAP7_75t_R g211901__7410 (.A1(n_3265),
    .A2(n_1835),
    .B1(n_1751),
    .B2(n_1821),
    .C(n_2155),
    .Y(n_8010));
 INVxp67_ASAP7_75t_R g211902 (.A(n_8007),
    .Y(n_8008));
 INVxp33_ASAP7_75t_R g211903 (.A(n_8005),
    .Y(n_8006));
 INVxp67_ASAP7_75t_R g211904 (.A(n_8002),
    .Y(n_8003));
 INVxp67_ASAP7_75t_R g211905 (.A(n_8000),
    .Y(n_8001));
 INVxp33_ASAP7_75t_R g211906 (.A(n_7998),
    .Y(n_7999));
 INVxp33_ASAP7_75t_R g211907 (.A(n_7996),
    .Y(n_7997));
 INVxp33_ASAP7_75t_R g211908 (.A(n_7990),
    .Y(n_7991));
 NAND2xp33_ASAP7_75t_R g211909__6417 (.A(n_5432),
    .B(n_1832),
    .Y(n_7988));
 NOR2xp33_ASAP7_75t_L g211910__5477 (.A(n_1833),
    .B(n_5453),
    .Y(n_7987));
 NOR2xp33_ASAP7_75t_R g211911__2398 (.A(n_1825),
    .B(n_4305),
    .Y(n_7986));
 NOR2xp33_ASAP7_75t_R g211912__5107 (.A(n_2604),
    .B(n_1830),
    .Y(n_7985));
 NAND2xp33_ASAP7_75t_R g211913__6260 (.A(n_7953),
    .B(n_1517),
    .Y(n_7984));
 NAND2xp5_ASAP7_75t_R g211914__4319 (.A(n_1836),
    .B(n_3090),
    .Y(n_7983));
 NAND2xp5_ASAP7_75t_L g211915__8428 (.A(n_1824),
    .B(n_3015),
    .Y(n_7982));
 NAND2xp33_ASAP7_75t_R g211916__5526 (.A(n_3455),
    .B(n_7952),
    .Y(n_7981));
 NOR2xp33_ASAP7_75t_R g211917__6783 (.A(n_2515),
    .B(n_1823),
    .Y(n_8009));
 NOR2xp33_ASAP7_75t_L g211918__3680 (.A(n_1833),
    .B(n_4665),
    .Y(n_8007));
 NOR2xp33_ASAP7_75t_R g211919__1617 (.A(n_1823),
    .B(n_5425),
    .Y(n_8005));
 NAND2xp33_ASAP7_75t_R g211920__2802 (.A(n_1832),
    .B(n_3594),
    .Y(n_8004));
 NOR2xp33_ASAP7_75t_R g211921__1705 (.A(n_1829),
    .B(n_3469),
    .Y(n_8002));
 NAND2xp33_ASAP7_75t_R g211922__5122 (.A(n_1836),
    .B(n_3679),
    .Y(n_8000));
 NOR2xp33_ASAP7_75t_R g211923__8246 (.A(n_3455),
    .B(n_1835),
    .Y(n_7998));
 NAND2xp5_ASAP7_75t_R g211924__7098 (.A(n_1827),
    .B(n_4429),
    .Y(n_7996));
 NAND2xp5_ASAP7_75t_R g211925__6131 (.A(n_1822),
    .B(n_4665),
    .Y(n_7995));
 NAND2xp5_ASAP7_75t_L g211926__1881 (.A(n_2469),
    .B(n_1830),
    .Y(n_7994));
 AND2x2_ASAP7_75t_R g211927__5115 (.A(n_2470),
    .B(n_1828),
    .Y(n_7993));
 NAND2xp5_ASAP7_75t_R g211928__7482 (.A(n_2527),
    .B(n_7952),
    .Y(n_7992));
 NAND2xp5_ASAP7_75t_R g211929__4733 (.A(n_1832),
    .B(n_2527),
    .Y(n_7990));
 NOR2xp33_ASAP7_75t_L g211930__6161 (.A(n_1823),
    .B(n_3351),
    .Y(n_7989));
 INVxp67_ASAP7_75t_SL g211931 (.A(n_7978),
    .Y(n_7979));
 INVxp67_ASAP7_75t_R g211932 (.A(n_7972),
    .Y(n_7973));
 INVxp67_ASAP7_75t_R g211933 (.A(n_7968),
    .Y(n_7969));
 INVxp33_ASAP7_75t_R g211935 (.A(n_7965),
    .Y(n_7964));
 AOI22xp33_ASAP7_75t_L g211936__9315 (.A1(n_1820),
    .A2(n_3481),
    .B1(n_2138),
    .B2(n_2341),
    .Y(n_7963));
 AOI22xp33_ASAP7_75t_R g211937__9945 (.A1(n_1821),
    .A2(n_3679),
    .B1(sa23[3]),
    .B2(n_1750),
    .Y(n_7962));
 NOR2xp33_ASAP7_75t_R g211938__2883 (.A(n_1833),
    .B(n_3589),
    .Y(n_7961));
 NAND2xp33_ASAP7_75t_R g211939__2346 (.A(n_1836),
    .B(n_4135),
    .Y(n_7960));
 OAI211xp5_ASAP7_75t_R g211940__1666 (.A1(n_2724),
    .A2(n_2528),
    .B(n_1537),
    .C(n_1821),
    .Y(n_7959));
 AO21x1_ASAP7_75t_R g211941__7410 (.A1(n_2193),
    .A2(n_1750),
    .B(n_1825),
    .Y(n_7958));
 OAI21xp33_ASAP7_75t_R g211942__6417 (.A1(n_1688),
    .A2(n_2160),
    .B(n_1836),
    .Y(n_7957));
 AOI21xp33_ASAP7_75t_R g211943__5477 (.A1(n_2527),
    .A2(n_1916),
    .B(n_1825),
    .Y(n_7956));
 OAI22xp33_ASAP7_75t_R g211944__2398 (.A1(n_4744),
    .A2(n_1821),
    .B1(n_5368),
    .B2(n_1820),
    .Y(n_7955));
 AND2x2_ASAP7_75t_L g211945__5107 (.A(n_1830),
    .B(n_5374),
    .Y(n_7980));
 NOR2xp33_ASAP7_75t_SL g211946__6260 (.A(n_1826),
    .B(n_4336),
    .Y(n_7978));
 NOR2xp33_ASAP7_75t_R g211947__4319 (.A(n_2289),
    .B(n_1833),
    .Y(n_7977));
 AOI21xp5_ASAP7_75t_R g211948__8428 (.A1(n_4305),
    .A2(n_1687),
    .B(n_7951),
    .Y(n_7976));
 OAI21xp5_ASAP7_75t_R g211949__5526 (.A1(n_2138),
    .A2(n_2528),
    .B(n_1827),
    .Y(n_7975));
 NOR2xp33_ASAP7_75t_L g211950__6783 (.A(n_1837),
    .B(n_3305),
    .Y(n_7974));
 AOI21xp5_ASAP7_75t_L g211951__3680 (.A1(n_2527),
    .A2(n_3363),
    .B(n_1835),
    .Y(n_7972));
 OAI21xp33_ASAP7_75t_R g211952__1617 (.A1(n_2515),
    .A2(n_2528),
    .B(n_1832),
    .Y(n_7971));
 NAND2xp5_ASAP7_75t_R g211953__2802 (.A(n_1822),
    .B(n_4305),
    .Y(n_7970));
 NOR2xp33_ASAP7_75t_L g211954__1705 (.A(n_1823),
    .B(n_3589),
    .Y(n_7968));
 NOR2xp33_ASAP7_75t_R g211955__5122 (.A(n_1829),
    .B(n_3870),
    .Y(n_7967));
 NAND2xp5_ASAP7_75t_L g211956__8246 (.A(n_1827),
    .B(n_5528),
    .Y(n_7966));
 NAND2xp5_ASAP7_75t_L g211957__7098 (.A(n_1836),
    .B(n_3016),
    .Y(n_1838));
 NAND2xp5_ASAP7_75t_R g211958__6131 (.A(n_1832),
    .B(n_3266),
    .Y(n_7965));
 INVx2_ASAP7_75t_R g211971 (.A(n_1836),
    .Y(n_1837));
 INVx2_ASAP7_75t_SL g211977 (.A(n_1836),
    .Y(n_1835));
 INVx1_ASAP7_75t_SL g211984 (.A(n_1835),
    .Y(n_1834));
 INVx1_ASAP7_75t_SL g212003 (.A(n_1830),
    .Y(n_1831));
 INVx2_ASAP7_75t_SL g212006 (.A(n_1833),
    .Y(n_1830));
 INVx2_ASAP7_75t_L g212007 (.A(n_1833),
    .Y(n_1832));
 INVxp67_ASAP7_75t_R g212015 (.A(n_1828),
    .Y(n_1829));
 INVx2_ASAP7_75t_SL g212020 (.A(n_1826),
    .Y(n_1827));
 INVx2_ASAP7_75t_SL g212024 (.A(n_7953),
    .Y(n_1826));
 INVx1_ASAP7_75t_SL g212027 (.A(n_7953),
    .Y(n_1825));
 BUFx3_ASAP7_75t_L g212036 (.A(n_1828),
    .Y(n_7953));
 NOR2xp33_ASAP7_75t_R g212037__1881 (.A(n_1821),
    .B(n_5497),
    .Y(n_7954));
 AND2x2_ASAP7_75t_SL g212038__5115 (.A(sa23[6]),
    .B(n_1983),
    .Y(n_1836));
 OR2x4_ASAP7_75t_SL g212039__7482 (.A(sa23[6]),
    .B(sa23[3]),
    .Y(n_1833));
 AND2x2_ASAP7_75t_SL g212040__4733 (.A(sa23[6]),
    .B(sa23[3]),
    .Y(n_1828));
 INVx1_ASAP7_75t_SL g212045 (.A(n_1822),
    .Y(n_7951));
 BUFx2_ASAP7_75t_L g212051 (.A(n_7952),
    .Y(n_1822));
 INVx2_ASAP7_75t_SL g212060 (.A(n_7952),
    .Y(n_1823));
 INVxp67_ASAP7_75t_SL g212061 (.A(n_1823),
    .Y(n_1824));
 A2O1A1Ixp33_ASAP7_75t_R g212065__6161 (.A1(sa23[3]),
    .A2(n_4056),
    .B(n_5357),
    .C(n_1820),
    .Y(n_7950));
 NOR2xp33_ASAP7_75t_R g212066__9315 (.A(n_1821),
    .B(n_3871),
    .Y(n_7949));
 OA21x2_ASAP7_75t_R g212067__9945 (.A1(n_2335),
    .A2(n_3305),
    .B(n_1821),
    .Y(n_7948));
 O2A1O1Ixp33_ASAP7_75t_R g212068__2883 (.A1(n_1983),
    .A2(n_2470),
    .B(n_2334),
    .C(n_1820),
    .Y(n_7947));
 AND2x2_ASAP7_75t_SL g212069__2346 (.A(n_7946),
    .B(sa23[3]),
    .Y(n_7952));
 INVx2_ASAP7_75t_L g212083 (.A(n_1821),
    .Y(n_1820));
 BUFx2_ASAP7_75t_L g212090 (.A(sa23[6]),
    .Y(n_1821));
 INVxp67_ASAP7_75t_L g212091 (.A(sa23[6]),
    .Y(n_7946));
 XNOR2xp5_ASAP7_75t_L g212099__1666 (.A(n_7610),
    .B(n_7943),
    .Y(n_7945));
 INVxp67_ASAP7_75t_SL g212105 (.A(n_8277),
    .Y(n_341));
 XNOR2xp5_ASAP7_75t_L g212107__7410 (.A(n_7931),
    .B(n_1800),
    .Y(n_7943));
 OAI21x1_ASAP7_75t_SL g212108__6417 (.A1(n_7932),
    .A2(n_1917),
    .B(n_7926),
    .Y(n_8277));
 OAI21x1_ASAP7_75t_SL g212112__5477 (.A1(n_7921),
    .A2(n_1917),
    .B(n_7925),
    .Y(n_8256));
 NAND3xp33_ASAP7_75t_SL g212117__2398 (.A(n_7904),
    .B(n_7935),
    .C(n_7888),
    .Y(n_8293));
 OAI21x1_ASAP7_75t_SL g212118__5107 (.A1(n_7927),
    .A2(n_1917),
    .B(n_7936),
    .Y(n_8329));
 AO211x2_ASAP7_75t_SL g212119__6260 (.A1(n_2694),
    .A2(n_7916),
    .B(n_7924),
    .C(n_7911),
    .Y(n_8330));
 OAI21x1_ASAP7_75t_SL g212120__4319 (.A1(n_7923),
    .A2(n_1917),
    .B(n_7922),
    .Y(n_8331));
 AOI221x1_ASAP7_75t_SL g212122__8428 (.A1(n_7872),
    .A2(n_3590),
    .B1(n_7907),
    .B2(n_2711),
    .C(n_7912),
    .Y(n_7936));
 A2O1A1Ixp33_ASAP7_75t_SL g212123__5526 (.A1(n_7898),
    .A2(n_7853),
    .B(n_7863),
    .C(sa20[5]),
    .Y(n_7935));
 OR3x2_ASAP7_75t_SL g212125__6783 (.A(n_7914),
    .B(n_7903),
    .C(n_7919),
    .Y(n_8255));
 AOI221xp5_ASAP7_75t_SL g212128__3680 (.A1(n_7857),
    .A2(n_2656),
    .B1(n_7881),
    .B2(n_2685),
    .C(n_7906),
    .Y(n_7932));
 XOR2xp5_ASAP7_75t_L g212129__1617 (.A(n_8274),
    .B(n_8266),
    .Y(n_7931));
 NAND4xp75_ASAP7_75t_SL g212130__2802 (.A(n_7915),
    .B(n_7900),
    .C(n_7790),
    .D(n_7846),
    .Y(n_8226));
 AO21x2_ASAP7_75t_SL g212131__1705 (.A1(n_1917),
    .A2(n_7913),
    .B(n_7905),
    .Y(n_8229));
 AOI21xp5_ASAP7_75t_SL g212136__5122 (.A1(n_7892),
    .A2(n_8179),
    .B(n_7917),
    .Y(n_7927));
 NAND4xp75_ASAP7_75t_SL g212137__8246 (.A(n_7701),
    .B(n_7697),
    .C(n_7893),
    .D(n_7844),
    .Y(n_8290));
 AO221x1_ASAP7_75t_SL g212138__7098 (.A1(n_7896),
    .A2(sa10[5]),
    .B1(n_7114),
    .B2(n_7652),
    .C(n_7765),
    .Y(n_8250));
 AO21x1_ASAP7_75t_SL g212139__6131 (.A1(n_7794),
    .A2(n_7871),
    .B(n_7908),
    .Y(n_8322));
 AND2x2_ASAP7_75t_SL g212140__1881 (.A(n_7901),
    .B(n_7909),
    .Y(n_7926));
 AOI21xp5_ASAP7_75t_SL g212141__5115 (.A1(n_7883),
    .A2(n_7860),
    .B(n_7918),
    .Y(n_7925));
 NAND3xp33_ASAP7_75t_SL g212142__7482 (.A(n_7877),
    .B(n_7891),
    .C(n_7889),
    .Y(n_7924));
 AOI221xp5_ASAP7_75t_SL g212143__4733 (.A1(n_7876),
    .A2(n_2284),
    .B1(n_7838),
    .B2(n_2685),
    .C(n_7902),
    .Y(n_7923));
 AOI221x1_ASAP7_75t_SL g212144__6161 (.A1(n_7854),
    .A2(n_3462),
    .B1(n_2694),
    .B2(n_7887),
    .C(n_7873),
    .Y(n_7922));
 AND4x1_ASAP7_75t_SL g212145__9315 (.A(n_7897),
    .B(n_7885),
    .C(n_7852),
    .D(n_7861),
    .Y(n_7921));
 OAI221xp5_ASAP7_75t_SL g212147__9945 (.A1(n_7705),
    .A2(n_7878),
    .B1(n_7733),
    .B2(n_3442),
    .C(n_7761),
    .Y(n_7919));
 AO22x1_ASAP7_75t_SL g212148__2883 (.A1(n_3384),
    .A2(n_7858),
    .B1(n_3462),
    .B2(n_7818),
    .Y(n_7918));
 A2O1A1Ixp33_ASAP7_75t_SL g212149__2346 (.A1(n_7810),
    .A2(n_7717),
    .B(n_2657),
    .C(n_7895),
    .Y(n_7917));
 OAI21xp5_ASAP7_75t_SL g212150__1666 (.A1(sa20[0]),
    .A2(n_7865),
    .B(n_7870),
    .Y(n_7916));
 OA332x1_ASAP7_75t_SL g212151__7410 (.A1(n_6140),
    .A2(n_7744),
    .A3(n_5316),
    .B1(n_5998),
    .B2(n_7791),
    .B3(n_5085),
    .C1(n_6657),
    .C2(n_7664),
    .Y(n_7915));
 AOI221xp5_ASAP7_75t_SL g212152__6417 (.A1(n_7806),
    .A2(n_8179),
    .B1(n_7859),
    .B2(n_1923),
    .C(n_2710),
    .Y(n_7914));
 OAI321xp33_ASAP7_75t_SL g212153__5477 (.A1(n_7698),
    .A2(n_7769),
    .A3(n_7770),
    .B1(n_7695),
    .B2(n_7845),
    .C(n_7884),
    .Y(n_7913));
 O2A1O1Ixp33_ASAP7_75t_SL g212154__2398 (.A1(n_1724),
    .A2(n_1809),
    .B(n_12816),
    .C(n_3383),
    .Y(n_7912));
 A2O1A1Ixp33_ASAP7_75t_SL g212155__5107 (.A1(n_7706),
    .A2(n_7800),
    .B(n_3479),
    .C(n_7886),
    .Y(n_7911));
 AO21x2_ASAP7_75t_SL g212156__6260 (.A1(sa10[5]),
    .A2(n_7787),
    .B(n_7890),
    .Y(n_8249));
 OAI331xp33_ASAP7_75t_SL g212158__4319 (.A1(n_7757),
    .A2(n_7793),
    .A3(n_7795),
    .B1(n_1923),
    .B2(n_7767),
    .B3(n_7824),
    .C1(n_2711),
    .Y(n_7909));
 OAI322xp33_ASAP7_75t_SL g212159__8428 (.A1(n_5457),
    .A2(n_4708),
    .A3(n_7686),
    .B1(n_7804),
    .B2(n_5314),
    .C1(n_6874),
    .C2(n_7660),
    .Y(n_7908));
 OAI22xp5_ASAP7_75t_SL g212160__5526 (.A1(n_1923),
    .A2(n_7815),
    .B1(n_8179),
    .B2(n_7855),
    .Y(n_7907));
 A2O1A1Ixp33_ASAP7_75t_SL g212161__6783 (.A1(n_7717),
    .A2(n_7823),
    .B(n_2233),
    .C(n_7874),
    .Y(n_7906));
 OAI211xp5_ASAP7_75t_SL g212162__3680 (.A1(n_3473),
    .A2(n_7822),
    .B(n_7882),
    .C(n_7833),
    .Y(n_7905));
 AOI211xp5_ASAP7_75t_SL g212163__1617 (.A1(n_7831),
    .A2(n_3472),
    .B(n_7812),
    .C(n_7869),
    .Y(n_7904));
 OAI221xp5_ASAP7_75t_SL g212164__2802 (.A1(n_7834),
    .A2(n_7784),
    .B1(n_7796),
    .B2(n_3473),
    .C(n_7880),
    .Y(n_7903));
 OAI22xp5_ASAP7_75t_SL g212165__1705 (.A1(n_2233),
    .A2(n_7817),
    .B1(n_2657),
    .B2(n_7866),
    .Y(n_7902));
 AOI22xp33_ASAP7_75t_SL g212166__5122 (.A1(n_3384),
    .A2(n_7864),
    .B1(n_3590),
    .B2(n_7819),
    .Y(n_7901));
 AO221x1_ASAP7_75t_SL g212167__8246 (.A1(n_4025),
    .A2(n_1449),
    .B1(n_7803),
    .B2(n_7676),
    .C(sa10[5]),
    .Y(n_7900));
 AO21x1_ASAP7_75t_SL g212168__7098 (.A1(sa10[5]),
    .A2(n_7771),
    .B(n_7894),
    .Y(n_8274));
 OAI21xp33_ASAP7_75t_R g212170__6131 (.A1(n_7681),
    .A2(n_7847),
    .B(n_1888),
    .Y(n_7898));
 A2O1A1Ixp33_ASAP7_75t_R g212171__1881 (.A1(n_1810),
    .A2(n_4390),
    .B(n_7827),
    .C(n_2656),
    .Y(n_7897));
 NAND3xp33_ASAP7_75t_SL g212172__5115 (.A(n_7821),
    .B(n_7781),
    .C(n_7637),
    .Y(n_7896));
 A2O1A1Ixp33_ASAP7_75t_SL g212173__7482 (.A1(n_2013),
    .A2(n_7710),
    .B(n_7809),
    .C(n_2232),
    .Y(n_7895));
 NAND4xp25_ASAP7_75t_SL g212174__4733 (.A(n_7690),
    .B(n_7743),
    .C(n_7680),
    .D(n_7687),
    .Y(n_7894));
 OA211x2_ASAP7_75t_SL g212175__6161 (.A1(n_7673),
    .A2(n_6646),
    .B(n_7843),
    .C(n_7848),
    .Y(n_7893));
 OAI321xp33_ASAP7_75t_SL g212176__9315 (.A1(n_7647),
    .A2(n_7745),
    .A3(n_7775),
    .B1(n_2613),
    .B2(n_7712),
    .C(n_7811),
    .Y(n_7892));
 OAI21xp33_ASAP7_75t_L g212177__9945 (.A1(n_7724),
    .A2(n_7828),
    .B(n_3472),
    .Y(n_7891));
 OAI21xp5_ASAP7_75t_SL g212178__2883 (.A1(n_7645),
    .A2(n_7617),
    .B(n_7867),
    .Y(n_7890));
 AO21x2_ASAP7_75t_SL g212179__2346 (.A1(sa10[5]),
    .A2(n_7836),
    .B(n_7850),
    .Y(n_8321));
 AOI21xp33_ASAP7_75t_L g212180__1666 (.A1(n_7839),
    .A2(n_3462),
    .B(n_7875),
    .Y(n_7889));
 OAI221xp5_ASAP7_75t_L g212181__7410 (.A1(n_7832),
    .A2(sa20[0]),
    .B1(n_4139),
    .B2(n_7712),
    .C(n_7825),
    .Y(n_7888));
 A2O1A1Ixp33_ASAP7_75t_SL g212182__6417 (.A1(n_2863),
    .A2(n_7708),
    .B(n_7816),
    .C(n_7862),
    .Y(n_7887));
 A2O1A1Ixp33_ASAP7_75t_L g212183__5477 (.A1(n_1807),
    .A2(n_4330),
    .B(n_7820),
    .C(n_3443),
    .Y(n_7886));
 A2O1A1Ixp33_ASAP7_75t_L g212184__2398 (.A1(n_2518),
    .A2(n_7704),
    .B(n_7829),
    .C(n_2284),
    .Y(n_7885));
 O2A1O1Ixp33_ASAP7_75t_L g212185__5107 (.A1(n_1805),
    .A2(n_1784),
    .B(n_7813),
    .C(n_7856),
    .Y(n_7884));
 AOI221xp5_ASAP7_75t_L g212186__6260 (.A1(n_1792),
    .A2(n_7703),
    .B1(n_7729),
    .B2(sa20[0]),
    .C(n_7789),
    .Y(n_7883));
 AOI22xp5_ASAP7_75t_SL g212187__4319 (.A1(n_3443),
    .A2(n_7837),
    .B1(n_3538),
    .B2(n_7801),
    .Y(n_7882));
 OAI222xp33_ASAP7_75t_SL g212188__8428 (.A1(n_7760),
    .A2(n_2106),
    .B1(n_5454),
    .B2(n_1806),
    .C1(n_3149),
    .C2(n_7658),
    .Y(n_7881));
 AOI22xp5_ASAP7_75t_SL g212189__5526 (.A1(n_3538),
    .A2(n_7814),
    .B1(n_3478),
    .B2(n_7826),
    .Y(n_7880));
 OAI211xp5_ASAP7_75t_R g212191__6783 (.A1(n_2499),
    .A2(n_7723),
    .B(n_7773),
    .C(n_7719),
    .Y(n_7878));
 A2O1A1Ixp33_ASAP7_75t_SL g212192__3680 (.A1(n_7623),
    .A2(n_5100),
    .B(n_7751),
    .C(n_3384),
    .Y(n_7877));
 NAND3xp33_ASAP7_75t_SL g212193__1617 (.A(n_7706),
    .B(n_7738),
    .C(n_7723),
    .Y(n_7876));
 O2A1O1Ixp33_ASAP7_75t_L g212194__2802 (.A1(n_2216),
    .A2(n_7654),
    .B(n_7749),
    .C(n_3537),
    .Y(n_7875));
 OAI21xp33_ASAP7_75t_L g212195__1705 (.A1(n_7734),
    .A2(n_7732),
    .B(n_2284),
    .Y(n_7874));
 AOI21xp5_ASAP7_75t_L g212196__5122 (.A1(n_7742),
    .A2(n_7785),
    .B(n_3383),
    .Y(n_7873));
 OR3x1_ASAP7_75t_SL g212197__8246 (.A(n_7754),
    .B(n_7695),
    .C(n_7696),
    .Y(n_7872));
 NAND5xp2_ASAP7_75t_SL g212198__7098 (.A(n_7633),
    .B(n_7642),
    .C(n_7691),
    .D(n_7650),
    .E(n_7631),
    .Y(n_7871));
 OAI221xp5_ASAP7_75t_SL g212199__6131 (.A1(n_7709),
    .A2(n_3504),
    .B1(n_4378),
    .B2(n_7658),
    .C(n_7802),
    .Y(n_7870));
 AOI321xp33_ASAP7_75t_R g212200__1881 (.A1(n_1718),
    .A2(n_1818),
    .A3(n_3348),
    .B1(n_7711),
    .B2(n_2452),
    .C(n_7746),
    .Y(n_7869));
 AOI22xp33_ASAP7_75t_SL g212202__7482 (.A1(n_7756),
    .A2(n_6170),
    .B1(n_6060),
    .B2(n_1339),
    .Y(n_7867));
 AOI221xp5_ASAP7_75t_SL g212203__4733 (.A1(n_3149),
    .A2(n_1808),
    .B1(n_2988),
    .B2(n_1807),
    .C(n_7851),
    .Y(n_7866));
 AO21x2_ASAP7_75t_SL g212204__6161 (.A1(sa10[5]),
    .A2(n_7748),
    .B(n_7849),
    .Y(n_8320));
 AOI221xp5_ASAP7_75t_L g212205__9315 (.A1(n_4400),
    .A2(n_7657),
    .B1(n_5382),
    .B2(n_1810),
    .C(n_7776),
    .Y(n_7865));
 A2O1A1Ixp33_ASAP7_75t_SL g212206__9945 (.A1(n_2452),
    .A2(n_4329),
    .B(n_7658),
    .C(n_7808),
    .Y(n_7864));
 NOR4xp25_ASAP7_75t_R g212207__2883 (.A(n_7702),
    .B(n_7741),
    .C(n_7711),
    .D(n_2233),
    .Y(n_7863));
 NAND2xp5_ASAP7_75t_SL g212208__2346 (.A(n_7797),
    .B(n_7799),
    .Y(n_7862));
 OAI211xp5_ASAP7_75t_L g212209__1666 (.A1(n_3271),
    .A2(n_1817),
    .B(n_7805),
    .C(n_2232),
    .Y(n_7861));
 OAI211xp5_ASAP7_75t_L g212210__7410 (.A1(n_2105),
    .A2(n_7654),
    .B(n_7840),
    .C(n_7721),
    .Y(n_7860));
 OAI211xp5_ASAP7_75t_SL g212211__6417 (.A1(n_1812),
    .A2(n_1792),
    .B(n_7763),
    .C(n_7722),
    .Y(n_7859));
 OAI21xp33_ASAP7_75t_L g212212__5477 (.A1(n_7653),
    .A2(n_5454),
    .B(n_7798),
    .Y(n_7858));
 OAI211xp5_ASAP7_75t_L g212213__2398 (.A1(n_1814),
    .A2(n_5516),
    .B(n_7830),
    .C(n_7721),
    .Y(n_7857));
 NOR3xp33_ASAP7_75t_L g212214__5107 (.A(n_7731),
    .B(n_7702),
    .C(n_7768),
    .Y(n_7856));
 AOI21xp5_ASAP7_75t_R g212215__6260 (.A1(n_5381),
    .A2(n_1813),
    .B(n_7807),
    .Y(n_7855));
 OAI221xp5_ASAP7_75t_R g212216__4319 (.A1(n_4392),
    .A2(n_1817),
    .B1(n_4417),
    .B2(n_1814),
    .C(n_7730),
    .Y(n_7854));
 AOI211xp5_ASAP7_75t_L g212217__8428 (.A1(n_7703),
    .A2(n_2871),
    .B(n_7783),
    .C(n_7779),
    .Y(n_7853));
 OAI211xp5_ASAP7_75t_L g212218__5526 (.A1(n_1805),
    .A2(n_4312),
    .B(n_7835),
    .C(n_7669),
    .Y(n_7852));
 INVxp67_ASAP7_75t_R g212219 (.A(n_7841),
    .Y(n_7851));
 OAI21xp5_ASAP7_75t_SL g212220__6783 (.A1(n_7628),
    .A2(n_7135),
    .B(n_7750),
    .Y(n_7850));
 A2O1A1Ixp33_ASAP7_75t_SL g212221__3680 (.A1(n_7618),
    .A2(n_7634),
    .B(n_2698),
    .C(n_7759),
    .Y(n_7849));
 A2O1A1Ixp33_ASAP7_75t_SL g212222__1617 (.A1(n_7659),
    .A2(n_4729),
    .B(n_7688),
    .C(n_8180),
    .Y(n_7848));
 OAI211xp5_ASAP7_75t_R g212223__2802 (.A1(n_1809),
    .A2(n_4417),
    .B(n_7725),
    .C(n_7684),
    .Y(n_7847));
 NAND3xp33_ASAP7_75t_R g212224__1705 (.A(n_7670),
    .B(n_6216),
    .C(n_6070),
    .Y(n_7846));
 OAI211xp5_ASAP7_75t_R g212225__5122 (.A1(n_7653),
    .A2(n_4431),
    .B(n_7782),
    .C(n_2685),
    .Y(n_7845));
 OR4x1_ASAP7_75t_R g212226__8246 (.A(n_3940),
    .B(n_3943),
    .C(n_4156),
    .D(n_7675),
    .Y(n_7844));
 NOR2xp33_ASAP7_75t_SL g212227__7098 (.A(n_7786),
    .B(n_7788),
    .Y(n_7843));
 A2O1A1Ixp33_ASAP7_75t_L g212228__6131 (.A1(sa20[3]),
    .A2(n_2182),
    .B(n_11524),
    .C(n_4695),
    .Y(n_7842));
 A2O1A1Ixp33_ASAP7_75t_L g212229__1881 (.A1(n_2106),
    .A2(n_1819),
    .B(n_7704),
    .C(sa20[4]),
    .Y(n_7841));
 OA211x2_ASAP7_75t_L g212230__5115 (.A1(n_1812),
    .A2(n_1784),
    .B(n_7719),
    .C(n_1888),
    .Y(n_7840));
 OAI211xp5_ASAP7_75t_L g212231__7482 (.A1(n_1806),
    .A2(n_4223),
    .B(n_7780),
    .C(n_7679),
    .Y(n_7839));
 OAI211xp5_ASAP7_75t_R g212232__4733 (.A1(n_7653),
    .A2(n_3911),
    .B(n_7699),
    .C(n_7778),
    .Y(n_7838));
 OAI221xp5_ASAP7_75t_L g212233__6161 (.A1(n_5059),
    .A2(n_1817),
    .B1(n_4515),
    .B2(n_1805),
    .C(n_7764),
    .Y(n_7837));
 NAND3xp33_ASAP7_75t_SL g212234__9315 (.A(n_7689),
    .B(n_7639),
    .C(n_7636),
    .Y(n_7836));
 AOI211xp5_ASAP7_75t_L g212235__9945 (.A1(n_4330),
    .A2(n_1818),
    .B(n_7713),
    .C(n_2686),
    .Y(n_7835));
 OAI221xp5_ASAP7_75t_R g212236__2883 (.A1(n_3463),
    .A2(n_1806),
    .B1(n_4340),
    .B2(n_7653),
    .C(n_3384),
    .Y(n_7834));
 OAI221xp5_ASAP7_75t_R g212237__2346 (.A1(n_5411),
    .A2(n_7653),
    .B1(n_4399),
    .B2(n_1817),
    .C(n_7740),
    .Y(n_7833));
 AOI211xp5_ASAP7_75t_L g212238__1666 (.A1(n_3271),
    .A2(n_1819),
    .B(n_7726),
    .C(n_7718),
    .Y(n_7832));
 A2O1A1Ixp33_ASAP7_75t_L g212239__7410 (.A1(sa20[3]),
    .A2(n_4391),
    .B(n_7638),
    .C(n_7762),
    .Y(n_7831));
 OAI21xp33_ASAP7_75t_R g212240__6417 (.A1(n_2613),
    .A2(n_1810),
    .B(n_7758),
    .Y(n_7830));
 OAI221xp5_ASAP7_75t_R g212241__5477 (.A1(n_4133),
    .A2(n_1812),
    .B1(n_3156),
    .B2(n_1805),
    .C(n_7722),
    .Y(n_7829));
 OAI221xp5_ASAP7_75t_R g212242__2398 (.A1(n_4694),
    .A2(n_7658),
    .B1(n_1805),
    .B2(n_2285),
    .C(n_7709),
    .Y(n_7828));
 OAI221xp5_ASAP7_75t_R g212243__5107 (.A1(n_4132),
    .A2(n_7654),
    .B1(n_3225),
    .B2(n_1805),
    .C(n_7694),
    .Y(n_7827));
 OAI221xp5_ASAP7_75t_SL g212244__6260 (.A1(n_4514),
    .A2(n_1809),
    .B1(n_1817),
    .B2(n_2500),
    .C(n_7716),
    .Y(n_7826));
 AOI221xp5_ASAP7_75t_R g212245__4319 (.A1(n_1804),
    .A2(n_2453),
    .B1(n_3632),
    .B2(n_7662),
    .C(n_5216),
    .Y(n_7825));
 O2A1O1Ixp33_ASAP7_75t_R g212246__8428 (.A1(n_2500),
    .A2(n_7653),
    .B(n_7720),
    .C(n_2344),
    .Y(n_7824));
 AOI322xp5_ASAP7_75t_L g212247__5526 (.A1(n_1819),
    .A2(n_3326),
    .A3(n_2613),
    .B1(n_7657),
    .B2(n_4341),
    .C1(n_3790),
    .C2(n_1804),
    .Y(n_7823));
 NOR3xp33_ASAP7_75t_L g212248__6783 (.A(n_7766),
    .B(n_7724),
    .C(n_7728),
    .Y(n_7822));
 AOI22xp33_ASAP7_75t_L g212249__3680 (.A1(n_7621),
    .A2(n_6550),
    .B1(n_7672),
    .B2(n_5564),
    .Y(n_7821));
 OAI221xp5_ASAP7_75t_L g212250__1617 (.A1(n_3927),
    .A2(n_7658),
    .B1(n_3691),
    .B2(n_1802),
    .C(n_7693),
    .Y(n_7820));
 OAI211xp5_ASAP7_75t_L g212251__2802 (.A1(n_2348),
    .A2(n_7654),
    .B(n_7747),
    .C(n_7727),
    .Y(n_7819));
 OAI221xp5_ASAP7_75t_SL g212252__1705 (.A1(n_7654),
    .A2(n_2989),
    .B1(n_1805),
    .B2(n_2517),
    .C(n_7772),
    .Y(n_7818));
 AOI221xp5_ASAP7_75t_SL g212253__5122 (.A1(n_4037),
    .A2(n_1819),
    .B1(n_1813),
    .B2(n_3299),
    .C(n_7755),
    .Y(n_7817));
 OR3x1_ASAP7_75t_SL g212254__8246 (.A(n_7713),
    .B(n_7774),
    .C(n_7692),
    .Y(n_7816));
 AOI221xp5_ASAP7_75t_SL g212255__7098 (.A1(n_4038),
    .A2(n_1818),
    .B1(n_1810),
    .B2(n_2217),
    .C(n_7752),
    .Y(n_7815));
 AO221x1_ASAP7_75t_SL g212256__6131 (.A1(n_2988),
    .A2(n_1808),
    .B1(n_2182),
    .B2(n_1819),
    .C(n_7739),
    .Y(n_7814));
 AOI221xp5_ASAP7_75t_R g212257__1881 (.A1(n_1810),
    .A2(n_3521),
    .B1(n_3600),
    .B2(n_1818),
    .C(n_7777),
    .Y(n_7813));
 AOI321xp33_ASAP7_75t_R g212258__5115 (.A1(n_4600),
    .A2(n_2384),
    .A3(n_1802),
    .B1(n_4741),
    .B2(n_7623),
    .C(n_3383),
    .Y(n_7812));
 AOI22xp5_ASAP7_75t_L g212259__7482 (.A1(n_5100),
    .A2(n_7662),
    .B1(n_4387),
    .B2(n_7703),
    .Y(n_7811));
 AOI21xp33_ASAP7_75t_R g212260__4733 (.A1(n_4312),
    .A2(n_1813),
    .B(n_7735),
    .Y(n_7810));
 OAI222xp33_ASAP7_75t_SL g212261__6161 (.A1(n_1814),
    .A2(n_2990),
    .B1(n_3124),
    .B2(n_1801),
    .C1(n_1805),
    .C2(n_1607),
    .Y(n_7809));
 AOI222xp33_ASAP7_75t_SL g212262__9315 (.A1(n_1810),
    .A2(sa20[7]),
    .B1(n_4515),
    .B2(n_1807),
    .C1(n_3463),
    .C2(n_1815),
    .Y(n_7808));
 OAI222xp33_ASAP7_75t_L g212263__9945 (.A1(n_3900),
    .A2(n_7653),
    .B1(n_7658),
    .B2(sa20[4]),
    .C1(n_2578),
    .C2(n_1801),
    .Y(n_7807));
 OAI322xp33_ASAP7_75t_L g212264__2883 (.A1(n_4340),
    .A2(n_3756),
    .A3(n_1801),
    .B1(n_2578),
    .B2(n_7654),
    .C1(n_1771),
    .C2(n_1802),
    .Y(n_7806));
 AOI221xp5_ASAP7_75t_L g212265__2346 (.A1(n_1815),
    .A2(sa20[4]),
    .B1(n_4378),
    .B2(n_1807),
    .C(n_7649),
    .Y(n_7805));
 AO221x1_ASAP7_75t_SL g212266__1666 (.A1(n_3940),
    .A2(n_2100),
    .B1(n_3891),
    .B2(n_2092),
    .C(n_7674),
    .Y(n_7804));
 OAI321xp33_ASAP7_75t_SL g212267__7410 (.A1(n_4356),
    .A2(n_3288),
    .A3(n_2430),
    .B1(n_1551),
    .B2(n_4062),
    .C(n_7682),
    .Y(n_7803));
 AOI221xp5_ASAP7_75t_L g212268__6417 (.A1(n_3721),
    .A2(n_1807),
    .B1(n_2517),
    .B2(n_1815),
    .C(n_1888),
    .Y(n_7802));
 OAI221xp5_ASAP7_75t_R g212269__5477 (.A1(n_5174),
    .A2(n_1802),
    .B1(n_4430),
    .B2(n_1805),
    .C(n_7792),
    .Y(n_7801));
 AOI322xp5_ASAP7_75t_L g212270__2398 (.A1(n_3300),
    .A2(n_7657),
    .A3(n_3348),
    .B1(n_1818),
    .B2(n_4401),
    .C1(n_5060),
    .C2(n_1810),
    .Y(n_7800));
 AOI221xp5_ASAP7_75t_L g212271__5107 (.A1(n_3720),
    .A2(n_1807),
    .B1(n_3899),
    .B2(n_1813),
    .C(sa20[0]),
    .Y(n_7799));
 AOI221xp5_ASAP7_75t_L g212272__6260 (.A1(n_4378),
    .A2(n_1802),
    .B1(n_1807),
    .B2(n_2613),
    .C(n_7678),
    .Y(n_7798));
 AOI22xp5_ASAP7_75t_R g212273__4319 (.A1(n_2216),
    .A2(n_7711),
    .B1(n_3910),
    .B2(n_1819),
    .Y(n_7797));
 AOI221xp5_ASAP7_75t_SL g212274__8428 (.A1(n_3504),
    .A2(n_1810),
    .B1(n_1815),
    .B2(n_2613),
    .C(n_7753),
    .Y(n_7796));
 OAI21xp33_ASAP7_75t_R g212275__5526 (.A1(n_2452),
    .A2(n_7653),
    .B(n_1923),
    .Y(n_7795));
 NAND2xp33_ASAP7_75t_R g212276__6783 (.A(n_2004),
    .B(n_7691),
    .Y(n_7794));
 NOR2xp33_ASAP7_75t_R g212277__3680 (.A(n_3207),
    .B(n_7707),
    .Y(n_7793));
 NAND2xp5_ASAP7_75t_L g212278__1617 (.A(n_2216),
    .B(n_7708),
    .Y(n_7792));
 NAND4xp25_ASAP7_75t_R g212279__2802 (.A(n_2761),
    .B(n_3284),
    .C(n_7621),
    .D(sa10[5]),
    .Y(n_7791));
 A2O1A1Ixp33_ASAP7_75t_SL g212280__1705 (.A1(n_7626),
    .A2(n_6486),
    .B(n_7648),
    .C(sa10[5]),
    .Y(n_7790));
 A2O1A1Ixp33_ASAP7_75t_R g212281__5122 (.A1(n_2379),
    .A2(n_3294),
    .B(n_7661),
    .C(n_2694),
    .Y(n_7789));
 OAI22xp33_ASAP7_75t_SL g212282__8246 (.A1(n_5657),
    .A2(n_7664),
    .B1(n_6095),
    .B2(n_7660),
    .Y(n_7788));
 NAND4xp25_ASAP7_75t_SL g212283__7098 (.A(n_7651),
    .B(n_7643),
    .C(n_7640),
    .D(n_7641),
    .Y(n_7787));
 AOI321xp33_ASAP7_75t_L g212284__6131 (.A1(n_3429),
    .A2(n_3321),
    .A3(n_2092),
    .B1(n_3940),
    .B2(n_2436),
    .C(n_7685),
    .Y(n_7786));
 AOI31xp33_ASAP7_75t_L g212285__1881 (.A1(n_3300),
    .A2(n_1808),
    .A3(n_2286),
    .B(n_7668),
    .Y(n_7785));
 OAI21xp33_ASAP7_75t_R g212286__5115 (.A1(n_1817),
    .A2(n_4271),
    .B(n_7720),
    .Y(n_7784));
 AO21x1_ASAP7_75t_L g212287__7482 (.A1(n_7662),
    .A2(n_5152),
    .B(n_1923),
    .Y(n_7783));
 A2O1A1Ixp33_ASAP7_75t_R g212288__4733 (.A1(n_1802),
    .A2(n_2871),
    .B(n_1804),
    .C(n_5385),
    .Y(n_7782));
 OAI211xp5_ASAP7_75t_SL g212289__6161 (.A1(n_2395),
    .A2(n_4323),
    .B(n_7671),
    .C(n_6210),
    .Y(n_7781));
 AOI21xp33_ASAP7_75t_L g212290__9315 (.A1(n_1808),
    .A2(n_3520),
    .B(n_7704),
    .Y(n_7780));
 NOR2xp33_ASAP7_75t_R g212291__9945 (.A(n_7712),
    .B(n_3601),
    .Y(n_7779));
 A2O1A1Ixp33_ASAP7_75t_R g212292__2883 (.A1(n_1802),
    .A2(n_2517),
    .B(n_1807),
    .C(n_3520),
    .Y(n_7778));
 OAI21xp33_ASAP7_75t_R g212293__2346 (.A1(n_3156),
    .A2(n_1814),
    .B(n_2656),
    .Y(n_7777));
 O2A1O1Ixp33_ASAP7_75t_R g212294__1666 (.A1(n_1801),
    .A2(n_2182),
    .B(n_1806),
    .C(n_1862),
    .Y(n_7776));
 OAI21xp33_ASAP7_75t_R g212295__7410 (.A1(n_1817),
    .A2(n_4036),
    .B(n_1888),
    .Y(n_7775));
 OAI21xp33_ASAP7_75t_R g212296__6417 (.A1(n_3270),
    .A2(n_1814),
    .B(sa20[0]),
    .Y(n_7774));
 OA21x2_ASAP7_75t_L g212297__5477 (.A1(n_7653),
    .A2(n_2989),
    .B(n_3590),
    .Y(n_7773));
 AOI21xp5_ASAP7_75t_R g212298__2398 (.A1(n_3136),
    .A2(n_1808),
    .B(n_7702),
    .Y(n_7772));
 OAI221xp5_ASAP7_75t_L g212299__5107 (.A1(n_7035),
    .A2(n_7627),
    .B1(n_6802),
    .B2(n_7620),
    .C(n_7632),
    .Y(n_7771));
 AO21x1_ASAP7_75t_R g212300__6260 (.A1(n_1813),
    .A2(n_3900),
    .B(n_7718),
    .Y(n_7770));
 OAI21xp33_ASAP7_75t_R g212301__4319 (.A1(n_1806),
    .A2(n_4615),
    .B(n_2284),
    .Y(n_7769));
 A2O1A1Ixp33_ASAP7_75t_R g212302__8428 (.A1(sa20[4]),
    .A2(n_2106),
    .B(n_1805),
    .C(n_2232),
    .Y(n_7768));
 O2A1O1Ixp33_ASAP7_75t_R g212303__5526 (.A1(n_7623),
    .A2(n_2181),
    .B(n_1817),
    .C(n_2348),
    .Y(n_7767));
 AO21x1_ASAP7_75t_R g212304__6783 (.A1(n_1819),
    .A2(n_3900),
    .B(n_7692),
    .Y(n_7766));
 OAI22xp5_ASAP7_75t_SL g212305__3680 (.A1(n_7660),
    .A2(n_6717),
    .B1(n_7666),
    .B2(n_5876),
    .Y(n_7765));
 A2O1A1Ixp33_ASAP7_75t_R g212306__1617 (.A1(n_1801),
    .A2(n_2105),
    .B(n_1815),
    .C(n_4312),
    .Y(n_7764));
 INVxp67_ASAP7_75t_SL g212307 (.A(n_7737),
    .Y(n_7763));
 INVxp67_ASAP7_75t_R g212308 (.A(n_7736),
    .Y(n_7762));
 AOI22xp5_ASAP7_75t_SL g212309__2802 (.A1(n_7657),
    .A2(n_5815),
    .B1(n_1818),
    .B2(n_5230),
    .Y(n_7761));
 AOI31xp33_ASAP7_75t_L g212310__1705 (.A1(n_4329),
    .A2(n_2452),
    .A3(n_1801),
    .B(n_1810),
    .Y(n_7760));
 AOI22xp5_ASAP7_75t_SL g212311__5122 (.A1(n_7665),
    .A2(n_6633),
    .B1(n_7659),
    .B2(n_6103),
    .Y(n_7759));
 A2O1A1Ixp33_ASAP7_75t_R g212312__8246 (.A1(n_2613),
    .A2(n_3300),
    .B(n_7653),
    .C(n_7694),
    .Y(n_7758));
 OAI22xp33_ASAP7_75t_R g212313__7098 (.A1(n_7654),
    .A2(n_4600),
    .B1(n_7623),
    .B2(n_5385),
    .Y(n_7757));
 AOI211xp5_ASAP7_75t_R g212314__6131 (.A1(n_3121),
    .A2(n_2488),
    .B(n_7683),
    .C(n_4610),
    .Y(n_7756));
 OAI21xp33_ASAP7_75t_L g212315__1881 (.A1(n_1812),
    .A2(n_4392),
    .B(n_7716),
    .Y(n_7755));
 OAI21xp5_ASAP7_75t_SL g212316__5115 (.A1(n_7658),
    .A2(n_4388),
    .B(n_7693),
    .Y(n_7754));
 OAI21xp33_ASAP7_75t_L g212317__7482 (.A1(n_1801),
    .A2(n_4390),
    .B(n_7677),
    .Y(n_7753));
 OAI22xp5_ASAP7_75t_L g212318__4733 (.A1(n_1814),
    .A2(n_5308),
    .B1(n_1805),
    .B2(n_3697),
    .Y(n_7752));
 A2O1A1Ixp33_ASAP7_75t_L g212319__6161 (.A1(n_3300),
    .A2(n_4329),
    .B(n_1805),
    .C(n_7700),
    .Y(n_7751));
 AOI22xp5_ASAP7_75t_SL g212320__9315 (.A1(n_7659),
    .A2(n_6788),
    .B1(n_7667),
    .B2(n_6677),
    .Y(n_7750));
 AOI222xp33_ASAP7_75t_SL g212321__9945 (.A1(n_3271),
    .A2(sa20[3]),
    .B1(n_3521),
    .B2(n_1801),
    .C1(n_2344),
    .C2(n_2106),
    .Y(n_7749));
 OAI221xp5_ASAP7_75t_SL g212322__2883 (.A1(n_7004),
    .A2(sa10[2]),
    .B1(n_6467),
    .B2(n_7624),
    .C(n_7644),
    .Y(n_7748));
 AOI22xp33_ASAP7_75t_R g212323__2346 (.A1(n_1802),
    .A2(n_4431),
    .B1(n_1466),
    .B2(n_1807),
    .Y(n_7747));
 OAI221xp5_ASAP7_75t_R g212324__1666 (.A1(n_1806),
    .A2(sa20[4]),
    .B1(n_3694),
    .B2(n_1867),
    .C(n_3462),
    .Y(n_7746));
 O2A1O1Ixp33_ASAP7_75t_R g212325__7410 (.A1(n_1802),
    .A2(n_2217),
    .B(n_7654),
    .C(n_4389),
    .Y(n_7745));
 OAI211xp5_ASAP7_75t_R g212326__6417 (.A1(n_1379),
    .A2(n_4669),
    .B(n_3204),
    .C(n_7665),
    .Y(n_7744));
 OAI321xp33_ASAP7_75t_L g212327__5477 (.A1(n_5992),
    .A2(n_5005),
    .A3(sa10[2]),
    .B1(n_6189),
    .B2(n_7646),
    .C(n_2697),
    .Y(n_7743));
 AOI22xp33_ASAP7_75t_L g212328__2398 (.A1(n_1802),
    .A2(n_4388),
    .B1(sa20[7]),
    .B2(n_1819),
    .Y(n_7742));
 OAI22xp33_ASAP7_75t_R g212329__5107 (.A1(n_7654),
    .A2(n_3453),
    .B1(n_3612),
    .B2(n_1805),
    .Y(n_7741));
 AOI211xp5_ASAP7_75t_R g212330__6260 (.A1(n_1804),
    .A2(n_2181),
    .B(n_3327),
    .C(n_3479),
    .Y(n_7740));
 AO32x1_ASAP7_75t_SL g212331__4319 (.A1(n_1815),
    .A2(n_1606),
    .A3(n_1862),
    .B1(n_1724),
    .B2(n_1807),
    .Y(n_7739));
 AOI22xp33_ASAP7_75t_R g212332__8428 (.A1(n_4391),
    .A2(n_1808),
    .B1(n_1818),
    .B2(n_2013),
    .Y(n_7738));
 OAI22xp5_ASAP7_75t_L g212333__5526 (.A1(n_1806),
    .A2(n_3927),
    .B1(n_1814),
    .B2(n_3136),
    .Y(n_7737));
 OAI22xp33_ASAP7_75t_L g212334__6783 (.A1(n_1806),
    .A2(n_4417),
    .B1(n_3691),
    .B2(n_7658),
    .Y(n_7736));
 OAI22xp33_ASAP7_75t_R g212335__3680 (.A1(n_1801),
    .A2(n_1724),
    .B1(n_2217),
    .B2(n_1806),
    .Y(n_7735));
 OAI22xp33_ASAP7_75t_R g212336__1617 (.A1(n_2871),
    .A2(n_1817),
    .B1(n_1709),
    .B2(n_1814),
    .Y(n_7734));
 AOI22xp33_ASAP7_75t_R g212337__2802 (.A1(n_1810),
    .A2(n_4616),
    .B1(n_1807),
    .B2(n_4036),
    .Y(n_7733));
 OAI22xp33_ASAP7_75t_R g212338__1705 (.A1(n_3348),
    .A2(n_1809),
    .B1(n_2862),
    .B2(n_1806),
    .Y(n_7732));
 AO32x1_ASAP7_75t_L g212339__5122 (.A1(n_4380),
    .A2(n_1808),
    .A3(n_3294),
    .B1(n_4037),
    .B2(n_1815),
    .Y(n_7731));
 AOI22xp33_ASAP7_75t_L g212340__8246 (.A1(n_4400),
    .A2(n_1804),
    .B1(n_1810),
    .B2(n_2500),
    .Y(n_7730));
 OAI22xp33_ASAP7_75t_R g212341__7098 (.A1(n_1809),
    .A2(n_4038),
    .B1(n_2518),
    .B2(n_1806),
    .Y(n_7729));
 INVxp33_ASAP7_75t_R g212342 (.A(n_7727),
    .Y(n_7728));
 INVxp33_ASAP7_75t_R g212343 (.A(n_7725),
    .Y(n_7726));
 INVxp67_ASAP7_75t_R g212345 (.A(n_7709),
    .Y(n_7710));
 INVxp67_ASAP7_75t_R g212346 (.A(n_7708),
    .Y(n_7707));
 INVx1_ASAP7_75t_SL g212347 (.A(n_7705),
    .Y(n_7706));
 NAND3xp33_ASAP7_75t_L g212348__6131 (.A(n_6978),
    .B(n_7630),
    .C(n_1528),
    .Y(n_7701));
 NAND2xp33_ASAP7_75t_R g212349__1881 (.A(n_1819),
    .B(n_4139),
    .Y(n_7700));
 NAND2xp33_ASAP7_75t_R g212350__5115 (.A(n_1815),
    .B(n_3911),
    .Y(n_7699));
 AND2x2_ASAP7_75t_R g212351__7482 (.A(n_1818),
    .B(n_1792),
    .Y(n_7698));
 NAND3xp33_ASAP7_75t_SL g212352__4733 (.A(n_6978),
    .B(n_6872),
    .C(n_7630),
    .Y(n_7697));
 NAND2xp33_ASAP7_75t_R g212353__6161 (.A(n_1810),
    .B(n_3697),
    .Y(n_7727));
 NAND2xp33_ASAP7_75t_R g212354__9315 (.A(n_1815),
    .B(n_4636),
    .Y(n_7725));
 AND2x2_ASAP7_75t_L g212355__9945 (.A(n_7657),
    .B(n_5411),
    .Y(n_7724));
 NAND2xp33_ASAP7_75t_R g212356__2883 (.A(n_1815),
    .B(n_2518),
    .Y(n_7723));
 NAND2xp33_ASAP7_75t_R g212357__2346 (.A(n_1819),
    .B(n_3453),
    .Y(n_7722));
 OR2x2_ASAP7_75t_R g212358__1666 (.A(n_1806),
    .B(n_4392),
    .Y(n_7721));
 NAND2xp5_ASAP7_75t_L g212359__7410 (.A(n_1813),
    .B(n_3600),
    .Y(n_7720));
 NOR2xp33_ASAP7_75t_R g212360__6417 (.A(n_1806),
    .B(n_3463),
    .Y(n_7696));
 NAND2xp5_ASAP7_75t_R g212361__5477 (.A(n_1819),
    .B(n_3632),
    .Y(n_7719));
 NOR2xp33_ASAP7_75t_R g212362__2398 (.A(n_2348),
    .B(n_1812),
    .Y(n_7718));
 NAND2xp5_ASAP7_75t_R g212363__5107 (.A(n_1810),
    .B(n_5381),
    .Y(n_7717));
 NAND2xp5_ASAP7_75t_L g212364__6260 (.A(n_1807),
    .B(n_4339),
    .Y(n_7716));
 NOR2xp33_ASAP7_75t_R g212365__223004 (.A(n_1815),
    .B(n_2182),
    .Y(n_11524));
 NOR2xp33_ASAP7_75t_R g212366__8428 (.A(n_1812),
    .B(n_4636),
    .Y(n_7713));
 NAND2xp5_ASAP7_75t_R g212367__5526 (.A(sa20[0]),
    .B(n_1808),
    .Y(n_7712));
 NOR2xp33_ASAP7_75t_L g212368__6783 (.A(n_7653),
    .B(n_3271),
    .Y(n_7711));
 NAND2xp5_ASAP7_75t_R g212369__3680 (.A(n_1808),
    .B(n_2578),
    .Y(n_7709));
 NOR2xp33_ASAP7_75t_SL g212370__1617 (.A(n_2453),
    .B(n_7658),
    .Y(n_7708));
 NOR2x1_ASAP7_75t_L g212371__2802 (.A(n_1806),
    .B(n_5516),
    .Y(n_7705));
 NOR2xp67_ASAP7_75t_R g212372__1705 (.A(n_1466),
    .B(n_1814),
    .Y(n_7704));
 NOR2xp33_ASAP7_75t_R g212373__5122 (.A(n_1888),
    .B(n_7654),
    .Y(n_7703));
 NOR2x1_ASAP7_75t_L g212374__8246 (.A(n_7658),
    .B(n_2988),
    .Y(n_7702));
 A2O1A1Ixp33_ASAP7_75t_L g212375__7098 (.A1(n_1550),
    .A2(n_5121),
    .B(n_6443),
    .C(n_7663),
    .Y(n_7690));
 AOI22xp33_ASAP7_75t_SL g212376__6131 (.A1(n_7625),
    .A2(n_6659),
    .B1(n_7626),
    .B2(n_6339),
    .Y(n_7689));
 O2A1O1Ixp33_ASAP7_75t_L g212377__1881 (.A1(n_1972),
    .A2(n_4029),
    .B(n_5347),
    .C(n_7664),
    .Y(n_7688));
 A2O1A1Ixp33_ASAP7_75t_R g212378__5115 (.A1(n_1935),
    .A2(n_4578),
    .B(n_5255),
    .C(n_7665),
    .Y(n_7687));
 NAND3xp33_ASAP7_75t_R g212379__7482 (.A(n_4137),
    .B(n_7629),
    .C(n_1528),
    .Y(n_7686));
 OAI221xp5_ASAP7_75t_SL g212380__4733 (.A1(n_3685),
    .A2(n_8178),
    .B1(n_2395),
    .B2(sa10[4]),
    .C(n_7667),
    .Y(n_7685));
 OAI21xp33_ASAP7_75t_R g212381__6161 (.A1(sa20[7]),
    .A2(n_2612),
    .B(n_1807),
    .Y(n_7684));
 OAI21xp33_ASAP7_75t_L g212382__9315 (.A1(n_2430),
    .A2(n_2971),
    .B(n_7665),
    .Y(n_7683));
 AOI211xp5_ASAP7_75t_L g212383__9945 (.A1(n_3587),
    .A2(n_1449),
    .B(n_3943),
    .C(n_7620),
    .Y(n_7682));
 AOI21xp33_ASAP7_75t_R g212384__2883 (.A1(n_3532),
    .A2(n_4312),
    .B(n_7658),
    .Y(n_7681));
 A2O1A1Ixp33_ASAP7_75t_R g212386__2346 (.A1(n_2092),
    .A2(n_5260),
    .B(n_5800),
    .C(n_7659),
    .Y(n_7680));
 OAI21xp33_ASAP7_75t_R g212387__1666 (.A1(n_1607),
    .A2(n_2499),
    .B(n_1819),
    .Y(n_7679));
 AOI21xp33_ASAP7_75t_R g212388__7410 (.A1(n_3294),
    .A2(n_2613),
    .B(n_7654),
    .Y(n_7678));
 OAI21xp33_ASAP7_75t_R g212389__6417 (.A1(n_2453),
    .A2(n_2612),
    .B(n_1804),
    .Y(n_7677));
 OAI221xp5_ASAP7_75t_R g212390__5477 (.A1(n_1665),
    .A2(n_3593),
    .B1(n_2041),
    .B2(n_3102),
    .C(n_7635),
    .Y(n_7676));
 OAI211xp5_ASAP7_75t_R g212391__2398 (.A1(n_2395),
    .A2(n_3617),
    .B(n_7619),
    .C(sa10[5]),
    .Y(n_7675));
 OAI211xp5_ASAP7_75t_R g212392__5107 (.A1(n_2395),
    .A2(n_3664),
    .B(n_7629),
    .C(n_1527),
    .Y(n_7674));
 OAI221xp5_ASAP7_75t_L g212393__6260 (.A1(n_5632),
    .A2(n_1527),
    .B1(n_2395),
    .B2(n_2436),
    .C(n_7629),
    .Y(n_7673));
 AOI221xp5_ASAP7_75t_R g212394__4319 (.A1(n_1549),
    .A2(sa10[4]),
    .B1(n_3273),
    .B2(n_2092),
    .C(n_7620),
    .Y(n_7672));
 AOI211xp5_ASAP7_75t_SL g212395__8428 (.A1(n_4316),
    .A2(n_2092),
    .B(n_5457),
    .C(n_7627),
    .Y(n_7671));
 AOI211xp5_ASAP7_75t_R g212396__5526 (.A1(n_4577),
    .A2(n_1664),
    .B(n_7627),
    .C(sa10[5]),
    .Y(n_7670));
 AOI21xp33_ASAP7_75t_R g212397__6783 (.A1(n_2500),
    .A2(n_4312),
    .B(n_7654),
    .Y(n_7695));
 NAND2xp5_ASAP7_75t_R g212398__3680 (.A(n_3294),
    .B(n_1819),
    .Y(n_7694));
 OAI21xp33_ASAP7_75t_R g212399__1617 (.A1(n_2577),
    .A2(n_2517),
    .B(n_1808),
    .Y(n_7693));
 AOI21xp33_ASAP7_75t_R g212400__2802 (.A1(n_2105),
    .A2(n_2578),
    .B(n_1805),
    .Y(n_7692));
 OAI31xp33_ASAP7_75t_L g212401__1705 (.A1(n_5626),
    .A2(n_5136),
    .A3(n_5196),
    .B(n_7667),
    .Y(n_7691));
 INVxp67_ASAP7_75t_R g212402 (.A(n_7668),
    .Y(n_7669));
 INVxp33_ASAP7_75t_R g212403 (.A(n_7667),
    .Y(n_7666));
 INVxp33_ASAP7_75t_R g212404 (.A(n_7664),
    .Y(n_7663));
 INVxp67_ASAP7_75t_L g212405 (.A(n_7662),
    .Y(n_7661));
 INVx1_ASAP7_75t_L g212406 (.A(n_7660),
    .Y(n_7659));
 INVx2_ASAP7_75t_SL g212407 (.A(n_1819),
    .Y(n_7658));
 INVx1_ASAP7_75t_R g212423 (.A(n_1819),
    .Y(n_1817));
 INVx1_ASAP7_75t_L g212426 (.A(n_7658),
    .Y(n_1818));
 INVx3_ASAP7_75t_SL g212431 (.A(n_1815),
    .Y(n_1814));
 INVxp67_ASAP7_75t_R g212433 (.A(n_1814),
    .Y(n_7657));
 INVx1_ASAP7_75t_L g212450 (.A(n_7654),
    .Y(n_1813));
 INVx2_ASAP7_75t_L g212454 (.A(n_1815),
    .Y(n_7654));
 INVx2_ASAP7_75t_L g212459 (.A(n_1810),
    .Y(n_7653));
 INVxp67_ASAP7_75t_SL g212464 (.A(n_1810),
    .Y(n_1812));
 INVx1_ASAP7_75t_L g212473 (.A(n_1808),
    .Y(n_1809));
 INVx2_ASAP7_75t_L g212487 (.A(n_1807),
    .Y(n_1806));
 HB1xp67_ASAP7_75t_SL g212489 (.A(n_1807),
    .Y(n_1804));
 INVx2_ASAP7_75t_L g212493 (.A(n_1807),
    .Y(n_1805));
 AOI31xp33_ASAP7_75t_L g212501__5122 (.A1(n_5746),
    .A2(n_5496),
    .A3(n_1527),
    .B(n_7628),
    .Y(n_7652));
 OAI21xp5_ASAP7_75t_L g212502__8246 (.A1(n_5907),
    .A2(n_5692),
    .B(n_7619),
    .Y(n_7651));
 A2O1A1Ixp33_ASAP7_75t_L g212503__7098 (.A1(n_1663),
    .A2(n_3891),
    .B(n_6036),
    .C(n_7626),
    .Y(n_7650));
 NOR2xp33_ASAP7_75t_R g212504__6131 (.A(n_1802),
    .B(n_2863),
    .Y(n_7649));
 AOI21xp33_ASAP7_75t_L g212505__1881 (.A1(n_4923),
    .A2(n_5715),
    .B(n_7620),
    .Y(n_7648));
 NOR2xp33_ASAP7_75t_R g212506__5115 (.A(n_1801),
    .B(n_5385),
    .Y(n_7647));
 NOR2xp33_ASAP7_75t_SL g212507__7482 (.A(n_1802),
    .B(n_5385),
    .Y(n_7668));
 NOR2xp33_ASAP7_75t_SL g212508__4733 (.A(sa10[5]),
    .B(n_7620),
    .Y(n_7667));
 NOR2xp33_ASAP7_75t_SL g212509__6161 (.A(sa10[5]),
    .B(n_7622),
    .Y(n_7665));
 NAND2xp5_ASAP7_75t_R g212510__9315 (.A(sa10[5]),
    .B(n_7625),
    .Y(n_7664));
 NOR2xp33_ASAP7_75t_SL g212511__9945 (.A(n_1801),
    .B(n_1888),
    .Y(n_7662));
 NAND2xp5_ASAP7_75t_L g212512__2883 (.A(n_2004),
    .B(n_7625),
    .Y(n_7660));
 AND2x2_ASAP7_75t_SL g212513__2346 (.A(sa20[6]),
    .B(n_1867),
    .Y(n_1819));
 AND2x4_ASAP7_75t_SL g212514__1666 (.A(n_1803),
    .B(sa20[3]),
    .Y(n_1815));
 AND2x4_ASAP7_75t_SL g212515__7410 (.A(n_1803),
    .B(n_1867),
    .Y(n_1810));
 AND2x2_ASAP7_75t_SL g212516__6417 (.A(sa20[6]),
    .B(sa20[3]),
    .Y(n_1807));
 OAI211xp5_ASAP7_75t_L g212517__5477 (.A1(n_3713),
    .A2(n_2961),
    .B(n_5544),
    .C(sa10[2]),
    .Y(n_7646));
 OAI21xp5_ASAP7_75t_L g212518__2398 (.A1(sa10[2]),
    .A2(n_6253),
    .B(n_2697),
    .Y(n_7645));
 A2O1A1Ixp33_ASAP7_75t_L g212519__5107 (.A1(n_1921),
    .A2(n_2975),
    .B(n_5608),
    .C(n_7619),
    .Y(n_7644));
 OAI21xp5_ASAP7_75t_L g212520__6260 (.A1(n_5813),
    .A2(n_5532),
    .B(n_7621),
    .Y(n_7643));
 AO21x1_ASAP7_75t_L g212521__4319 (.A1(n_4785),
    .A2(n_6170),
    .B(n_7622),
    .Y(n_7642));
 A2O1A1Ixp33_ASAP7_75t_L g212522__8428 (.A1(n_2110),
    .A2(n_3668),
    .B(n_5624),
    .C(n_7626),
    .Y(n_7641));
 A2O1A1Ixp33_ASAP7_75t_L g212523__5526 (.A1(n_1935),
    .A2(n_3992),
    .B(n_5700),
    .C(n_7625),
    .Y(n_7640));
 AO21x1_ASAP7_75t_L g212524__6783 (.A1(n_6250),
    .A2(n_6170),
    .B(n_7622),
    .Y(n_7639));
 OAI21xp33_ASAP7_75t_R g212525__3680 (.A1(sa20[3]),
    .A2(n_4391),
    .B(n_7623),
    .Y(n_7638));
 A2O1A1Ixp33_ASAP7_75t_SL g212526__1617 (.A1(n_1664),
    .A2(n_3993),
    .B(n_5978),
    .C(n_7625),
    .Y(n_7637));
 A2O1A1Ixp33_ASAP7_75t_R g212527__2802 (.A1(n_1449),
    .A2(n_4316),
    .B(n_5574),
    .C(n_7619),
    .Y(n_7636));
 AOI21xp33_ASAP7_75t_R g212528__1705 (.A1(n_3541),
    .A2(n_1374),
    .B(n_7624),
    .Y(n_7635));
 OAI31xp33_ASAP7_75t_R g212529__5122 (.A1(n_5931),
    .A2(n_5833),
    .A3(sa10[2]),
    .B(n_7616),
    .Y(n_7634));
 A2O1A1Ixp33_ASAP7_75t_SL g212530__8246 (.A1(n_1663),
    .A2(n_4412),
    .B(n_6447),
    .C(n_7619),
    .Y(n_7633));
 OAI31xp33_ASAP7_75t_R g212531__7098 (.A1(n_4711),
    .A2(n_4671),
    .A3(n_4087),
    .B(n_7621),
    .Y(n_7632));
 A2O1A1Ixp33_ASAP7_75t_R g212532__6131 (.A1(n_2100),
    .A2(n_2940),
    .B(n_5811),
    .C(n_7625),
    .Y(n_7631));
 INVxp33_ASAP7_75t_R g212533 (.A(n_7629),
    .Y(n_7628));
 INVxp67_ASAP7_75t_R g212534 (.A(n_7627),
    .Y(n_7626));
 INVxp33_ASAP7_75t_R g212535 (.A(n_7625),
    .Y(n_7624));
 INVxp67_ASAP7_75t_L g212539 (.A(n_1802),
    .Y(n_7623));
 INVx2_ASAP7_75t_SL g212546 (.A(n_1801),
    .Y(n_1802));
 BUFx2_ASAP7_75t_L g212551 (.A(n_1803),
    .Y(n_1801));
 INVx1_ASAP7_75t_SL g212552 (.A(sa20[6]),
    .Y(n_1803));
 NOR2xp33_ASAP7_75t_R g212553__1881 (.A(sa10[2]),
    .B(n_2004),
    .Y(n_7630));
 NOR2xp33_ASAP7_75t_R g212554__5115 (.A(sa10[2]),
    .B(sa10[5]),
    .Y(n_7629));
 NAND2xp5_ASAP7_75t_L g212555__7482 (.A(n_7615),
    .B(n_1527),
    .Y(n_7627));
 AND2x2_ASAP7_75t_SL g212556__4733 (.A(sa10[2]),
    .B(n_1528),
    .Y(n_7625));
 INVxp67_ASAP7_75t_R g212558 (.A(n_7622),
    .Y(n_7621));
 INVx1_ASAP7_75t_R g212559 (.A(n_7620),
    .Y(n_7619));
 A2O1A1Ixp33_ASAP7_75t_R g212560__6161 (.A1(n_1552),
    .A2(n_5384),
    .B(n_5342),
    .C(sa10[2]),
    .Y(n_7618));
 O2A1O1Ixp33_ASAP7_75t_SL g212561__9315 (.A1(n_2430),
    .A2(n_5401),
    .B(n_5581),
    .C(n_7615),
    .Y(n_7617));
 A2O1A1Ixp33_ASAP7_75t_R g212562__9945 (.A1(n_2728),
    .A2(n_2525),
    .B(n_8180),
    .C(sa10[2]),
    .Y(n_7616));
 NAND2xp5_ASAP7_75t_SL g212563__2883 (.A(n_7615),
    .B(n_1528),
    .Y(n_7622));
 OR2x2_ASAP7_75t_SL g212564__2346 (.A(n_7615),
    .B(sa10[0]),
    .Y(n_7620));
 INVx1_ASAP7_75t_L g212565 (.A(sa10[2]),
    .Y(n_7615));
 XNOR2xp5_ASAP7_75t_SL g212567__1666 (.A(n_7612),
    .B(n_8218),
    .Y(n_7614));
 XOR2xp5_ASAP7_75t_SL g212568__7410 (.A(n_7611),
    .B(n_7608),
    .Y(n_7613));
 XOR2xp5_ASAP7_75t_SL g212569__6417 (.A(n_7609),
    .B(n_8279),
    .Y(n_7612));
 XNOR2xp5_ASAP7_75t_L g212581__5477 (.A(n_7605),
    .B(n_8313),
    .Y(n_7611));
 OAI22xp5_ASAP7_75t_L g212582__2398 (.A1(n_158),
    .A2(n_7606),
    .B1(n_8270),
    .B2(n_7607),
    .Y(n_7610));
 XNOR2xp5_ASAP7_75t_SL g212606__5107 (.A(n_7592),
    .B(n_8260),
    .Y(n_7609));
 XNOR2xp5_ASAP7_75t_SL g212607__6260 (.A(n_7593),
    .B(n_8336),
    .Y(n_7608));
 OAI22xp5_ASAP7_75t_SL g212608__4319 (.A1(n_8267),
    .A2(n_364),
    .B1(n_228),
    .B2(n_8271),
    .Y(n_8218));
 INVxp67_ASAP7_75t_R g212641 (.A(n_7606),
    .Y(n_7607));
 OAI22xp5_ASAP7_75t_L g212673__8428 (.A1(n_8801),
    .A2(n_8258),
    .B1(w3[14]),
    .B2(n_242),
    .Y(n_7606));
 XOR2xp5_ASAP7_75t_R g212674__5526 (.A(n_203),
    .B(w0[18]),
    .Y(n_7605));
 INVxp33_ASAP7_75t_R g212678 (.A(n_1800),
    .Y(n_7602));
 HB1xp67_ASAP7_75t_R g212680 (.A(n_8282),
    .Y(n_1800));
 AO21x1_ASAP7_75t_SL g212688__6783 (.A1(n_8213),
    .A2(n_7528),
    .B(n_7482),
    .Y(n_8281));
 OAI21x1_ASAP7_75t_SL g212689__3680 (.A1(n_7522),
    .A2(n_2033),
    .B(n_7433),
    .Y(n_8280));
 AO21x2_ASAP7_75t_SL g212690__1617 (.A1(n_8203),
    .A2(n_7529),
    .B(n_7439),
    .Y(n_8282));
 INVx2_ASAP7_75t_SL g212694 (.A(n_8273),
    .Y(n_351));
 INVx2_ASAP7_75t_SL g212699 (.A(n_8271),
    .Y(n_364));
 OAI22xp5_ASAP7_75t_L g212700__2802 (.A1(n_235),
    .A2(n_62),
    .B1(n_8300),
    .B2(n_324),
    .Y(n_7593));
 OAI22xp5_ASAP7_75t_SL g212701__1705 (.A1(n_2035),
    .A2(n_8252),
    .B1(w0[14]),
    .B2(n_361),
    .Y(n_7592));
 AO221x2_ASAP7_75t_SL g212702__5122 (.A1(n_1912),
    .A2(n_7446),
    .B1(n_8190),
    .B2(n_7461),
    .C(n_6932),
    .Y(n_8272));
 AO21x2_ASAP7_75t_SL g212703__8246 (.A1(sa22[5]),
    .A2(n_7479),
    .B(n_7460),
    .Y(n_8323));
 OAI21x1_ASAP7_75t_SL g212704__7098 (.A1(n_7480),
    .A2(n_1873),
    .B(n_7435),
    .Y(n_8345));
 AO221x2_ASAP7_75t_SL g212705__6131 (.A1(n_1878),
    .A2(n_7427),
    .B1(n_7471),
    .B2(n_8207),
    .C(n_6933),
    .Y(n_8273));
 AO211x2_ASAP7_75t_SL g212706__1881 (.A1(n_1913),
    .A2(n_7467),
    .B(n_6938),
    .C(n_7525),
    .Y(n_8269));
 AO21x2_ASAP7_75t_SL g212707__5115 (.A1(n_8209),
    .A2(n_8992),
    .B(n_7523),
    .Y(n_8312));
 AO211x2_ASAP7_75t_SL g212708__7482 (.A1(n_2022),
    .A2(n_7481),
    .B(n_6943),
    .C(n_7524),
    .Y(n_8270));
 AO21x2_ASAP7_75t_SL g212709__4733 (.A1(n_8182),
    .A2(n_7526),
    .B(n_7436),
    .Y(n_8271));
 INVxp33_ASAP7_75t_R g212712 (.A(n_7588),
    .Y(n_7589));
 HB1xp67_ASAP7_75t_R g212713 (.A(n_8240),
    .Y(n_7588));
 INVxp33_ASAP7_75t_R g212717 (.A(n_7584),
    .Y(n_7585));
 HB1xp67_ASAP7_75t_R g212718 (.A(n_8264),
    .Y(n_7584));
 OAI21x1_ASAP7_75t_SL g212722__6161 (.A1(n_7438),
    .A2(n_8202),
    .B(n_7380),
    .Y(n_8299));
 AO221x2_ASAP7_75t_SL g212723__9315 (.A1(n_7263),
    .A2(n_2705),
    .B1(n_7374),
    .B2(sa33[5]),
    .C(n_7062),
    .Y(n_8259));
 OAI21x1_ASAP7_75t_SL g212724__9945 (.A1(n_7218),
    .A2(n_1913),
    .B(n_7527),
    .Y(n_8240));
 AO21x2_ASAP7_75t_SL g212725__2883 (.A1(sa21[5]),
    .A2(n_7455),
    .B(n_7432),
    .Y(n_8278));
 AO21x2_ASAP7_75t_SL g212726__2346 (.A1(sa22[5]),
    .A2(n_7442),
    .B(n_7477),
    .Y(n_8275));
 AO221x2_ASAP7_75t_SL g212727__1666 (.A1(n_7411),
    .A2(n_8197),
    .B1(n_7383),
    .B2(n_2022),
    .C(n_6474),
    .Y(n_8310));
 AO221x2_ASAP7_75t_SL g212728__7410 (.A1(n_7376),
    .A2(n_1878),
    .B1(n_7396),
    .B2(n_7353),
    .C(n_6708),
    .Y(n_8318));
 NAND4xp75_ASAP7_75t_SL g212729__6417 (.A(n_7453),
    .B(n_7325),
    .C(n_7097),
    .D(n_6652),
    .Y(n_8264));
 AO21x2_ASAP7_75t_SL g212730__5477 (.A1(sa33[5]),
    .A2(n_7430),
    .B(n_7322),
    .Y(n_8335));
 AO211x2_ASAP7_75t_SL g212731__2398 (.A1(sa21[5]),
    .A2(n_7365),
    .B(n_7086),
    .C(n_7444),
    .Y(n_8258));
 AO221x2_ASAP7_75t_SL g212732__5107 (.A1(n_7316),
    .A2(n_2003),
    .B1(n_7364),
    .B2(sa33[5]),
    .C(n_6799),
    .Y(n_8336));
 INVxp33_ASAP7_75t_R g212740 (.A(n_7573),
    .Y(n_7574));
 HB1xp67_ASAP7_75t_R g212741 (.A(n_8246),
    .Y(n_7573));
 AO21x2_ASAP7_75t_SL g212747__6260 (.A1(n_1540),
    .A2(n_7434),
    .B(n_7321),
    .Y(n_8295));
 AO211x2_ASAP7_75t_SL g212748__4319 (.A1(n_1865),
    .A2(n_7359),
    .B(n_7300),
    .C(n_7413),
    .Y(n_8244));
 AO211x2_ASAP7_75t_SL g212749__8428 (.A1(sa01[5]),
    .A2(n_7331),
    .B(n_7255),
    .C(n_7268),
    .Y(n_8238));
 AO221x2_ASAP7_75t_SL g212750__5526 (.A1(n_7354),
    .A2(n_7192),
    .B1(n_7375),
    .B2(sa02[5]),
    .C(n_6711),
    .Y(n_169));
 AO21x2_ASAP7_75t_SL g212751__6783 (.A1(n_1865),
    .A2(n_7441),
    .B(n_7420),
    .Y(n_8311));
 AO21x2_ASAP7_75t_SL g212752__3680 (.A1(sa21[5]),
    .A2(n_7454),
    .B(n_7326),
    .Y(n_8332));
 NAND4xp75_ASAP7_75t_SL g212753__1617 (.A(n_7469),
    .B(n_7337),
    .C(n_7093),
    .D(n_6411),
    .Y(n_8246));
 AO21x2_ASAP7_75t_SL g212754__2802 (.A1(sa01[5]),
    .A2(n_7428),
    .B(n_7459),
    .Y(n_8268));
 AO211x2_ASAP7_75t_SL g212755__1705 (.A1(n_1865),
    .A2(n_7332),
    .B(n_6999),
    .C(n_7224),
    .Y(n_8243));
 AO221x2_ASAP7_75t_SL g212756__5122 (.A1(n_7370),
    .A2(sa22[5]),
    .B1(n_7330),
    .B2(n_1879),
    .C(n_6700),
    .Y(n_8325));
 AO21x2_ASAP7_75t_SL g212757__8246 (.A1(sa33[5]),
    .A2(n_7431),
    .B(n_7462),
    .Y(n_8279));
 AO221x2_ASAP7_75t_SL g212758__7098 (.A1(n_7392),
    .A2(n_7470),
    .B1(n_7249),
    .B2(sa00[5]),
    .C(n_7005),
    .Y(n_8267));
 INVxp33_ASAP7_75t_R g212761 (.A(n_7564),
    .Y(n_7565));
 HB1xp67_ASAP7_75t_R g212762 (.A(n_8291),
    .Y(n_7564));
 INVxp33_ASAP7_75t_R g212768 (.A(n_8225),
    .Y(n_7560));
 INVxp33_ASAP7_75t_R g212773 (.A(n_8309),
    .Y(n_7556));
 INVxp33_ASAP7_75t_R g212774 (.A(n_7554),
    .Y(n_7555));
 HB1xp67_ASAP7_75t_R g212775 (.A(n_8227),
    .Y(n_7554));
 INVxp33_ASAP7_75t_R g212780 (.A(n_8232),
    .Y(n_7550));
 INVxp33_ASAP7_75t_R g212781 (.A(n_7548),
    .Y(n_7549));
 HB1xp67_ASAP7_75t_R g212782 (.A(n_8248),
    .Y(n_7548));
 INVxp33_ASAP7_75t_R g212783 (.A(n_7546),
    .Y(n_7547));
 HB1xp67_ASAP7_75t_R g212784 (.A(n_8235),
    .Y(n_7546));
 INVxp33_ASAP7_75t_R g212788 (.A(n_7541),
    .Y(n_7542));
 HB1xp67_ASAP7_75t_R g212789 (.A(n_178),
    .Y(n_7541));
 INVxp33_ASAP7_75t_R g212790 (.A(n_7539),
    .Y(n_7540));
 HB1xp67_ASAP7_75t_R g212791 (.A(n_8230),
    .Y(n_7539));
 INVx2_ASAP7_75t_SL g212792 (.A(n_7537),
    .Y(n_332));
 INVxp33_ASAP7_75t_R g212797 (.A(n_8339),
    .Y(n_7533));
 OAI21xp5_ASAP7_75t_SL g212801__6131 (.A1(n_1873),
    .A2(n_7314),
    .B(n_7394),
    .Y(n_7529));
 OAI21xp5_ASAP7_75t_SL g212802__1881 (.A1(n_1895),
    .A2(n_7320),
    .B(n_7398),
    .Y(n_7528));
 AOI321xp33_ASAP7_75t_SL g212803__5115 (.A1(n_7132),
    .A2(n_6537),
    .A3(n_5259),
    .B1(n_6743),
    .B2(n_3439),
    .C(n_6375),
    .Y(n_7527));
 OAI22xp5_ASAP7_75t_SL g212804__7482 (.A1(n_8209),
    .A2(n_7318),
    .B1(n_1865),
    .B2(n_7234),
    .Y(n_7526));
 AOI21xp5_ASAP7_75t_SL g212805__4733 (.A1(n_7397),
    .A2(n_7296),
    .B(n_1913),
    .Y(n_7525));
 O2A1O1Ixp33_ASAP7_75t_SL g212806__6161 (.A1(n_1510),
    .A2(n_7231),
    .B(n_6919),
    .C(n_2022),
    .Y(n_7524));
 A2O1A1Ixp33_ASAP7_75t_SL g212807__9315 (.A1(n_7074),
    .A2(n_7273),
    .B(n_8209),
    .C(n_6720),
    .Y(n_7523));
 AOI221xp5_ASAP7_75t_SL g212808__9945 (.A1(n_6695),
    .A2(n_2189),
    .B1(n_7000),
    .B2(n_2673),
    .C(n_7333),
    .Y(n_7522));
 NAND2x1_ASAP7_75t_SL g212809__2883 (.A(n_7336),
    .B(n_7458),
    .Y(n_8346));
 NAND4xp75_ASAP7_75t_SL g212810__2346 (.A(n_7217),
    .B(n_7267),
    .C(n_7269),
    .D(n_6617),
    .Y(n_8285));
 NAND3x1_ASAP7_75t_SL g212811__1666 (.A(n_7391),
    .B(n_7216),
    .C(n_7254),
    .Y(n_8291));
 NAND2x1_ASAP7_75t_SL g212812__7410 (.A(n_7466),
    .B(n_7323),
    .Y(n_8303));
 AO211x2_ASAP7_75t_SL g212813__6417 (.A1(n_2022),
    .A2(n_7301),
    .B(n_7106),
    .C(n_7406),
    .Y(n_8242));
 NAND3x2_ASAP7_75t_SL g212814__5477 (.B(n_7219),
    .C(n_7285),
    .Y(n_8296),
    .A(n_7386));
 AO221x2_ASAP7_75t_SL g212815__2398 (.A1(n_7334),
    .A2(n_8207),
    .B1(n_7236),
    .B2(n_1878),
    .C(n_7282),
    .Y(n_8225));
 AO21x2_ASAP7_75t_SL g212816__5107 (.A1(sa30[5]),
    .A2(n_7351),
    .B(n_7361),
    .Y(n_8262));
 AO21x2_ASAP7_75t_SL g212817__6260 (.A1(sa30[5]),
    .A2(n_7324),
    .B(n_7408),
    .Y(n_8338));
 AO211x2_ASAP7_75t_SL g212818__4319 (.A1(sa01[5]),
    .A2(n_7309),
    .B(n_7089),
    .C(n_7221),
    .Y(n_131));
 AO21x2_ASAP7_75t_SL g212819__8428 (.A1(n_2022),
    .A2(n_7350),
    .B(n_7313),
    .Y(n_8309));
 NAND4xp75_ASAP7_75t_SL g212820__5526 (.A(n_7080),
    .B(n_7274),
    .C(n_7373),
    .D(n_7229),
    .Y(n_8227));
 OAI21x1_ASAP7_75t_SL g212821__6783 (.A1(n_7329),
    .A2(sa02[5]),
    .B(n_7429),
    .Y(n_8305));
 OAI21x1_ASAP7_75t_SL g212822__3680 (.A1(n_7307),
    .A2(sa02[5]),
    .B(n_7348),
    .Y(n_8221));
 AO21x2_ASAP7_75t_SL g212823__1617 (.A1(sa00[5]),
    .A2(n_7379),
    .B(n_7412),
    .Y(n_8301));
 AO211x2_ASAP7_75t_SL g212824__2802 (.A1(n_2033),
    .A2(n_7308),
    .B(n_7237),
    .C(n_7261),
    .Y(n_8232));
 OAI21x1_ASAP7_75t_SL g212825__1705 (.A1(n_8207),
    .A2(n_7220),
    .B(n_7440),
    .Y(n_8248));
 NAND3x2_ASAP7_75t_SL g212826__5122 (.B(n_7404),
    .C(n_7407),
    .Y(n_8235),
    .A(n_7437));
 OAI21x1_ASAP7_75t_SL g212827__8246 (.A1(n_7369),
    .A2(sa32[5]),
    .B(n_7312),
    .Y(n_8234));
 NAND2x2_ASAP7_75t_SL g212828__7098 (.A(n_7423),
    .B(n_7465),
    .Y(n_8247));
 AO211x2_ASAP7_75t_SL g212829__6131 (.A1(n_1895),
    .A2(n_7385),
    .B(n_7228),
    .C(n_7280),
    .Y(n_178));
 OAI21x1_ASAP7_75t_SL g212830__1881 (.A1(n_7416),
    .A2(sa21[5]),
    .B(n_7382),
    .Y(n_8230));
 OAI21x1_ASAP7_75t_SL g212831__5115 (.A1(n_7343),
    .A2(n_1879),
    .B(n_7403),
    .Y(n_7537));
 OAI21x1_ASAP7_75t_SL g212832__7482 (.A1(n_7244),
    .A2(n_8202),
    .B(n_7457),
    .Y(n_8236));
 OAI21x1_ASAP7_75t_SL g212833__4733 (.A1(n_8183),
    .A2(n_7338),
    .B(n_7352),
    .Y(n_8333));
 OAI21x1_ASAP7_75t_SL g212834__6161 (.A1(n_7426),
    .A2(n_1878),
    .B(n_7367),
    .Y(n_8317));
 AO21x2_ASAP7_75t_SL g212835__9315 (.A1(sa30[5]),
    .A2(n_7345),
    .B(n_7390),
    .Y(n_8339));
 OAI21x1_ASAP7_75t_SL g212836__9945 (.A1(n_8190),
    .A2(n_7372),
    .B(n_7357),
    .Y(n_8315));
 AO211x2_ASAP7_75t_SL g212837__2883 (.A1(sa32[5]),
    .A2(n_7328),
    .B(n_7084),
    .C(n_7417),
    .Y(n_8266));
 AO221x1_ASAP7_75t_SL g212838__2346 (.A1(n_7340),
    .A2(sa00[5]),
    .B1(n_7190),
    .B2(n_2692),
    .C(n_7272),
    .Y(n_8300));
 INVxp33_ASAP7_75t_R g212841 (.A(n_7518),
    .Y(n_7519));
 HB1xp67_ASAP7_75t_R g212842 (.A(n_8298),
    .Y(n_7518));
 INVxp33_ASAP7_75t_R g212847 (.A(n_7513),
    .Y(n_7514));
 HB1xp67_ASAP7_75t_R g212848 (.A(n_8294),
    .Y(n_7513));
 INVxp33_ASAP7_75t_R g212855 (.A(n_8340),
    .Y(n_7507));
 INVxp33_ASAP7_75t_R g212860 (.A(n_7502),
    .Y(n_7503));
 HB1xp67_ASAP7_75t_R g212861 (.A(n_8219),
    .Y(n_7502));
 INVxp33_ASAP7_75t_R g212869 (.A(n_7494),
    .Y(n_7495));
 HB1xp67_ASAP7_75t_R g212870 (.A(n_69),
    .Y(n_7494));
 INVxp33_ASAP7_75t_R g212872 (.A(n_7491),
    .Y(n_7492));
 HB1xp67_ASAP7_75t_R g212873 (.A(n_8241),
    .Y(n_7491));
 INVx1_ASAP7_75t_L g212884 (.A(n_62),
    .Y(n_324));
 HB1xp67_ASAP7_75t_SL g212885 (.A(n_8324),
    .Y(n_62));
 A2O1A1Ixp33_ASAP7_75t_SL g212886__1666 (.A1(n_6849),
    .A2(n_7266),
    .B(n_1895),
    .C(n_7003),
    .Y(n_7482));
 OAI21xp5_ASAP7_75t_SL g212887__7410 (.A1(n_1510),
    .A2(n_7319),
    .B(n_7227),
    .Y(n_7481));
 AOI221xp5_ASAP7_75t_SL g212888__6417 (.A1(n_6601),
    .A2(n_2608),
    .B1(n_7209),
    .B2(n_1981),
    .C(n_6945),
    .Y(n_7480));
 OAI211xp5_ASAP7_75t_SL g212889__5477 (.A1(sa22[2]),
    .A2(n_7206),
    .B(n_6774),
    .C(n_6661),
    .Y(n_7479));
 OAI221xp5_ASAP7_75t_SL g212891__5107 (.A1(n_6491),
    .A2(n_3359),
    .B1(n_7233),
    .B2(n_2695),
    .C(n_6857),
    .Y(n_7477));
 AO221x2_ASAP7_75t_SL g212892__6260 (.A1(n_7356),
    .A2(n_8190),
    .B1(n_1912),
    .B2(n_7235),
    .C(n_6354),
    .Y(n_8245));
 AO21x2_ASAP7_75t_SL g212893__4319 (.A1(n_1878),
    .A2(n_7362),
    .B(n_7293),
    .Y(n_8319));
 OAI21x1_ASAP7_75t_SL g212894__8428 (.A1(n_7414),
    .A2(sa32[2]),
    .B(n_7395),
    .Y(n_8298));
 OAI21x1_ASAP7_75t_SL g212895__5526 (.A1(n_7393),
    .A2(n_2003),
    .B(n_7456),
    .Y(n_8337));
 OAI21x1_ASAP7_75t_SL g212896__6783 (.A1(n_8183),
    .A2(n_7371),
    .B(n_7422),
    .Y(n_8334));
 AO211x2_ASAP7_75t_SL g212897__3680 (.A1(n_8197),
    .A2(n_7387),
    .B(n_7368),
    .C(n_7230),
    .Y(n_8222));
 NAND4xp75_ASAP7_75t_SL g212898__1617 (.A(n_7223),
    .B(n_7304),
    .C(n_7245),
    .D(n_7292),
    .Y(n_8294));
 AO211x2_ASAP7_75t_SL g212899__2802 (.A1(sa32[5]),
    .A2(n_7246),
    .B(n_6370),
    .C(n_7306),
    .Y(n_8265));
 OAI21x1_ASAP7_75t_SL g212900__1705 (.A1(n_7415),
    .A2(n_8202),
    .B(n_7358),
    .Y(n_8283));
 AO21x2_ASAP7_75t_SL g212901__5122 (.A1(sa31[5]),
    .A2(n_7388),
    .B(n_7418),
    .Y(n_8343));
 OAI21x1_ASAP7_75t_SL g212902__8246 (.A1(n_2022),
    .A2(n_7341),
    .B(n_7472),
    .Y(n_8308));
 AO21x2_ASAP7_75t_SL g212903__7098 (.A1(sa30[5]),
    .A2(n_7378),
    .B(n_7421),
    .Y(n_8340));
 AO21x2_ASAP7_75t_SL g212904__6131 (.A1(n_1884),
    .A2(n_7311),
    .B(n_7445),
    .Y(n_8220));
 OAI21xp5_ASAP7_75t_SL g212905__1881 (.A1(n_7188),
    .A2(n_7025),
    .B(n_7463),
    .Y(n_8286));
 AO21x2_ASAP7_75t_SL g212906__5115 (.A1(sa31[5]),
    .A2(n_7344),
    .B(n_7381),
    .Y(n_8342));
 OAI21x1_ASAP7_75t_SL g212907__7482 (.A1(n_7355),
    .A2(sa00[5]),
    .B(n_7305),
    .Y(n_8219));
 AO211x2_ASAP7_75t_SL g212908__4733 (.A1(n_1895),
    .A2(n_7299),
    .B(n_6896),
    .C(n_7399),
    .Y(n_129));
 AO21x2_ASAP7_75t_SL g212909__6161 (.A1(sa01[5]),
    .A2(n_7317),
    .B(n_7464),
    .Y(n_8302));
 OAI21x1_ASAP7_75t_SL g212910__9315 (.A1(sa02[5]),
    .A2(n_7400),
    .B(n_7443),
    .Y(n_8239));
 OAI21x1_ASAP7_75t_SL g212911__9945 (.A1(n_7349),
    .A2(n_8190),
    .B(n_7405),
    .Y(n_8316));
 AO221x2_ASAP7_75t_SL g212912__2883 (.A1(n_7215),
    .A2(n_1895),
    .B1(n_7270),
    .B2(sa31[5]),
    .C(n_6827),
    .Y(n_8263));
 NAND4xp75_ASAP7_75t_SL g212913__2346 (.A(n_7419),
    .B(n_7222),
    .C(n_7271),
    .D(n_7070),
    .Y(n_69));
 AO21x2_ASAP7_75t_SL g212914__1666 (.A1(n_8190),
    .A2(n_7360),
    .B(n_7335),
    .Y(n_8314));
 AO221x2_ASAP7_75t_SL g212915__7410 (.A1(n_7377),
    .A2(n_8197),
    .B1(n_7242),
    .B2(n_2022),
    .C(n_6664),
    .Y(n_8241));
 OAI21x1_ASAP7_75t_SL g212916__6417 (.A1(n_7327),
    .A2(sa11[2]),
    .B(n_7363),
    .Y(n_8287));
 OAI21x1_ASAP7_75t_SL g212917__5477 (.A1(n_7384),
    .A2(n_1913),
    .B(n_7425),
    .Y(n_8307));
 AO22x2_ASAP7_75t_SL g212918__2398 (.A1(n_2003),
    .A2(n_7310),
    .B1(sa33[5]),
    .B2(n_7286),
    .Y(n_8231));
 AO221x2_ASAP7_75t_SL g212919__5107 (.A1(n_7339),
    .A2(sa01[5]),
    .B1(n_7248),
    .B2(n_1884),
    .C(n_7143),
    .Y(n_8304));
 AO21x2_ASAP7_75t_SL g212920__6260 (.A1(sa32[5]),
    .A2(n_7366),
    .B(n_7468),
    .Y(n_8344));
 AO21x2_ASAP7_75t_SL g212921__4319 (.A1(n_1865),
    .A2(n_7402),
    .B(n_7424),
    .Y(n_8313));
 AO21x1_ASAP7_75t_SL g212922__8428 (.A1(sa33[5]),
    .A2(n_7315),
    .B(n_7401),
    .Y(n_8260));
 AO21x2_ASAP7_75t_SL g212923__5526 (.A1(sa22[5]),
    .A2(n_7346),
    .B(n_7389),
    .Y(n_8252));
 NAND4xp75_ASAP7_75t_SL g212924__6783 (.A(n_8993),
    .B(n_7208),
    .C(n_7187),
    .D(n_6989),
    .Y(n_8324));
 INVxp33_ASAP7_75t_R g212926 (.A(n_7474),
    .Y(n_7475));
 HB1xp67_ASAP7_75t_R g212927 (.A(n_8284),
    .Y(n_7474));
 O2A1O1Ixp5_ASAP7_75t_SL g212929__3680 (.A1(n_6985),
    .A2(n_6577),
    .B(n_2362),
    .C(n_7145),
    .Y(n_7472));
 A2O1A1Ixp33_ASAP7_75t_SL g212930__1617 (.A1(n_6906),
    .A2(n_7196),
    .B(n_1966),
    .C(n_6591),
    .Y(n_7471));
 AOI31xp33_ASAP7_75t_SL g212931__2802 (.A1(n_7191),
    .A2(n_6908),
    .A3(n_8202),
    .B(sa00[0]),
    .Y(n_7470));
 A2O1A1Ixp33_ASAP7_75t_SL g212932__1705 (.A1(n_2611),
    .A2(n_6248),
    .B(n_7303),
    .C(n_1912),
    .Y(n_7469));
 A2O1A1Ixp33_ASAP7_75t_SL g212933__5122 (.A1(n_7194),
    .A2(n_7095),
    .B(sa32[5]),
    .C(n_6446),
    .Y(n_7468));
 A2O1A1Ixp33_ASAP7_75t_SL g212934__8246 (.A1(n_6909),
    .A2(n_7197),
    .B(sa02[0]),
    .C(n_6573),
    .Y(n_7467));
 OAI21x1_ASAP7_75t_SL g212935__7098 (.A1(n_7078),
    .A2(n_7297),
    .B(sa01[5]),
    .Y(n_7466));
 OAI21x1_ASAP7_75t_SL g212936__6131 (.A1(n_7251),
    .A2(n_6834),
    .B(n_8207),
    .Y(n_7465));
 OAI21xp5_ASAP7_75t_SL g212937__1881 (.A1(n_2701),
    .A2(n_7259),
    .B(n_7136),
    .Y(n_7464));
 AOI311xp33_ASAP7_75t_SL g212938__5115 (.A1(n_6826),
    .A2(n_6526),
    .A3(n_2712),
    .B(n_7050),
    .C(n_7278),
    .Y(n_7463));
 A2O1A1Ixp33_ASAP7_75t_SL g212939__7482 (.A1(n_6907),
    .A2(n_7193),
    .B(n_2706),
    .C(n_7112),
    .Y(n_7462));
 A2O1A1Ixp33_ASAP7_75t_SL g212940__4733 (.A1(n_6905),
    .A2(n_7195),
    .B(sa12[0]),
    .C(n_6502),
    .Y(n_7461));
 OAI21xp5_ASAP7_75t_SL g212941__6161 (.A1(n_2695),
    .A2(n_7260),
    .B(n_7033),
    .Y(n_7460));
 OAI21xp5_ASAP7_75t_SL g212942__9315 (.A1(n_2701),
    .A2(n_7238),
    .B(n_7085),
    .Y(n_7459));
 OAI21xp5_ASAP7_75t_SL g212943__9945 (.A1(n_7121),
    .A2(n_7250),
    .B(sa32[5]),
    .Y(n_7458));
 AOI321xp33_ASAP7_75t_SL g212944__2883 (.A1(n_7101),
    .A2(n_6532),
    .A3(n_6076),
    .B1(n_6738),
    .B2(n_3378),
    .C(n_6367),
    .Y(n_7457));
 AOI31xp67_ASAP7_75t_SL g212945__2346 (.A1(n_7141),
    .A2(n_7053),
    .A3(n_2719),
    .B(n_7043),
    .Y(n_7456));
 NAND3xp33_ASAP7_75t_SL g212946__1666 (.A(n_7239),
    .B(n_7173),
    .C(n_7038),
    .Y(n_7455));
 A2O1A1Ixp33_ASAP7_75t_SL g212947__7410 (.A1(n_6971),
    .A2(n_7014),
    .B(sa21[2]),
    .C(n_7015),
    .Y(n_7454));
 AO21x1_ASAP7_75t_SL g212948__6417 (.A1(n_6715),
    .A2(n_7211),
    .B(n_1895),
    .Y(n_7453));
 OR2x6_ASAP7_75t_SL g212949__5477 (.A(n_7410),
    .B(n_7347),
    .Y(n_8261));
 NAND4xp25_ASAP7_75t_SL g212950__2398 (.A(n_7241),
    .B(n_7291),
    .C(n_7252),
    .D(n_7063),
    .Y(n_8284));
 OR3x2_ASAP7_75t_SL g212951__5107 (.A(n_7298),
    .B(n_7256),
    .C(n_7295),
    .Y(n_37));
 INVxp33_ASAP7_75t_R g212953 (.A(n_7450),
    .Y(n_7451));
 HB1xp67_ASAP7_75t_R g212954 (.A(n_8289),
    .Y(n_7450));
 INVxp33_ASAP7_75t_R g212956 (.A(n_7447),
    .Y(n_7448));
 OAI311xp33_ASAP7_75t_SL g212958__6260 (.A1(n_7031),
    .A2(n_7016),
    .A3(sa12[0]),
    .B1(n_5911),
    .C1(n_7073),
    .Y(n_7446));
 OAI321xp33_ASAP7_75t_SL g212959__4319 (.A1(n_6807),
    .A2(n_2151),
    .A3(n_1884),
    .B1(n_2376),
    .B2(n_7213),
    .C(n_6884),
    .Y(n_7445));
 AO32x1_ASAP7_75t_SL g212960__8428 (.A1(n_7110),
    .A2(n_6878),
    .A3(n_6062),
    .B1(n_6112),
    .B2(n_3466),
    .Y(n_7444));
 O2A1O1Ixp5_ASAP7_75t_SL g212961__5526 (.A1(n_7091),
    .A2(n_7179),
    .B(sa02[5]),
    .C(n_6653),
    .Y(n_7443));
 OAI211xp5_ASAP7_75t_SL g212962__6783 (.A1(n_2672),
    .A2(n_7029),
    .B(n_7232),
    .C(n_7059),
    .Y(n_7442));
 OAI21xp5_ASAP7_75t_SL g212963__3680 (.A1(sa11[2]),
    .A2(n_7210),
    .B(n_7169),
    .Y(n_7441));
 AOI321xp33_ASAP7_75t_SL g212964__1617 (.A1(n_7129),
    .A2(n_6534),
    .A3(n_5360),
    .B1(n_6727),
    .B2(n_3430),
    .C(n_6404),
    .Y(n_7440));
 A2O1A1Ixp33_ASAP7_75t_SL g212965__2802 (.A1(n_6475),
    .A2(n_7055),
    .B(n_1873),
    .C(n_7066),
    .Y(n_7439));
 AOI211xp5_ASAP7_75t_SL g212966__1705 (.A1(n_7203),
    .A2(n_1531),
    .B(n_6898),
    .C(n_6922),
    .Y(n_7438));
 AND4x2_ASAP7_75t_SL g212967__5122 (.A(n_7279),
    .B(n_7287),
    .C(n_7058),
    .D(n_6882),
    .Y(n_7437));
 A2O1A1Ixp33_ASAP7_75t_SL g212968__8246 (.A1(n_6847),
    .A2(n_7077),
    .B(n_8209),
    .C(n_7142),
    .Y(n_7436));
 O2A1O1Ixp5_ASAP7_75t_SL g212969__7098 (.A1(n_6963),
    .A2(n_7013),
    .B(n_2722),
    .C(n_7036),
    .Y(n_7435));
 OAI22xp5_ASAP7_75t_SL g212970__6131 (.A1(n_2003),
    .A2(n_7205),
    .B1(sa33[5]),
    .B2(n_7168),
    .Y(n_7434));
 AOI221x1_ASAP7_75t_SL g212971__1881 (.A1(n_6522),
    .A2(n_3353),
    .B1(n_7024),
    .B2(n_2696),
    .C(n_6864),
    .Y(n_7433));
 OAI221xp5_ASAP7_75t_SL g212972__5115 (.A1(n_6516),
    .A2(n_3336),
    .B1(n_7022),
    .B2(n_2717),
    .C(n_6921),
    .Y(n_7432));
 OAI211xp5_ASAP7_75t_SL g212973__7482 (.A1(n_2663),
    .A2(n_6998),
    .B(n_7240),
    .C(n_7065),
    .Y(n_7431));
 OAI21xp5_ASAP7_75t_SL g212974__4733 (.A1(sa33[2]),
    .A2(n_7258),
    .B(n_7020),
    .Y(n_7430));
 AOI21x1_ASAP7_75t_SL g212975__6161 (.A1(n_7207),
    .A2(n_2369),
    .B(n_7202),
    .Y(n_7429));
 OAI221xp5_ASAP7_75t_SL g212976__9315 (.A1(n_6994),
    .A2(n_2665),
    .B1(n_6691),
    .B2(n_2602),
    .C(n_7262),
    .Y(n_7428));
 OAI211xp5_ASAP7_75t_SL g212977__9945 (.A1(n_2661),
    .A2(n_6993),
    .B(n_7243),
    .C(n_7071),
    .Y(n_7427));
 AO21x2_ASAP7_75t_SL g212978__2883 (.A1(n_8190),
    .A2(n_7276),
    .B(n_7342),
    .Y(n_8224));
 NAND4xp25_ASAP7_75t_SL g212979__2346 (.A(n_7158),
    .B(n_7264),
    .C(n_7265),
    .D(n_7039),
    .Y(n_8289));
 AO22x2_ASAP7_75t_SL g212980__1666 (.A1(n_8209),
    .A2(n_7281),
    .B1(n_1865),
    .B2(n_7283),
    .Y(n_357));
 AO211x2_ASAP7_75t_SL g212981__7410 (.A1(sa21[5]),
    .A2(n_7247),
    .B(n_7019),
    .C(n_7204),
    .Y(n_7447));
 AOI321xp33_ASAP7_75t_SL g212982__6417 (.A1(n_6417),
    .A2(n_6881),
    .A3(n_8188),
    .B1(n_6621),
    .B2(n_2220),
    .C(n_6570),
    .Y(n_7426));
 AOI221x1_ASAP7_75t_SL g212983__5477 (.A1(n_6658),
    .A2(n_3439),
    .B1(n_7103),
    .B2(n_7138),
    .C(n_6376),
    .Y(n_7425));
 OAI211xp5_ASAP7_75t_SL g212984__2398 (.A1(n_7098),
    .A2(n_7155),
    .B(n_6901),
    .C(n_6421),
    .Y(n_7424));
 AND3x1_ASAP7_75t_SL g212985__5107 (.A(n_7075),
    .B(n_7122),
    .C(n_6812),
    .Y(n_7423));
 AOI21xp5_ASAP7_75t_SL g212986__6260 (.A1(n_7072),
    .A2(n_7154),
    .B(n_7289),
    .Y(n_7422));
 OAI21xp5_ASAP7_75t_SL g212987__4319 (.A1(n_7144),
    .A2(n_7102),
    .B(n_7225),
    .Y(n_7421));
 OAI211xp5_ASAP7_75t_SL g212988__8428 (.A1(n_2723),
    .A2(n_7151),
    .B(n_6820),
    .C(n_6843),
    .Y(n_7420));
 A2O1A1Ixp33_ASAP7_75t_SL g212989__5526 (.A1(n_8213),
    .A2(n_6912),
    .B(n_6958),
    .C(n_2700),
    .Y(n_7419));
 OAI21xp5_ASAP7_75t_SL g212990__6783 (.A1(n_6964),
    .A2(n_7099),
    .B(n_7275),
    .Y(n_7418));
 A2O1A1Ixp33_ASAP7_75t_SL g212991__3680 (.A1(n_1980),
    .A2(n_6760),
    .B(n_6929),
    .C(n_6372),
    .Y(n_7417));
 AOI211xp5_ASAP7_75t_SL g212992__1617 (.A1(n_6543),
    .A2(n_6228),
    .B(n_7087),
    .C(n_6674),
    .Y(n_7416));
 AOI21xp5_ASAP7_75t_SL g212993__2802 (.A1(n_7118),
    .A2(n_7189),
    .B(n_6453),
    .Y(n_7415));
 O2A1O1Ixp33_ASAP7_75t_SL g212994__1705 (.A1(n_1980),
    .A2(n_6890),
    .B(n_7083),
    .C(n_7288),
    .Y(n_7414));
 NOR3xp33_ASAP7_75t_SL g212995__5122 (.A(n_7100),
    .B(n_6541),
    .C(n_4859),
    .Y(n_7413));
 OAI21xp5_ASAP7_75t_SL g212996__8246 (.A1(n_2691),
    .A2(n_7199),
    .B(n_7146),
    .Y(n_7412));
 A2O1A1Ixp33_ASAP7_75t_SL g212997__7098 (.A1(n_6433),
    .A2(n_6835),
    .B(n_3229),
    .C(n_6962),
    .Y(n_7411));
 AOI21xp5_ASAP7_75t_SL g212998__6131 (.A1(n_6981),
    .A2(n_7157),
    .B(n_2033),
    .Y(n_7410));
 AO21x1_ASAP7_75t_SL g213000__5115 (.A1(n_2696),
    .A2(n_7001),
    .B(n_7125),
    .Y(n_7408));
 A2O1A1Ixp33_ASAP7_75t_SL g213001__7482 (.A1(n_2678),
    .A2(n_5889),
    .B(n_7149),
    .C(sa00[5]),
    .Y(n_7407));
 OAI31xp33_ASAP7_75t_SL g213002__4733 (.A1(n_6928),
    .A2(n_6546),
    .A3(n_6085),
    .B(n_6348),
    .Y(n_7406));
 AND2x2_ASAP7_75t_SL g213003__6161 (.A(n_7294),
    .B(n_7148),
    .Y(n_7405));
 OA21x2_ASAP7_75t_SL g213004__9315 (.A1(n_8202),
    .A2(n_7140),
    .B(n_6775),
    .Y(n_7404));
 AOI221x1_ASAP7_75t_SL g213005__9945 (.A1(n_6639),
    .A2(n_6176),
    .B1(n_7133),
    .B2(n_6953),
    .C(n_6665),
    .Y(n_7403));
 NAND2xp5_ASAP7_75t_SL g213006__2883 (.A(n_6863),
    .B(n_7277),
    .Y(n_7402));
 OAI221xp5_ASAP7_75t_SL g213007__2346 (.A1(n_7060),
    .A2(n_6975),
    .B1(n_6726),
    .B2(n_3408),
    .C(n_6692),
    .Y(n_7401));
 AOI21xp5_ASAP7_75t_SL g213008__1666 (.A1(n_7088),
    .A2(n_7181),
    .B(n_6854),
    .Y(n_7400));
 A2O1A1Ixp33_ASAP7_75t_SL g213009__7410 (.A1(n_6927),
    .A2(n_6868),
    .B(n_2699),
    .C(n_6892),
    .Y(n_7399));
 A2O1A1Ixp33_ASAP7_75t_SL g213010__6417 (.A1(sa31[2]),
    .A2(n_6768),
    .B(n_6915),
    .C(n_1895),
    .Y(n_7398));
 AOI221xp5_ASAP7_75t_SL g213011__5477 (.A1(n_6937),
    .A2(n_2224),
    .B1(n_6773),
    .B2(n_2596),
    .C(n_6853),
    .Y(n_7397));
 AOI31xp33_ASAP7_75t_SL g213012__2398 (.A1(n_7183),
    .A2(n_6949),
    .A3(n_6563),
    .B(n_1878),
    .Y(n_7396));
 AOI221x1_ASAP7_75t_SL g213013__5107 (.A1(n_3688),
    .A2(n_6730),
    .B1(n_6163),
    .B2(n_3963),
    .C(n_7134),
    .Y(n_7395));
 A2O1A1Ixp33_ASAP7_75t_L g213014__6260 (.A1(sa32[2]),
    .A2(n_6756),
    .B(n_6900),
    .C(n_1873),
    .Y(n_7394));
 AOI221xp5_ASAP7_75t_SL g213015__4319 (.A1(n_6750),
    .A2(n_2163),
    .B1(n_6615),
    .B2(n_2264),
    .C(n_7007),
    .Y(n_7393));
 OAI211xp5_ASAP7_75t_SL g213016__8428 (.A1(sa00[2]),
    .A2(n_6704),
    .B(n_7107),
    .C(sa00[5]),
    .Y(n_7392));
 AOI31xp33_ASAP7_75t_SL g213017__5526 (.A1(n_6828),
    .A2(n_6805),
    .A3(n_2693),
    .B(n_6521),
    .Y(n_7391));
 NAND2xp5_ASAP7_75t_SL g213018__6783 (.A(n_7212),
    .B(n_7302),
    .Y(n_7390));
 OAI21xp33_ASAP7_75t_L g213019__3680 (.A1(n_6973),
    .A2(n_7054),
    .B(n_8994),
    .Y(n_7389));
 OAI221xp5_ASAP7_75t_SL g213020__1617 (.A1(n_6613),
    .A2(n_2625),
    .B1(n_6746),
    .B2(n_2626),
    .C(n_7009),
    .Y(n_7388));
 OAI311xp33_ASAP7_75t_SL g213021__2802 (.A1(n_6220),
    .A2(n_6020),
    .A3(n_5865),
    .B1(n_6690),
    .C1(n_7104),
    .Y(n_7387));
 OA21x2_ASAP7_75t_SL g213022__1705 (.A1(n_3680),
    .A2(n_6729),
    .B(n_7290),
    .Y(n_7386));
 OAI211xp5_ASAP7_75t_SL g213023__5122 (.A1(n_6219),
    .A2(n_6574),
    .B(n_7117),
    .C(n_6678),
    .Y(n_7385));
 AOI221xp5_ASAP7_75t_SL g213024__8246 (.A1(n_6762),
    .A2(n_2224),
    .B1(n_6606),
    .B2(n_2180),
    .C(n_7126),
    .Y(n_7384));
 OAI211xp5_ASAP7_75t_SL g213025__7098 (.A1(n_2125),
    .A2(n_6609),
    .B(n_7012),
    .C(n_6910),
    .Y(n_7383));
 AOI21xp5_ASAP7_75t_SL g213026__6131 (.A1(n_7079),
    .A2(n_2718),
    .B(n_7018),
    .Y(n_7382));
 A2O1A1Ixp33_ASAP7_75t_SL g213027__1881 (.A1(n_6916),
    .A2(n_6844),
    .B(n_2688),
    .C(n_7214),
    .Y(n_7381));
 AOI21xp5_ASAP7_75t_SL g213028__5115 (.A1(n_6917),
    .A2(n_7137),
    .B(n_7048),
    .Y(n_7380));
 NAND4xp25_ASAP7_75t_SL g213029__7482 (.A(n_6791),
    .B(n_6913),
    .C(n_7051),
    .D(n_6627),
    .Y(n_7379));
 OAI211xp5_ASAP7_75t_SL g213030__4733 (.A1(n_2272),
    .A2(n_6614),
    .B(n_7006),
    .C(n_7037),
    .Y(n_7378));
 OAI21xp33_ASAP7_75t_SL g213031__6161 (.A1(n_7045),
    .A2(n_6861),
    .B(n_6871),
    .Y(n_7377));
 OAI211xp5_ASAP7_75t_SL g213032__9315 (.A1(n_2565),
    .A2(n_6618),
    .B(n_7068),
    .C(n_7166),
    .Y(n_7376));
 OAI211xp5_ASAP7_75t_SL g213033__9945 (.A1(n_2595),
    .A2(n_6620),
    .B(n_7164),
    .C(n_7064),
    .Y(n_7375));
 OAI221xp5_ASAP7_75t_SL g213034__2883 (.A1(n_6363),
    .A2(n_2164),
    .B1(n_6503),
    .B2(n_2582),
    .C(n_7284),
    .Y(n_7374));
 OAI21xp5_ASAP7_75t_SL g213035__2346 (.A1(n_7111),
    .A2(n_6676),
    .B(n_1879),
    .Y(n_7373));
 AOI211x1_ASAP7_75t_SL g213036__1666 (.A1(n_6947),
    .A2(n_2094),
    .B(n_7172),
    .C(n_6780),
    .Y(n_7372));
 AOI221xp5_ASAP7_75t_SL g213037__7410 (.A1(n_6747),
    .A2(n_2632),
    .B1(n_6611),
    .B2(n_2649),
    .C(n_7108),
    .Y(n_7371));
 NAND3xp33_ASAP7_75t_SL g213038__6417 (.A(n_6841),
    .B(n_7127),
    .C(n_7040),
    .Y(n_7370));
 AND4x1_ASAP7_75t_SL g213039__5477 (.A(n_6681),
    .B(n_6956),
    .C(n_6687),
    .D(n_6437),
    .Y(n_7369));
 O2A1O1Ixp33_ASAP7_75t_SL g213040__2398 (.A1(n_6671),
    .A2(n_1510),
    .B(n_6294),
    .C(n_2361),
    .Y(n_7368));
 OA22x2_ASAP7_75t_SL g213041__5107 (.A1(n_2363),
    .A2(n_6997),
    .B1(n_8207),
    .B2(n_7200),
    .Y(n_7367));
 NAND3xp33_ASAP7_75t_SL g213042__6260 (.A(n_7094),
    .B(n_6840),
    .C(n_7041),
    .Y(n_7366));
 OAI211xp5_ASAP7_75t_SL g213043__4319 (.A1(n_1700),
    .A2(n_6440),
    .B(n_6986),
    .C(n_7027),
    .Y(n_7365));
 NAND4xp25_ASAP7_75t_SL g213044__8428 (.A(n_7056),
    .B(n_6789),
    .C(n_6764),
    .D(n_6925),
    .Y(n_7364));
 OA331x1_ASAP7_75t_SL g213045__5526 (.A1(n_5963),
    .A2(n_2190),
    .A3(n_8209),
    .B1(n_6744),
    .B2(n_2541),
    .B3(n_8209),
    .C1(n_7186),
    .Y(n_7363));
 NAND3xp33_ASAP7_75t_SL g213046__6783 (.A(n_6763),
    .B(n_7011),
    .C(n_7028),
    .Y(n_7362));
 OAI221xp5_ASAP7_75t_SL g213047__3680 (.A1(n_7113),
    .A2(n_7061),
    .B1(n_6130),
    .B2(n_3445),
    .C(n_6980),
    .Y(n_7361));
 OAI321xp33_ASAP7_75t_SL g213048__1617 (.A1(n_6970),
    .A2(n_6416),
    .A3(sa12[0]),
    .B1(n_2610),
    .B2(n_6093),
    .C(n_6811),
    .Y(n_7360));
 OAI311xp33_ASAP7_75t_SL g213049__2802 (.A1(n_6215),
    .A2(n_6511),
    .A3(n_5157),
    .B1(n_6865),
    .C1(n_7067),
    .Y(n_7359));
 AOI221x1_ASAP7_75t_SL g213050__1705 (.A1(n_3673),
    .A2(n_6737),
    .B1(n_6701),
    .B2(n_6648),
    .C(n_7152),
    .Y(n_7358));
 AOI321xp33_ASAP7_75t_SL g213051__5122 (.A1(n_6960),
    .A2(n_6902),
    .A3(n_2687),
    .B1(n_6752),
    .B2(n_3404),
    .C(n_6728),
    .Y(n_7357));
 A2O1A1Ixp33_ASAP7_75t_SL g213052__8246 (.A1(sa12[2]),
    .A2(n_6431),
    .B(n_7123),
    .C(n_6623),
    .Y(n_7356));
 AOI311xp33_ASAP7_75t_SL g213053__7098 (.A1(n_5887),
    .A2(n_6533),
    .A3(n_2678),
    .B(n_7201),
    .C(n_6683),
    .Y(n_7355));
 AOI321xp33_ASAP7_75t_SL g213054__6131 (.A1(n_6950),
    .A2(n_6346),
    .A3(n_2595),
    .B1(n_2652),
    .B2(n_1857),
    .C(sa02[5]),
    .Y(n_7354));
 A2O1A1Ixp33_ASAP7_75t_SL g213055__1881 (.A1(n_1495),
    .A2(n_6668),
    .B(n_8188),
    .C(n_2661),
    .Y(n_7353));
 AOI221x1_ASAP7_75t_SL g213056__5115 (.A1(n_6567),
    .A2(n_3466),
    .B1(n_7180),
    .B2(n_2682),
    .C(n_7175),
    .Y(n_7352));
 OAI221xp5_ASAP7_75t_SL g213057__7482 (.A1(n_6769),
    .A2(n_5179),
    .B1(n_6265),
    .B2(n_2628),
    .C(n_7177),
    .Y(n_7351));
 OAI211xp5_ASAP7_75t_SL g213058__4733 (.A1(n_2125),
    .A2(n_6946),
    .B(n_7161),
    .C(n_6777),
    .Y(n_7350));
 AOI221xp5_ASAP7_75t_SL g213059__6161 (.A1(n_6761),
    .A2(n_1608),
    .B1(n_6625),
    .B2(n_2094),
    .C(n_7010),
    .Y(n_7349));
 AOI221x1_ASAP7_75t_SL g213060__9315 (.A1(n_6605),
    .A2(n_3568),
    .B1(n_2369),
    .B2(n_7057),
    .C(n_7198),
    .Y(n_7348));
 AO21x1_ASAP7_75t_SL g213061__9945 (.A1(n_2696),
    .A2(n_7147),
    .B(n_7160),
    .Y(n_7347));
 OAI211xp5_ASAP7_75t_SL g213062__2883 (.A1(n_1696),
    .A2(n_6244),
    .B(n_7171),
    .C(n_6990),
    .Y(n_7346));
 OAI211xp5_ASAP7_75t_SL g213063__2346 (.A1(n_2272),
    .A2(n_6941),
    .B(n_7167),
    .C(n_6816),
    .Y(n_7345));
 NAND3xp33_ASAP7_75t_SL g213064__1666 (.A(n_7046),
    .B(n_7165),
    .C(n_6866),
    .Y(n_7344));
 NOR4xp75_ASAP7_75t_SL g213065__7410 (.A(n_7184),
    .B(n_6931),
    .C(n_6942),
    .D(n_6873),
    .Y(n_7343));
 OAI322xp33_ASAP7_75t_SL g213066__6417 (.A1(n_6721),
    .A2(n_6793),
    .A3(n_2359),
    .B1(n_3663),
    .B2(n_6662),
    .C1(n_6530),
    .C2(n_3661),
    .Y(n_7342));
 O2A1O1Ixp33_ASAP7_75t_SL g213067__5477 (.A1(n_6926),
    .A2(n_6887),
    .B(n_1509),
    .C(n_7049),
    .Y(n_7341));
 OAI211xp5_ASAP7_75t_SL g213068__2398 (.A1(n_2257),
    .A2(n_6944),
    .B(n_7150),
    .C(n_6767),
    .Y(n_7340));
 OAI211xp5_ASAP7_75t_SL g213069__5107 (.A1(n_2151),
    .A2(n_6924),
    .B(n_6772),
    .C(n_7008),
    .Y(n_7339));
 AOI221xp5_ASAP7_75t_SL g213070__6260 (.A1(n_6616),
    .A2(n_2630),
    .B1(n_6948),
    .B2(n_2649),
    .C(n_7162),
    .Y(n_7338));
 NAND4xp25_ASAP7_75t_SL g213071__4319 (.A(n_6957),
    .B(n_6536),
    .C(n_6150),
    .D(n_2687),
    .Y(n_7337));
 O2A1O1Ixp33_ASAP7_75t_L g213072__8428 (.A1(n_6846),
    .A2(n_6590),
    .B(n_2720),
    .C(n_7253),
    .Y(n_7336));
 OAI22xp5_ASAP7_75t_SL g213073__5526 (.A1(n_2359),
    .A2(n_6996),
    .B1(n_8190),
    .B2(n_7139),
    .Y(n_7335));
 OAI311xp33_ASAP7_75t_SL g213074__6783 (.A1(n_6499),
    .A2(n_5888),
    .A3(n_2661),
    .B1(n_7092),
    .C1(n_6679),
    .Y(n_7334));
 OAI22xp5_ASAP7_75t_SL g213075__3680 (.A1(n_2628),
    .A2(n_7026),
    .B1(n_2272),
    .B2(n_5900),
    .Y(n_7333));
 OAI221xp5_ASAP7_75t_SL g213076__1617 (.A1(n_6381),
    .A2(n_2190),
    .B1(n_6366),
    .B2(n_2238),
    .C(n_7226),
    .Y(n_7332));
 NAND4xp25_ASAP7_75t_SL g213077__2802 (.A(n_6934),
    .B(n_6781),
    .C(n_7185),
    .D(n_6412),
    .Y(n_7331));
 A2O1A1Ixp33_ASAP7_75t_SL g213078__1705 (.A1(n_6434),
    .A2(n_6696),
    .B(sa22[2]),
    .C(n_6965),
    .Y(n_7330));
 AOI321xp33_ASAP7_75t_SL g213079__5122 (.A1(n_6325),
    .A2(n_6770),
    .A3(n_1857),
    .B1(n_6619),
    .B2(n_2180),
    .C(n_6571),
    .Y(n_7329));
 OAI221xp5_ASAP7_75t_SL g213080__8246 (.A1(n_6742),
    .A2(n_5154),
    .B1(n_6242),
    .B2(n_2609),
    .C(n_7174),
    .Y(n_7328));
 AOI32xp33_ASAP7_75t_SL g213081__7098 (.A1(n_7159),
    .A2(n_6796),
    .A3(n_1865),
    .B1(n_6983),
    .B2(n_8209),
    .Y(n_7327));
 OAI211xp5_ASAP7_75t_SL g213082__6131 (.A1(sa21[0]),
    .A2(n_6992),
    .B(n_6869),
    .C(n_6845),
    .Y(n_7326));
 NAND4xp25_ASAP7_75t_SL g213083__1881 (.A(n_6959),
    .B(n_6518),
    .C(n_6072),
    .D(n_2689),
    .Y(n_7325));
 OAI21xp5_ASAP7_75t_SL g213084__5115 (.A1(sa30[2]),
    .A2(n_6988),
    .B(n_7017),
    .Y(n_7324));
 AOI221xp5_ASAP7_75t_SL g213085__7482 (.A1(n_7153),
    .A2(n_2707),
    .B1(n_6771),
    .B2(n_3399),
    .C(n_6968),
    .Y(n_7323));
 OAI221xp5_ASAP7_75t_SL g213086__4733 (.A1(n_7002),
    .A2(n_2706),
    .B1(n_6100),
    .B2(n_3408),
    .C(n_6876),
    .Y(n_7322));
 OAI311xp33_ASAP7_75t_SL g213087__6161 (.A1(n_6733),
    .A2(n_2582),
    .A3(n_2003),
    .B1(n_6814),
    .C1(n_7130),
    .Y(n_7321));
 AOI22xp33_ASAP7_75t_SL g213088__9315 (.A1(sa31[2]),
    .A2(n_7082),
    .B1(n_1926),
    .B2(n_6702),
    .Y(n_7320));
 AOI22xp5_ASAP7_75t_SL g213089__9945 (.A1(n_1532),
    .A2(n_7119),
    .B1(n_1533),
    .B2(n_6705),
    .Y(n_7319));
 AOI22xp5_ASAP7_75t_SL g213090__2883 (.A1(sa11[2]),
    .A2(n_6685),
    .B1(n_2005),
    .B2(n_6995),
    .Y(n_7318));
 OAI21xp5_ASAP7_75t_SL g213091__2346 (.A1(sa01[2]),
    .A2(n_6982),
    .B(n_7023),
    .Y(n_7317));
 OAI22xp33_ASAP7_75t_SL g213092__1666 (.A1(sa33[2]),
    .A2(n_7047),
    .B1(n_2582),
    .B2(n_6751),
    .Y(n_7316));
 NAND4xp25_ASAP7_75t_L g213093__7410 (.A(n_6731),
    .B(n_7042),
    .C(n_6856),
    .D(n_6476),
    .Y(n_7315));
 AOI22xp33_ASAP7_75t_SL g213094__6417 (.A1(sa32[2]),
    .A2(n_7076),
    .B1(n_1981),
    .B2(n_6703),
    .Y(n_7314));
 OAI221xp5_ASAP7_75t_SL g213095__5477 (.A1(n_7170),
    .A2(n_6803),
    .B1(n_6713),
    .B2(n_3452),
    .C(n_6712),
    .Y(n_7313));
 AOI322xp5_ASAP7_75t_SL g213096__2398 (.A1(n_7021),
    .A2(sa32[5]),
    .A3(n_1981),
    .B1(n_3674),
    .B2(n_6833),
    .C1(n_6638),
    .C2(n_3688),
    .Y(n_7312));
 OAI211xp5_ASAP7_75t_SL g213097__5107 (.A1(n_6222),
    .A2(n_6495),
    .B(n_7105),
    .C(n_6535),
    .Y(n_7311));
 OAI211xp5_ASAP7_75t_SL g213098__6260 (.A1(n_5958),
    .A2(n_6399),
    .B(n_7052),
    .C(n_6879),
    .Y(n_7310));
 OAI221xp5_ASAP7_75t_SL g213099__4319 (.A1(n_6361),
    .A2(n_2151),
    .B1(n_6525),
    .B2(n_2602),
    .C(n_7120),
    .Y(n_7309));
 OAI211xp5_ASAP7_75t_SL g213100__8428 (.A1(n_6224),
    .A2(n_6557),
    .B(n_7115),
    .C(n_6675),
    .Y(n_7308));
 AOI211xp5_ASAP7_75t_SL g213101__5526 (.A1(n_6564),
    .A2(n_6230),
    .B(n_7109),
    .C(n_6673),
    .Y(n_7307));
 A2O1A1Ixp33_ASAP7_75t_SL g213102__6783 (.A1(n_3774),
    .A2(n_6779),
    .B(n_6976),
    .C(n_6842),
    .Y(n_7306));
 OA331x1_ASAP7_75t_SL g213103__3680 (.A1(n_6806),
    .A2(n_8202),
    .A3(n_2183),
    .B1(n_6991),
    .B2(n_8202),
    .B3(sa00[2]),
    .C1(n_6783),
    .Y(n_7305));
 OAI21xp5_ASAP7_75t_SL g213104__1617 (.A1(n_6855),
    .A2(n_6398),
    .B(n_2682),
    .Y(n_7304));
 OAI311xp33_ASAP7_75t_SL g213105__2802 (.A1(n_6209),
    .A2(n_6246),
    .A3(n_5173),
    .B1(n_5582),
    .C1(n_6786),
    .Y(n_7303));
 A2O1A1Ixp33_ASAP7_75t_SL g213106__1705 (.A1(n_1870),
    .A2(n_6455),
    .B(n_6589),
    .C(n_2690),
    .Y(n_7302));
 NAND4xp25_ASAP7_75t_SL g213107__5122 (.A(n_6714),
    .B(n_6838),
    .C(n_6877),
    .D(n_6405),
    .Y(n_7301));
 OAI21xp5_ASAP7_75t_SL g213108__8246 (.A1(n_3411),
    .A2(n_6736),
    .B(n_6365),
    .Y(n_7300));
 NAND4xp25_ASAP7_75t_SL g213109__7098 (.A(n_6862),
    .B(n_6830),
    .C(n_6961),
    .D(n_6553),
    .Y(n_7299));
 OAI211xp5_ASAP7_75t_SL g213110__6131 (.A1(n_3663),
    .A2(n_6723),
    .B(n_6920),
    .C(n_6753),
    .Y(n_7298));
 OAI211xp5_ASAP7_75t_SL g213111__1881 (.A1(n_2665),
    .A2(n_6384),
    .B(n_6817),
    .C(n_6790),
    .Y(n_7297));
 A2O1A1Ixp33_ASAP7_75t_L g213112__5115 (.A1(n_1422),
    .A2(n_5480),
    .B(n_6670),
    .C(n_2653),
    .Y(n_7296));
 AOI311xp33_ASAP7_75t_L g213113__7482 (.A1(n_4162),
    .A2(n_2414),
    .A3(sa12[0]),
    .B(n_6565),
    .C(n_6914),
    .Y(n_7295));
 OAI21xp5_ASAP7_75t_SL g213114__4733 (.A1(n_6353),
    .A2(n_6694),
    .B(n_2687),
    .Y(n_7294));
 OAI211xp5_ASAP7_75t_SL g213115__6161 (.A1(n_2703),
    .A2(n_6951),
    .B(n_6808),
    .C(n_6698),
    .Y(n_7293));
 A2O1A1O1Ixp25_ASAP7_75t_SL g213116__9315 (.A1(n_1627),
    .A2(n_1781),
    .B(n_6317),
    .C(n_3579),
    .D(n_6082),
    .Y(n_7292));
 OA22x2_ASAP7_75t_SL g213117__9945 (.A1(n_6706),
    .A2(n_6886),
    .B1(n_3608),
    .B2(n_6732),
    .Y(n_7291));
 AOI332xp33_ASAP7_75t_SL g213118__2883 (.A1(n_5162),
    .A2(n_5257),
    .A3(n_5708),
    .B1(n_5206),
    .B2(n_5013),
    .B3(n_4093),
    .C1(n_5925),
    .C2(n_4886),
    .Y(n_7290));
 OAI22xp5_ASAP7_75t_SL g213119__2346 (.A1(n_3467),
    .A2(n_6709),
    .B1(n_3336),
    .B2(n_6655),
    .Y(n_7289));
 AOI221xp5_ASAP7_75t_SL g213120__1666 (.A1(n_6385),
    .A2(n_8203),
    .B1(n_1980),
    .B2(n_6441),
    .C(sa32[5]),
    .Y(n_7288));
 NAND4xp25_ASAP7_75t_SL g213121__7410 (.A(n_6979),
    .B(n_5740),
    .C(n_6145),
    .D(n_2721),
    .Y(n_7287));
 OAI211xp5_ASAP7_75t_SL g213122__6417 (.A1(n_6859),
    .A2(n_6804),
    .B(n_6885),
    .C(n_6966),
    .Y(n_7286));
 OAI21x1_ASAP7_75t_SL g213123__5477 (.A1(n_6870),
    .A2(n_6410),
    .B(n_2690),
    .Y(n_7285));
 AOI22xp33_ASAP7_75t_SL g213124__2398 (.A1(n_2264),
    .A2(n_6952),
    .B1(n_2664),
    .B2(n_6334),
    .Y(n_7284));
 OAI211xp5_ASAP7_75t_SL g213125__5107 (.A1(n_6800),
    .A2(n_6836),
    .B(n_6832),
    .C(n_6967),
    .Y(n_7283));
 O2A1O1Ixp33_ASAP7_75t_L g213126__6260 (.A1(n_1966),
    .A2(n_6515),
    .B(n_6292),
    .C(n_2363),
    .Y(n_7282));
 OAI211xp5_ASAP7_75t_SL g213127__4319 (.A1(n_6229),
    .A2(n_6531),
    .B(n_7128),
    .C(n_6680),
    .Y(n_7281));
 A2O1A1O1Ixp25_ASAP7_75t_SL g213128__8428 (.A1(n_5944),
    .A2(n_5672),
    .B(n_1866),
    .C(n_6296),
    .D(n_2699),
    .Y(n_7280));
 NAND3xp33_ASAP7_75t_L g213129__5526 (.A(n_6979),
    .B(n_2721),
    .C(n_1531),
    .Y(n_7279));
 OAI22xp5_ASAP7_75t_SL g213130__6783 (.A1(n_6725),
    .A2(n_3550),
    .B1(n_6478),
    .B2(n_3452),
    .Y(n_7278));
 AOI221xp5_ASAP7_75t_SL g213131__3680 (.A1(n_6595),
    .A2(n_2670),
    .B1(n_6718),
    .B2(n_2191),
    .C(n_6622),
    .Y(n_7277));
 OAI211xp5_ASAP7_75t_SL g213132__1617 (.A1(n_6227),
    .A2(n_6545),
    .B(n_7116),
    .C(n_6682),
    .Y(n_7276));
 AOI22xp33_ASAP7_75t_SL g213133__2802 (.A1(n_3456),
    .A2(n_6710),
    .B1(n_3403),
    .B2(n_6660),
    .Y(n_7275));
 A2O1A1Ixp33_ASAP7_75t_SL g213134__1705 (.A1(n_8217),
    .A2(n_6415),
    .B(n_6298),
    .C(n_2375),
    .Y(n_7274));
 AOI211xp5_ASAP7_75t_SL g213135__5122 (.A1(n_6394),
    .A2(n_2670),
    .B(n_6785),
    .C(n_6784),
    .Y(n_7273));
 A2O1A1Ixp33_ASAP7_75t_SL g213136__8246 (.A1(n_5967),
    .A2(n_6389),
    .B(n_3377),
    .C(n_6739),
    .Y(n_7272));
 OAI211xp5_ASAP7_75t_SL g213137__7098 (.A1(n_6481),
    .A2(n_8213),
    .B(n_2689),
    .C(n_6977),
    .Y(n_7271));
 OAI221xp5_ASAP7_75t_SL g213138__6131 (.A1(n_6377),
    .A2(n_2626),
    .B1(n_6351),
    .B2(n_2625),
    .C(n_7090),
    .Y(n_7270));
 OAI211xp5_ASAP7_75t_SL g213139__1881 (.A1(sa02[0]),
    .A2(n_6391),
    .B(n_6798),
    .C(n_2709),
    .Y(n_7269));
 AOI21xp5_ASAP7_75t_SL g213140__5115 (.A1(n_6776),
    .A2(sa01[0]),
    .B(n_6974),
    .Y(n_7268));
 OAI21xp5_ASAP7_75t_SL g213141__7482 (.A1(sa02[0]),
    .A2(n_6897),
    .B(n_7032),
    .Y(n_7267));
 A2O1A1Ixp33_ASAP7_75t_R g213142__4733 (.A1(n_1547),
    .A2(n_5521),
    .B(n_6795),
    .C(n_2615),
    .Y(n_7266));
 OAI21xp5_ASAP7_75t_SL g213143__6161 (.A1(n_1966),
    .A2(n_6899),
    .B(n_7034),
    .Y(n_7265));
 OAI211xp5_ASAP7_75t_L g213144__9315 (.A1(n_1966),
    .A2(n_6359),
    .B(n_6801),
    .C(n_2702),
    .Y(n_7264));
 OAI32xp33_ASAP7_75t_L g213145__9945 (.A1(n_5961),
    .A2(n_6241),
    .A3(n_1540),
    .B1(n_3760),
    .B2(n_6328),
    .Y(n_7263));
 O2A1O1Ixp33_ASAP7_75t_R g213146__2883 (.A1(n_5513),
    .A2(n_6295),
    .B(n_2152),
    .C(n_6473),
    .Y(n_7262));
 O2A1O1Ixp33_ASAP7_75t_L g213147__2346 (.A1(n_6497),
    .A2(sa30[0]),
    .B(n_6270),
    .C(n_2381),
    .Y(n_7261));
 AOI22xp33_ASAP7_75t_L g213148__1666 (.A1(n_5235),
    .A2(n_6969),
    .B1(sa22[2]),
    .B2(n_6271),
    .Y(n_7260));
 O2A1O1Ixp33_ASAP7_75t_SL g213149__7410 (.A1(sa01[2]),
    .A2(n_6566),
    .B(n_5243),
    .C(n_6649),
    .Y(n_7259));
 AOI322xp5_ASAP7_75t_L g213150__6417 (.A1(n_2402),
    .A2(n_2570),
    .A3(sa33[0]),
    .B1(n_6519),
    .B2(n_5880),
    .C1(n_6288),
    .C2(sa33[0]),
    .Y(n_7258));
 AOI211xp5_ASAP7_75t_SL g213152__5477 (.A1(n_6889),
    .A2(n_1965),
    .B(n_6792),
    .C(n_5012),
    .Y(n_7256));
 OAI21xp5_ASAP7_75t_SL g213153__2398 (.A1(n_3508),
    .A2(n_6141),
    .B(n_7096),
    .Y(n_7255));
 OAI221xp5_ASAP7_75t_SL g213154__5107 (.A1(sa22[0]),
    .A2(n_6735),
    .B1(n_6360),
    .B2(n_8217),
    .C(n_2375),
    .Y(n_7254));
 OAI21xp5_ASAP7_75t_SL g213155__6260 (.A1(n_3400),
    .A2(n_6745),
    .B(n_6724),
    .Y(n_7253));
 AOI322xp5_ASAP7_75t_SL g213156__4319 (.A1(n_5727),
    .A2(n_5158),
    .A3(n_3507),
    .B1(sa01[5]),
    .B2(n_6561),
    .C1(n_3399),
    .C2(n_6485),
    .Y(n_7252));
 AOI221xp5_ASAP7_75t_SL g213157__8428 (.A1(n_1494),
    .A2(n_6299),
    .B1(n_6819),
    .B2(n_1495),
    .C(n_1966),
    .Y(n_7251));
 A2O1A1Ixp33_ASAP7_75t_SL g213158__5526 (.A1(n_6258),
    .A2(n_6175),
    .B(n_2266),
    .C(n_6765),
    .Y(n_7250));
 A2O1A1Ixp33_ASAP7_75t_SL g213159__6783 (.A1(n_6107),
    .A2(n_6479),
    .B(n_1698),
    .C(n_6848),
    .Y(n_7249));
 OAI22xp5_ASAP7_75t_SL g213160__3680 (.A1(sa01[2]),
    .A2(n_6930),
    .B1(n_2602),
    .B2(n_6420),
    .Y(n_7248));
 NAND3xp33_ASAP7_75t_SL g213161__1617 (.A(n_7044),
    .B(n_6858),
    .C(n_6936),
    .Y(n_7247));
 NAND4xp25_ASAP7_75t_SL g213162__2802 (.A(n_6935),
    .B(n_6644),
    .C(n_6860),
    .D(n_6954),
    .Y(n_7246));
 AOI321xp33_ASAP7_75t_SL g213163__1705 (.A1(n_5617),
    .A2(n_3914),
    .A3(n_3945),
    .B1(n_6500),
    .B2(n_4245),
    .C(n_6243),
    .Y(n_7245));
 AND4x1_ASAP7_75t_SL g213164__5122 (.A(n_6955),
    .B(n_6809),
    .C(n_6940),
    .D(n_6459),
    .Y(n_7244));
 O2A1O1Ixp33_ASAP7_75t_SL g213165__8246 (.A1(n_5518),
    .A2(n_6254),
    .B(n_2202),
    .C(n_6850),
    .Y(n_7243));
 NAND2xp5_ASAP7_75t_SL g213166__7098 (.A(n_7030),
    .B(n_6984),
    .Y(n_7242));
 OR3x1_ASAP7_75t_SL g213167__6131 (.A(n_6824),
    .B(n_6722),
    .C(n_2376),
    .Y(n_7241));
 O2A1O1Ixp33_ASAP7_75t_L g213168__1881 (.A1(n_5495),
    .A2(n_6300),
    .B(n_2163),
    .C(n_6851),
    .Y(n_7240));
 AOI22xp33_ASAP7_75t_SL g213169__5115 (.A1(n_2630),
    .A2(n_6741),
    .B1(n_2649),
    .B2(n_6118),
    .Y(n_7239));
 AOI22xp5_ASAP7_75t_L g213170__7482 (.A1(sa01[2]),
    .A2(n_6757),
    .B1(n_1915),
    .B2(n_6607),
    .Y(n_7238));
 OAI22xp5_ASAP7_75t_SL g213171__4733 (.A1(n_3680),
    .A2(n_6634),
    .B1(n_3684),
    .B2(n_6813),
    .Y(n_7237));
 OAI22xp5_ASAP7_75t_SL g213172__6161 (.A1(n_2565),
    .A2(n_6641),
    .B1(n_2201),
    .B2(n_6818),
    .Y(n_7236));
 NAND2xp5_ASAP7_75t_L g213173__9315 (.A(n_7156),
    .B(n_6987),
    .Y(n_7235));
 O2A1O1Ixp33_ASAP7_75t_SL g213174__9945 (.A1(n_6352),
    .A2(n_6198),
    .B(sa11[2]),
    .C(n_6904),
    .Y(n_7234));
 AOI21xp5_ASAP7_75t_SL g213175__2883 (.A1(n_6758),
    .A2(sa22[2]),
    .B(n_6911),
    .Y(n_7233));
 AOI22xp5_ASAP7_75t_SL g213176__2346 (.A1(n_2599),
    .A2(n_6716),
    .B1(n_2259),
    .B2(n_5869),
    .Y(n_7232));
 AOI22xp33_ASAP7_75t_SL g213177__1666 (.A1(n_1532),
    .A2(n_6754),
    .B1(n_1533),
    .B2(n_6604),
    .Y(n_7231));
 A2O1A1Ixp33_ASAP7_75t_SL g213178__7410 (.A1(n_5712),
    .A2(n_6496),
    .B(n_3577),
    .C(n_6839),
    .Y(n_7230));
 AOI22xp5_ASAP7_75t_SL g213179__6417 (.A1(n_3631),
    .A2(n_6637),
    .B1(n_3618),
    .B2(n_6810),
    .Y(n_7229));
 OAI21xp5_ASAP7_75t_SL g213180__5477 (.A1(n_3576),
    .A2(n_6815),
    .B(n_11517),
    .Y(n_7228));
 AOI21xp5_ASAP7_75t_SL g213181__2398 (.A1(n_6693),
    .A2(n_2601),
    .B(n_6852),
    .Y(n_7227));
 AOI22xp33_ASAP7_75t_L g213182__5107 (.A1(n_6867),
    .A2(n_2542),
    .B1(n_6138),
    .B2(n_2670),
    .Y(n_7226));
 AOI222xp33_ASAP7_75t_SL g213183__6260 (.A1(n_5724),
    .A2(n_3444),
    .B1(n_6656),
    .B2(n_3353),
    .C1(n_5615),
    .C2(n_3444),
    .Y(n_7225));
 AOI221xp5_ASAP7_75t_SL g213184__4319 (.A1(n_6504),
    .A2(n_2005),
    .B1(n_6568),
    .B2(sa11[2]),
    .C(n_2723),
    .Y(n_7224));
 AO21x1_ASAP7_75t_SL g213185__8428 (.A1(n_1968),
    .A2(n_6903),
    .B(n_7069),
    .Y(n_7223));
 AOI321xp33_ASAP7_75t_SL g213186__5526 (.A1(n_4479),
    .A2(n_3509),
    .A3(n_2398),
    .B1(n_6707),
    .B2(n_3509),
    .C(n_6822),
    .Y(n_7222));
 AOI221xp5_ASAP7_75t_SL g213187__6783 (.A1(n_6277),
    .A2(n_1915),
    .B1(n_6548),
    .B2(sa01[2]),
    .C(n_2701),
    .Y(n_7221));
 AOI211xp5_ASAP7_75t_SL g213188__3680 (.A1(n_6528),
    .A2(n_6240),
    .B(n_7176),
    .C(n_6880),
    .Y(n_7220));
 AO221x1_ASAP7_75t_SL g213189__1617 (.A1(n_6891),
    .A2(n_1870),
    .B1(n_6355),
    .B2(sa30[0]),
    .C(n_2381),
    .Y(n_7219));
 AOI211xp5_ASAP7_75t_SL g213190__2802 (.A1(n_6527),
    .A2(n_6239),
    .B(n_7178),
    .C(n_6883),
    .Y(n_7218));
 AOI21xp5_ASAP7_75t_SL g213191__1705 (.A1(n_6797),
    .A2(n_3568),
    .B(n_7131),
    .Y(n_7217));
 AOI211xp5_ASAP7_75t_SL g213192__5122 (.A1(n_6759),
    .A2(n_3631),
    .B(n_6918),
    .C(n_6669),
    .Y(n_7216));
 OAI211xp5_ASAP7_75t_SL g213193__8246 (.A1(n_6651),
    .A2(n_6172),
    .B(n_6686),
    .C(n_6592),
    .Y(n_7215));
 AOI21xp5_ASAP7_75t_SL g213194__7098 (.A1(n_6748),
    .A2(n_3403),
    .B(n_6939),
    .Y(n_7214));
 AOI22xp33_ASAP7_75t_SL g213195__6131 (.A1(n_1877),
    .A2(n_6672),
    .B1(n_6144),
    .B2(n_5962),
    .Y(n_7213));
 AOI22xp33_ASAP7_75t_SL g213196__1881 (.A1(n_3353),
    .A2(n_6755),
    .B1(n_3444),
    .B2(n_6514),
    .Y(n_7212));
 AOI221xp5_ASAP7_75t_SL g213197__5115 (.A1(n_6249),
    .A2(n_2615),
    .B1(n_6558),
    .B2(n_2624),
    .C(n_6505),
    .Y(n_7211));
 AOI22xp33_ASAP7_75t_SL g213198__7482 (.A1(n_6719),
    .A2(n_6199),
    .B1(sa11[0]),
    .B2(n_6326),
    .Y(n_7210));
 AO332x1_ASAP7_75t_SL g213199__4733 (.A1(n_6028),
    .A2(n_5502),
    .A3(n_6146),
    .B1(n_2546),
    .B2(n_1349),
    .B3(n_1980),
    .C1(n_6245),
    .C2(n_1980),
    .Y(n_7209));
 OA211x2_ASAP7_75t_SL g213200__6161 (.A1(n_3359),
    .A2(n_6749),
    .B(n_6972),
    .C(n_6766),
    .Y(n_7208));
 OAI322xp33_ASAP7_75t_SL g213201__9315 (.A1(n_6190),
    .A2(n_6010),
    .A3(n_4940),
    .B1(n_6274),
    .B2(n_1857),
    .C1(n_3602),
    .C2(n_4532),
    .Y(n_7207));
 AOI332xp33_ASAP7_75t_SL g213202__9945 (.A1(n_6349),
    .A2(n_5505),
    .A3(n_8217),
    .B1(n_1415),
    .B2(n_2548),
    .B3(sa22[0]),
    .C1(n_6251),
    .C2(sa22[0]),
    .Y(n_7206));
 AOI22xp5_ASAP7_75t_SL g213203__2883 (.A1(n_1869),
    .A2(n_6888),
    .B1(sa33[0]),
    .B2(n_6380),
    .Y(n_7205));
 AOI221xp5_ASAP7_75t_SL g213204__2346 (.A1(n_6309),
    .A2(n_1925),
    .B1(n_6794),
    .B2(sa21[2]),
    .C(n_2717),
    .Y(n_7204));
 OAI21xp33_ASAP7_75t_L g213205__1666 (.A1(n_8196),
    .A2(n_6324),
    .B(n_6825),
    .Y(n_7203));
 AO21x1_ASAP7_75t_SL g213206__7410 (.A1(n_3568),
    .A2(n_6419),
    .B(n_6893),
    .Y(n_7202));
 NAND2xp5_ASAP7_75t_SL g213207__6417 (.A(n_6414),
    .B(n_6689),
    .Y(n_7201));
 AOI21xp5_ASAP7_75t_SL g213208__5477 (.A1(n_6463),
    .A2(n_2566),
    .B(n_6875),
    .Y(n_7200));
 O2A1O1Ixp33_ASAP7_75t_SL g213209__2398 (.A1(n_1417),
    .A2(n_3875),
    .B(n_6460),
    .C(n_6493),
    .Y(n_7199));
 AOI21xp5_ASAP7_75t_L g213210__5107 (.A1(n_4937),
    .A2(n_6257),
    .B(n_3561),
    .Y(n_7198));
 OAI21xp33_ASAP7_75t_R g213211__6260 (.A1(n_6374),
    .A2(n_6190),
    .B(n_2034),
    .Y(n_7197));
 OAI21xp5_ASAP7_75t_L g213212__4319 (.A1(n_6358),
    .A2(n_6192),
    .B(n_1495),
    .Y(n_7196));
 OAI21xp33_ASAP7_75t_L g213213__8428 (.A1(n_6356),
    .A2(n_6194),
    .B(sa12[2]),
    .Y(n_7195));
 OAI31xp33_ASAP7_75t_R g213214__5526 (.A1(n_5491),
    .A2(n_5946),
    .A3(n_3822),
    .B(n_2608),
    .Y(n_7194));
 A2O1A1Ixp33_ASAP7_75t_L g213215__6783 (.A1(n_1346),
    .A2(n_5396),
    .B(n_6347),
    .C(sa33[2]),
    .Y(n_7193));
 NAND4xp25_ASAP7_75t_R g213216__3680 (.A(n_6148),
    .B(n_5971),
    .C(n_4841),
    .D(n_2034),
    .Y(n_7192));
 OAI21xp5_ASAP7_75t_SL g213217__1617 (.A1(n_6369),
    .A2(n_5881),
    .B(sa00[2]),
    .Y(n_7191));
 OAI22xp33_ASAP7_75t_SL g213218__2802 (.A1(sa00[0]),
    .A2(n_6520),
    .B1(n_4800),
    .B2(n_5802),
    .Y(n_7190));
 OAI31xp33_ASAP7_75t_L g213219__1705 (.A1(n_5996),
    .A2(n_6137),
    .A3(n_5416),
    .B(n_8196),
    .Y(n_7189));
 AOI31xp33_ASAP7_75t_L g213220__5122 (.A1(n_6078),
    .A2(n_5968),
    .A3(n_5250),
    .B(n_1510),
    .Y(n_7188));
 NAND3xp33_ASAP7_75t_L g213221__8246 (.A(n_6513),
    .B(n_2693),
    .C(n_8217),
    .Y(n_7187));
 OA33x2_ASAP7_75t_SL g213222__7098 (.A1(n_4838),
    .A2(n_5166),
    .A3(n_6059),
    .B1(n_3411),
    .B2(n_5223),
    .B3(n_6106),
    .Y(n_7186));
 OAI31xp33_ASAP7_75t_L g213223__6131 (.A1(n_5176),
    .A2(n_6142),
    .A3(n_1770),
    .B(n_2603),
    .Y(n_7185));
 AOI31xp33_ASAP7_75t_SL g213224__1881 (.A1(n_5936),
    .A2(n_4953),
    .A3(n_2750),
    .B(n_1696),
    .Y(n_7184));
 OAI21xp33_ASAP7_75t_SL g213225__5115 (.A1(n_6233),
    .A2(n_6450),
    .B(n_2566),
    .Y(n_7183));
 NAND2xp33_ASAP7_75t_R g213226__7482 (.A(n_2542),
    .B(n_6823),
    .Y(n_7182));
 OAI21xp33_ASAP7_75t_L g213227__4733 (.A1(n_5964),
    .A2(n_6237),
    .B(n_2034),
    .Y(n_7181));
 OAI22xp5_ASAP7_75t_SL g213228__6161 (.A1(sa21[0]),
    .A2(n_6508),
    .B1(n_5699),
    .B2(n_5743),
    .Y(n_7180));
 OAI22xp33_ASAP7_75t_SL g213229__9315 (.A1(n_2595),
    .A2(n_6439),
    .B1(n_2652),
    .B2(n_6501),
    .Y(n_7179));
 OAI21xp33_ASAP7_75t_SL g213230__9945 (.A1(n_2179),
    .A2(n_6429),
    .B(n_6667),
    .Y(n_7178));
 AOI22xp33_ASAP7_75t_SL g213231__2883 (.A1(n_2273),
    .A2(n_6368),
    .B1(n_4731),
    .B2(n_5559),
    .Y(n_7177));
 OAI21xp5_ASAP7_75t_SL g213232__2346 (.A1(n_2221),
    .A2(n_6428),
    .B(n_6234),
    .Y(n_7176));
 AOI31xp33_ASAP7_75t_SL g213233__1666 (.A1(n_6168),
    .A2(n_5896),
    .A3(n_4842),
    .B(n_3336),
    .Y(n_7175));
 AOI22xp33_ASAP7_75t_SL g213234__7410 (.A1(n_2267),
    .A2(n_6554),
    .B1(n_4721),
    .B2(n_5566),
    .Y(n_7174));
 A2O1A1Ixp33_ASAP7_75t_SL g213235__6417 (.A1(n_2135),
    .A2(n_5991),
    .B(n_6238),
    .C(n_2668),
    .Y(n_7173));
 NAND2xp5_ASAP7_75t_L g213236__5477 (.A(n_6923),
    .B(n_6778),
    .Y(n_7172));
 AOI22xp33_ASAP7_75t_SL g213237__2398 (.A1(n_2259),
    .A2(n_6432),
    .B1(n_4733),
    .B2(n_5569),
    .Y(n_7171));
 A2O1A1Ixp33_ASAP7_75t_L g213238__5107 (.A1(n_5194),
    .A2(n_5806),
    .B(n_1509),
    .C(n_2712),
    .Y(n_7170));
 AOI22xp33_ASAP7_75t_SL g213239__6260 (.A1(n_2542),
    .A2(n_6333),
    .B1(n_2191),
    .B2(n_6457),
    .Y(n_7169));
 OAI22xp33_ASAP7_75t_L g213240__4319 (.A1(sa33[0]),
    .A2(n_6362),
    .B1(n_1869),
    .B2(n_6166),
    .Y(n_7168));
 AOI22xp33_ASAP7_75t_SL g213241__8428 (.A1(n_2189),
    .A2(n_6383),
    .B1(n_2673),
    .B2(n_5863),
    .Y(n_7167));
 AOI22xp33_ASAP7_75t_SL g213242__5526 (.A1(n_2202),
    .A2(n_6407),
    .B1(n_2662),
    .B2(n_6342),
    .Y(n_7166));
 AOI22xp33_ASAP7_75t_SL g213243__6783 (.A1(n_2627),
    .A2(n_6393),
    .B1(n_2646),
    .B2(n_5861),
    .Y(n_7165));
 AOI22xp33_ASAP7_75t_SL g213244__3680 (.A1(n_2224),
    .A2(n_6408),
    .B1(n_2653),
    .B2(n_6341),
    .Y(n_7164));
 A2O1A1Ixp33_ASAP7_75t_SL g213245__1617 (.A1(n_5135),
    .A2(n_5536),
    .B(n_2204),
    .C(n_6588),
    .Y(n_7163));
 OAI22xp5_ASAP7_75t_SL g213246__2802 (.A1(n_2631),
    .A2(n_6409),
    .B1(n_2667),
    .B2(n_5862),
    .Y(n_7162));
 AOI22xp5_ASAP7_75t_SL g213247__1705 (.A1(n_2277),
    .A2(n_6403),
    .B1(n_2676),
    .B2(n_6329),
    .Y(n_7161));
 OAI21xp33_ASAP7_75t_SL g213248__5122 (.A1(n_6435),
    .A2(n_6171),
    .B(n_6734),
    .Y(n_7160));
 OAI21xp33_ASAP7_75t_L g213249__8246 (.A1(n_5895),
    .A2(n_6327),
    .B(n_5028),
    .Y(n_7159));
 A2O1A1Ixp33_ASAP7_75t_SL g213250__7098 (.A1(n_1404),
    .A2(n_5842),
    .B(n_5641),
    .C(n_3646),
    .Y(n_7158));
 AOI22xp5_ASAP7_75t_SL g213251__6131 (.A1(n_2629),
    .A2(n_6462),
    .B1(n_2673),
    .B2(n_6378),
    .Y(n_7157));
 AOI22xp33_ASAP7_75t_SL g213252__1881 (.A1(n_2611),
    .A2(n_6436),
    .B1(n_2679),
    .B2(n_6340),
    .Y(n_7156));
 O2A1O1Ixp33_ASAP7_75t_SL g213253__5115 (.A1(n_2187),
    .A2(n_3860),
    .B(n_6323),
    .C(sa11[0]),
    .Y(n_7155));
 A2O1A1Ixp33_ASAP7_75t_L g213254__7482 (.A1(n_2142),
    .A2(n_3913),
    .B(n_6322),
    .C(n_1968),
    .Y(n_7154));
 A2O1A1Ixp33_ASAP7_75t_SL g213255__4733 (.A1(n_6052),
    .A2(n_5787),
    .B(sa01[0]),
    .C(n_6585),
    .Y(n_7153));
 OAI33xp33_ASAP7_75t_SL g213256__6161 (.A1(n_4723),
    .A2(n_5994),
    .A3(n_5156),
    .B1(n_6105),
    .B2(n_5220),
    .B3(n_3377),
    .Y(n_7152));
 AOI22xp33_ASAP7_75t_SL g213257__9315 (.A1(n_2005),
    .A2(n_6549),
    .B1(sa11[2]),
    .B2(n_6512),
    .Y(n_7151));
 AOI22xp33_ASAP7_75t_SL g213258__9945 (.A1(n_1697),
    .A2(n_6647),
    .B1(n_6402),
    .B2(n_2678),
    .Y(n_7150));
 AOI31xp33_ASAP7_75t_SL g213259__2883 (.A1(n_4965),
    .A2(n_5854),
    .A3(n_1721),
    .B(n_1698),
    .Y(n_7149));
 O2A1O1Ixp33_ASAP7_75t_SL g213260__2346 (.A1(n_5735),
    .A2(n_6209),
    .B(n_3404),
    .C(n_6699),
    .Y(n_7148));
 OAI32xp33_ASAP7_75t_SL g213261__1666 (.A1(n_6129),
    .A2(n_5742),
    .A3(n_4253),
    .B1(n_6159),
    .B2(n_5680),
    .Y(n_7147));
 AOI211xp5_ASAP7_75t_SL g213262__7410 (.A1(n_6451),
    .A2(n_3378),
    .B(n_5701),
    .C(n_5629),
    .Y(n_7146));
 OAI22xp5_ASAP7_75t_L g213263__6417 (.A1(n_3550),
    .A2(n_6600),
    .B1(n_3577),
    .B2(n_6569),
    .Y(n_7145));
 O2A1O1Ixp33_ASAP7_75t_SL g213264__5477 (.A1(n_1434),
    .A2(n_3904),
    .B(n_6313),
    .C(sa30[0]),
    .Y(n_7144));
 O2A1O1Ixp33_ASAP7_75t_SL g213265__2398 (.A1(n_1590),
    .A2(n_4490),
    .B(n_6305),
    .C(n_3508),
    .Y(n_7143));
 AOI22xp5_ASAP7_75t_SL g213266__5107 (.A1(n_3410),
    .A2(n_6556),
    .B1(n_3583),
    .B2(n_6559),
    .Y(n_7142));
 A2O1A1Ixp33_ASAP7_75t_L g213267__6260 (.A1(n_1419),
    .A2(n_3878),
    .B(n_6306),
    .C(n_1869),
    .Y(n_7141));
 OAI31xp33_ASAP7_75t_SL g213268__4319 (.A1(n_5610),
    .A2(n_5408),
    .A3(n_4242),
    .B(n_2258),
    .Y(n_7140));
 AOI22xp33_ASAP7_75t_SL g213269__8428 (.A1(n_2611),
    .A2(n_6390),
    .B1(n_1608),
    .B2(n_5826),
    .Y(n_7139));
 A2O1A1Ixp33_ASAP7_75t_SL g213270__5526 (.A1(n_1444),
    .A2(n_3887),
    .B(n_6307),
    .C(n_1857),
    .Y(n_7138));
 OA21x2_ASAP7_75t_SL g213271__6783 (.A1(sa00[2]),
    .A2(n_6540),
    .B(n_2721),
    .Y(n_7137));
 O2A1O1Ixp33_ASAP7_75t_R g213272__3680 (.A1(n_5696),
    .A2(n_6222),
    .B(n_3544),
    .C(n_6584),
    .Y(n_7136));
 AOI21xp5_ASAP7_75t_SL g213273__1617 (.A1(n_6304),
    .A2(n_1527),
    .B(n_6583),
    .Y(n_7135));
 OAI22xp5_ASAP7_75t_SL g213274__2802 (.A1(n_5155),
    .A2(n_6438),
    .B1(n_3400),
    .B2(n_6480),
    .Y(n_7134));
 AOI21xp5_ASAP7_75t_SL g213275__1705 (.A1(n_6290),
    .A2(n_2026),
    .B(n_2695),
    .Y(n_7133));
 O2A1O1Ixp33_ASAP7_75t_L g213276__5122 (.A1(n_4946),
    .A2(n_5571),
    .B(sa02[0]),
    .C(n_2708),
    .Y(n_7132));
 A2O1A1Ixp33_ASAP7_75t_SL g213277__8246 (.A1(n_2439),
    .A2(n_1766),
    .B(n_6452),
    .C(n_6575),
    .Y(n_7131));
 AOI33xp33_ASAP7_75t_SL g213278__7098 (.A1(n_4767),
    .A2(n_5159),
    .A3(n_5983),
    .B1(n_6098),
    .B2(n_5205),
    .B3(n_3409),
    .Y(n_7130));
 O2A1O1Ixp33_ASAP7_75t_L g213279__6131 (.A1(n_4947),
    .A2(n_5587),
    .B(n_1966),
    .C(n_2703),
    .Y(n_7129));
 AOI32xp33_ASAP7_75t_SL g213280__1881 (.A1(n_6003),
    .A2(n_6017),
    .A3(n_5199),
    .B1(n_5943),
    .B2(n_5143),
    .Y(n_7128));
 AOI22xp33_ASAP7_75t_SL g213281__5115 (.A1(n_6319),
    .A2(n_2671),
    .B1(n_6332),
    .B2(n_2599),
    .Y(n_7127));
 OAI22xp5_ASAP7_75t_L g213282__7482 (.A1(n_2652),
    .A2(n_6320),
    .B1(n_2595),
    .B2(n_6331),
    .Y(n_7126));
 OAI22xp5_ASAP7_75t_SL g213283__4733 (.A1(n_3595),
    .A2(n_6624),
    .B1(n_3352),
    .B2(n_6413),
    .Y(n_7125));
 O2A1O1Ixp33_ASAP7_75t_SL g213284__6161 (.A1(n_5932),
    .A2(n_5772),
    .B(n_8182),
    .C(n_6587),
    .Y(n_7124));
 A2O1A1Ixp33_ASAP7_75t_SL g213285 (.A1(n_5289),
    .A2(n_5705),
    .B(sa12[2]),
    .C(n_1965),
    .Y(n_7123));
 AOI32xp33_ASAP7_75t_SL g213286 (.A1(n_5893),
    .A2(n_2662),
    .A3(n_1878),
    .B1(n_5910),
    .B2(n_3578),
    .Y(n_7122));
 A2O1A1Ixp33_ASAP7_75t_SL g213287 (.A1(n_5688),
    .A2(n_1797),
    .B(n_2609),
    .C(n_6586),
    .Y(n_7121));
 AOI22xp5_ASAP7_75t_SL g213288 (.A1(n_2245),
    .A2(n_6663),
    .B1(n_2666),
    .B2(n_6335),
    .Y(n_7120));
 OAI221xp5_ASAP7_75t_L g213289 (.A1(n_5866),
    .A2(n_1496),
    .B1(n_4367),
    .B2(n_1378),
    .C(n_5463),
    .Y(n_7119));
 A2O1A1O1Ixp25_ASAP7_75t_SL g213290 (.A1(n_1461),
    .A2(n_5198),
    .B(n_4876),
    .C(sa00[0]),
    .D(sa00[2]),
    .Y(n_7118));
 O2A1O1Ixp33_ASAP7_75t_SL g213291 (.A1(n_1644),
    .A2(n_3950),
    .B(n_6109),
    .C(n_6697),
    .Y(n_7117));
 AOI32xp33_ASAP7_75t_SL g213292 (.A1(n_6043),
    .A2(n_5197),
    .A3(n_5040),
    .B1(n_6165),
    .B2(n_5149),
    .Y(n_7116));
 AOI32xp33_ASAP7_75t_SL g213293 (.A1(n_6021),
    .A2(n_5193),
    .A3(n_5332),
    .B1(n_5985),
    .B2(n_5144),
    .Y(n_7115));
 A2O1A1Ixp33_ASAP7_75t_R g213294 (.A1(n_1552),
    .A2(n_5401),
    .B(n_6386),
    .C(n_1528),
    .Y(n_7114));
 OAI31xp33_ASAP7_75t_L g213295 (.A1(n_5747),
    .A2(n_5470),
    .A3(n_4555),
    .B(n_2690),
    .Y(n_7113));
 AOI22xp5_ASAP7_75t_SL g213296 (.A1(n_3409),
    .A2(n_6524),
    .B1(n_3548),
    .B2(n_6464),
    .Y(n_7112));
 OAI22xp5_ASAP7_75t_SL g213297 (.A1(n_5032),
    .A2(n_6458),
    .B1(n_5180),
    .B2(n_5972),
    .Y(n_7111));
 AOI21xp5_ASAP7_75t_SL g213298 (.A1(n_6392),
    .A2(sa21[0]),
    .B(n_2681),
    .Y(n_7110));
 OAI33xp33_ASAP7_75t_SL g213299 (.A1(n_5190),
    .A2(n_5030),
    .A3(n_6039),
    .B1(n_5153),
    .B2(n_4864),
    .B3(n_5343),
    .Y(n_7109));
 A2O1A1Ixp33_ASAP7_75t_SL g213300 (.A1(n_5293),
    .A2(n_5812),
    .B(n_2667),
    .C(n_6895),
    .Y(n_7108));
 OAI21xp33_ASAP7_75t_L g213301 (.A1(n_6252),
    .A2(n_5886),
    .B(sa00[2]),
    .Y(n_7107));
 O2A1O1Ixp33_ASAP7_75t_L g213302 (.A1(n_2066),
    .A2(n_5456),
    .B(n_6284),
    .C(n_3452),
    .Y(n_7106));
 O2A1O1Ixp33_ASAP7_75t_SL g213303 (.A1(n_1637),
    .A2(n_3991),
    .B(n_6108),
    .C(n_6688),
    .Y(n_7105));
 AOI33xp33_ASAP7_75t_SL g213304 (.A1(n_5019),
    .A2(n_5203),
    .A3(n_6019),
    .B1(n_4911),
    .B2(n_4959),
    .B3(n_5171),
    .Y(n_7104));
 O2A1O1Ixp33_ASAP7_75t_L g213305 (.A1(n_4925),
    .A2(n_6002),
    .B(sa02[0]),
    .C(n_2708),
    .Y(n_7103));
 A2O1A1Ixp33_ASAP7_75t_SL g213306 (.A1(n_4942),
    .A2(n_5973),
    .B(n_1870),
    .C(n_2690),
    .Y(n_7102));
 A2O1A1O1Ixp25_ASAP7_75t_R g213307 (.A1(n_1400),
    .A2(n_4146),
    .B(n_5914),
    .C(sa00[0]),
    .D(n_2691),
    .Y(n_7101));
 A2O1A1Ixp33_ASAP7_75t_L g213308 (.A1(n_5000),
    .A2(n_5580),
    .B(n_8182),
    .C(n_2716),
    .Y(n_7100));
 A2O1A1Ixp33_ASAP7_75t_SL g213309 (.A1(n_4961),
    .A2(n_5982),
    .B(n_8213),
    .C(n_2689),
    .Y(n_7099));
 A2O1A1Ixp33_ASAP7_75t_SL g213310 (.A1(n_4951),
    .A2(n_5975),
    .B(n_8182),
    .C(n_2716),
    .Y(n_7098));
 A2O1A1Ixp33_ASAP7_75t_L g213311 (.A1(n_1633),
    .A2(n_5455),
    .B(n_6283),
    .C(n_3403),
    .Y(n_7097));
 A2O1A1Ixp33_ASAP7_75t_L g213312 (.A1(n_1668),
    .A2(n_5476),
    .B(n_6286),
    .C(n_3399),
    .Y(n_7096));
 OAI21xp33_ASAP7_75t_L g213313 (.A1(n_6510),
    .A2(n_6562),
    .B(n_1981),
    .Y(n_7095));
 O2A1O1Ixp33_ASAP7_75t_SL g213314 (.A1(n_5284),
    .A2(n_5814),
    .B(n_2684),
    .C(n_6894),
    .Y(n_7094));
 A2O1A1Ixp33_ASAP7_75t_L g213315 (.A1(n_2414),
    .A2(n_5462),
    .B(n_6280),
    .C(n_3404),
    .Y(n_7093));
 AOI22xp5_ASAP7_75t_SL g213316 (.A1(n_5038),
    .A2(n_6471),
    .B1(n_5686),
    .B2(n_5589),
    .Y(n_7092));
 OAI22xp5_ASAP7_75t_SL g213317 (.A1(n_2225),
    .A2(n_6345),
    .B1(n_6418),
    .B2(n_2179),
    .Y(n_7091));
 AOI322xp5_ASAP7_75t_SL g213318 (.A1(n_3650),
    .A2(n_2646),
    .A3(n_2103),
    .B1(n_2646),
    .B2(n_5803),
    .C1(n_6461),
    .C2(n_2615),
    .Y(n_7090));
 OAI21xp5_ASAP7_75t_SL g213319 (.A1(n_6544),
    .A2(n_6186),
    .B(n_6666),
    .Y(n_7089));
 AOI21xp33_ASAP7_75t_L g213320 (.A1(n_6297),
    .A2(n_8208),
    .B(sa02[0]),
    .Y(n_7088));
 OAI21xp5_ASAP7_75t_SL g213321 (.A1(n_5951),
    .A2(n_6397),
    .B(n_6388),
    .Y(n_7087));
 O2A1O1Ixp33_ASAP7_75t_L g213322 (.A1(n_2424),
    .A2(n_5471),
    .B(n_6275),
    .C(n_3336),
    .Y(n_7086));
 AOI22xp5_ASAP7_75t_SL g213323 (.A1(n_3399),
    .A2(n_6492),
    .B1(n_3544),
    .B2(n_6371),
    .Y(n_7085));
 O2A1O1Ixp33_ASAP7_75t_L g213324 (.A1(n_1568),
    .A2(n_5458),
    .B(n_6276),
    .C(n_3400),
    .Y(n_7084));
 A2O1A1O1Ixp25_ASAP7_75t_SL g213325 (.A1(n_1498),
    .A2(n_5160),
    .B(n_5035),
    .C(n_1980),
    .D(n_1873),
    .Y(n_7083));
 OAI221xp5_ASAP7_75t_R g213326 (.A1(n_6162),
    .A2(n_1933),
    .B1(n_3861),
    .B2(n_1548),
    .C(n_6205),
    .Y(n_7082));
 NAND3xp33_ASAP7_75t_SL g213328 (.A(n_6217),
    .B(n_6551),
    .C(n_1879),
    .Y(n_7080));
 OAI21xp5_ASAP7_75t_SL g213329 (.A1(sa21[0]),
    .A2(n_6482),
    .B(n_6268),
    .Y(n_7079));
 AOI21xp5_ASAP7_75t_L g213330 (.A1(n_6185),
    .A2(n_6267),
    .B(n_2244),
    .Y(n_7078));
 A2O1A1Ixp33_ASAP7_75t_SL g213331 (.A1(n_2044),
    .A2(n_5126),
    .B(n_6488),
    .C(n_2542),
    .Y(n_7077));
 OAI221xp5_ASAP7_75t_SL g213332 (.A1(n_5867),
    .A2(n_1499),
    .B1(n_4352),
    .B2(n_1560),
    .C(n_6208),
    .Y(n_7076));
 AOI322xp5_ASAP7_75t_SL g213333 (.A1(n_6086),
    .A2(n_5345),
    .A3(n_5201),
    .B1(n_3578),
    .B2(n_5593),
    .C1(n_6444),
    .C2(n_3646),
    .Y(n_7075));
 AO21x1_ASAP7_75t_SL g213334 (.A1(n_6272),
    .A2(n_6181),
    .B(n_2238),
    .Y(n_7074));
 A2O1A1Ixp33_ASAP7_75t_L g213335 (.A1(n_2077),
    .A2(n_5123),
    .B(n_6466),
    .C(n_2611),
    .Y(n_7073));
 AOI21xp5_ASAP7_75t_L g213336 (.A1(sa21[0]),
    .A2(n_6430),
    .B(n_2681),
    .Y(n_7072));
 A2O1A1Ixp33_ASAP7_75t_L g213337 (.A1(n_1431),
    .A2(n_5474),
    .B(n_6468),
    .C(n_2566),
    .Y(n_7071));
 AOI22xp5_ASAP7_75t_SL g213338 (.A1(n_6572),
    .A2(n_3953),
    .B1(n_3403),
    .B2(n_6310),
    .Y(n_7070));
 A2O1A1Ixp33_ASAP7_75t_SL g213339 (.A1(n_5044),
    .A2(n_5966),
    .B(n_1968),
    .C(n_2718),
    .Y(n_7069));
 OAI21xp33_ASAP7_75t_L g213340 (.A1(n_6264),
    .A2(n_5879),
    .B(n_2220),
    .Y(n_7068));
 AOI22xp33_ASAP7_75t_SL g213341 (.A1(n_2239),
    .A2(n_6626),
    .B1(n_4057),
    .B2(n_4747),
    .Y(n_7067));
 AOI22xp33_ASAP7_75t_SL g213342 (.A1(n_3401),
    .A2(n_6498),
    .B1(n_3584),
    .B2(n_6350),
    .Y(n_7066));
 A2O1A1Ixp33_ASAP7_75t_SL g213343 (.A1(n_1419),
    .A2(n_5507),
    .B(n_6484),
    .C(n_2581),
    .Y(n_7065));
 OAI21xp33_ASAP7_75t_L g213344 (.A1(n_6184),
    .A2(n_6262),
    .B(n_2180),
    .Y(n_7064));
 A2O1A1Ixp33_ASAP7_75t_R g213345 (.A1(n_5111),
    .A2(n_6232),
    .B(n_1877),
    .C(n_3227),
    .Y(n_7063));
 OAI21xp5_ASAP7_75t_SL g213346 (.A1(n_6628),
    .A2(n_6188),
    .B(n_6837),
    .Y(n_7062));
 O2A1O1Ixp33_ASAP7_75t_L g213347 (.A1(n_2621),
    .A2(n_5512),
    .B(n_6396),
    .C(n_1870),
    .Y(n_7061));
 O2A1O1Ixp33_ASAP7_75t_L g213348 (.A1(n_1694),
    .A2(n_5508),
    .B(n_6395),
    .C(n_1869),
    .Y(n_7060));
 OAI21xp33_ASAP7_75t_R g213349 (.A1(n_6256),
    .A2(n_6207),
    .B(n_2203),
    .Y(n_7059));
 OAI211xp5_ASAP7_75t_SL g213350 (.A1(n_5904),
    .A2(n_5654),
    .B(n_2184),
    .C(sa00[5]),
    .Y(n_7058));
 OAI21xp33_ASAP7_75t_SL g213351 (.A1(sa02[0]),
    .A2(n_6445),
    .B(n_6293),
    .Y(n_7057));
 OAI21xp5_ASAP7_75t_R g213352 (.A1(n_6281),
    .A2(n_6188),
    .B(n_2264),
    .Y(n_7056));
 A2O1A1Ixp33_ASAP7_75t_L g213353 (.A1(n_1559),
    .A2(n_5526),
    .B(n_6469),
    .C(n_2608),
    .Y(n_7055));
 O2A1O1Ixp33_ASAP7_75t_R g213354 (.A1(n_1703),
    .A2(n_5511),
    .B(n_6382),
    .C(n_8217),
    .Y(n_7054));
 OAI31xp33_ASAP7_75t_R g213355 (.A1(n_5449),
    .A2(n_5537),
    .A3(n_4142),
    .B(sa33[0]),
    .Y(n_7053));
 AOI22xp5_ASAP7_75t_L g213356 (.A1(n_4974),
    .A2(n_6489),
    .B1(n_5142),
    .B2(n_5988),
    .Y(n_7052));
 A2O1A1Ixp33_ASAP7_75t_L g213357 (.A1(n_1400),
    .A2(n_4454),
    .B(n_6472),
    .C(n_2184),
    .Y(n_7051));
 OAI32xp33_ASAP7_75t_SL g213358 (.A1(n_5169),
    .A2(n_6001),
    .A3(n_4735),
    .B1(n_5034),
    .B2(n_5970),
    .Y(n_7050));
 A2O1A1Ixp33_ASAP7_75t_SL g213359 (.A1(n_5760),
    .A2(n_6221),
    .B(n_2125),
    .C(n_6640),
    .Y(n_7049));
 OAI22xp5_ASAP7_75t_SL g213360 (.A1(n_3554),
    .A2(n_6635),
    .B1(n_3377),
    .B2(n_6094),
    .Y(n_7048));
 AOI22xp33_ASAP7_75t_SL g213361 (.A1(n_5247),
    .A2(n_6303),
    .B1(n_1869),
    .B2(n_6442),
    .Y(n_7047));
 OAI21xp5_ASAP7_75t_L g213362 (.A1(n_6266),
    .A2(n_6172),
    .B(n_2624),
    .Y(n_7046));
 OAI21xp33_ASAP7_75t_L g213363 (.A1(n_1532),
    .A2(n_6273),
    .B(n_1509),
    .Y(n_7045));
 AOI22xp5_ASAP7_75t_SL g213364 (.A1(n_2630),
    .A2(n_6507),
    .B1(n_2668),
    .B2(n_6509),
    .Y(n_7044));
 A2O1A1Ixp33_ASAP7_75t_SL g213365 (.A1(n_5819),
    .A2(n_6212),
    .B(n_3408),
    .C(n_6684),
    .Y(n_7043));
 A2O1A1Ixp33_ASAP7_75t_L g213366 (.A1(n_2865),
    .A2(n_3960),
    .B(n_6379),
    .C(n_2581),
    .Y(n_7042));
 A2O1A1Ixp33_ASAP7_75t_SL g213367 (.A1(n_1349),
    .A2(n_4434),
    .B(n_6483),
    .C(n_2251),
    .Y(n_7041));
 OAI31xp33_ASAP7_75t_L g213368 (.A1(n_5554),
    .A2(n_5148),
    .A3(n_5446),
    .B(n_2203),
    .Y(n_7040));
 AOI333xp33_ASAP7_75t_SL g213369 (.A1(n_5976),
    .A2(n_3925),
    .A3(n_4703),
    .B1(n_5949),
    .B2(n_5225),
    .B3(n_3430),
    .C1(n_5146),
    .C2(n_5993),
    .C3(n_4724),
    .Y(n_7039));
 OAI21xp33_ASAP7_75t_R g213370 (.A1(n_5885),
    .A2(n_6449),
    .B(n_2632),
    .Y(n_7038));
 A2O1A1Ixp33_ASAP7_75t_L g213371 (.A1(n_1625),
    .A2(n_4444),
    .B(n_6454),
    .C(n_2189),
    .Y(n_7037));
 A2O1A1Ixp33_ASAP7_75t_SL g213372 (.A1(n_5684),
    .A2(n_6223),
    .B(n_3585),
    .C(n_6632),
    .Y(n_7036));
 AOI221xp5_ASAP7_75t_R g213373 (.A1(n_5461),
    .A2(n_1449),
    .B1(n_6006),
    .B2(n_2211),
    .C(n_3820),
    .Y(n_7035));
 A2O1A1O1Ixp25_ASAP7_75t_SL g213374 (.A1(n_1934),
    .A2(n_5187),
    .B(n_4258),
    .C(n_1966),
    .D(n_5334),
    .Y(n_7034));
 O2A1O1Ixp33_ASAP7_75t_SL g213375 (.A1(n_5703),
    .A2(n_6218),
    .B(n_3557),
    .C(n_6630),
    .Y(n_7033));
 A2O1A1O1Ixp25_ASAP7_75t_L g213376 (.A1(n_3034),
    .A2(n_1405),
    .B(n_5950),
    .C(sa02[0]),
    .D(n_5042),
    .Y(n_7032));
 AOI221xp5_ASAP7_75t_SL g213377 (.A1(n_5894),
    .A2(n_2132),
    .B1(n_2979),
    .B2(n_1370),
    .C(n_6523),
    .Y(n_7031));
 AOI22xp33_ASAP7_75t_SL g213378 (.A1(n_2601),
    .A2(n_6456),
    .B1(n_2676),
    .B2(n_6110),
    .Y(n_7030));
 AOI221xp5_ASAP7_75t_L g213379 (.A1(n_5940),
    .A2(n_1600),
    .B1(n_3103),
    .B2(n_1424),
    .C(n_5915),
    .Y(n_7029));
 A2O1A1Ixp33_ASAP7_75t_L g213380 (.A1(n_2421),
    .A2(n_1782),
    .B(n_6424),
    .C(n_2202),
    .Y(n_7028));
 AOI22xp33_ASAP7_75t_L g213381 (.A1(n_2649),
    .A2(n_6343),
    .B1(n_4737),
    .B2(n_5558),
    .Y(n_7027));
 AOI221xp5_ASAP7_75t_SL g213382 (.A1(n_5131),
    .A2(n_1435),
    .B1(n_5926),
    .B2(n_2751),
    .C(n_5470),
    .Y(n_7026));
 OAI221xp5_ASAP7_75t_L g213383 (.A1(n_6357),
    .A2(n_1509),
    .B1(n_3596),
    .B2(n_2847),
    .C(n_2362),
    .Y(n_7025));
 OAI22xp5_ASAP7_75t_SL g213384 (.A1(n_1924),
    .A2(n_6373),
    .B1(sa30[2]),
    .B2(n_6608),
    .Y(n_7024));
 AOI22xp33_ASAP7_75t_SL g213385 (.A1(n_2603),
    .A2(n_6645),
    .B1(n_2152),
    .B2(n_6099),
    .Y(n_7023));
 AOI22xp5_ASAP7_75t_SL g213386 (.A1(sa21[2]),
    .A2(n_6555),
    .B1(n_1925),
    .B2(n_6610),
    .Y(n_7022));
 OAI32xp33_ASAP7_75t_SL g213387 (.A1(n_6131),
    .A2(n_5084),
    .A3(n_5283),
    .B1(n_1980),
    .B2(n_6477),
    .Y(n_7021));
 AOI22xp5_ASAP7_75t_SL g213388 (.A1(n_2581),
    .A2(n_6642),
    .B1(n_2163),
    .B2(n_6315),
    .Y(n_7020));
 OAI21xp5_ASAP7_75t_SL g213389 (.A1(n_6629),
    .A2(n_6179),
    .B(n_6740),
    .Y(n_7019));
 OAI21xp5_ASAP7_75t_SL g213390 (.A1(n_3662),
    .A2(n_6287),
    .B(n_6821),
    .Y(n_7018));
 AOI22xp33_ASAP7_75t_SL g213391 (.A1(n_2629),
    .A2(n_6603),
    .B1(n_2189),
    .B2(n_6314),
    .Y(n_7017));
 AOI221xp5_ASAP7_75t_L g213392 (.A1(n_6157),
    .A2(n_1455),
    .B1(n_4348),
    .B2(n_2077),
    .C(n_6169),
    .Y(n_7016));
 AOI22xp5_ASAP7_75t_SL g213393 (.A1(n_2630),
    .A2(n_6643),
    .B1(n_2632),
    .B2(n_6312),
    .Y(n_7015));
 OAI21xp5_ASAP7_75t_SL g213394 (.A1(sa21[0]),
    .A2(n_6494),
    .B(n_3778),
    .Y(n_7014));
 A2O1A1Ixp33_ASAP7_75t_L g213395 (.A1(n_1981),
    .A2(n_5916),
    .B(n_5245),
    .C(n_6612),
    .Y(n_7013));
 AOI22xp5_ASAP7_75t_SL g213396 (.A1(n_2277),
    .A2(n_6401),
    .B1(n_2601),
    .B2(n_6330),
    .Y(n_7012));
 AOI22xp33_ASAP7_75t_SL g213397 (.A1(n_2662),
    .A2(n_6599),
    .B1(n_2566),
    .B2(n_5890),
    .Y(n_7011));
 OAI22xp33_ASAP7_75t_SL g213398 (.A1(n_2680),
    .A2(n_6598),
    .B1(n_2610),
    .B2(n_5892),
    .Y(n_7010));
 AOI22xp5_ASAP7_75t_SL g213399 (.A1(n_2646),
    .A2(n_6597),
    .B1(n_2615),
    .B2(n_5897),
    .Y(n_7009));
 AOI22xp33_ASAP7_75t_SL g213400 (.A1(n_2666),
    .A2(n_6596),
    .B1(n_2603),
    .B2(n_5903),
    .Y(n_7008));
 OAI22xp5_ASAP7_75t_SL g213401 (.A1(n_2663),
    .A2(n_6594),
    .B1(n_2582),
    .B2(n_6128),
    .Y(n_7007));
 AOI22xp5_ASAP7_75t_SL g213402 (.A1(n_2673),
    .A2(n_6593),
    .B1(n_2629),
    .B2(n_6127),
    .Y(n_7006));
 OAI22xp5_ASAP7_75t_SL g213403 (.A1(n_3377),
    .A2(n_6506),
    .B1(n_3554),
    .B2(n_6422),
    .Y(n_7005));
 AOI22xp33_ASAP7_75t_SL g213404 (.A1(n_6063),
    .A2(n_6636),
    .B1(n_1528),
    .B2(n_6302),
    .Y(n_7004));
 AOI32xp33_ASAP7_75t_SL g213405 (.A1(n_6560),
    .A2(n_2624),
    .A3(n_1895),
    .B1(n_6517),
    .B2(n_3403),
    .Y(n_7003));
 AOI22xp33_ASAP7_75t_SL g213406 (.A1(n_1540),
    .A2(n_6552),
    .B1(sa33[2]),
    .B2(n_6337),
    .Y(n_7002));
 OAI22xp5_ASAP7_75t_L g213407 (.A1(sa30[2]),
    .A2(n_6542),
    .B1(n_1924),
    .B2(n_6336),
    .Y(n_7001));
 OAI222xp33_ASAP7_75t_SL g213408 (.A1(n_5933),
    .A2(n_1599),
    .B1(n_5467),
    .B2(n_1639),
    .C1(n_1381),
    .C2(n_2991),
    .Y(n_7000));
 OAI22xp5_ASAP7_75t_L g213409 (.A1(n_6631),
    .A2(n_6182),
    .B1(n_5749),
    .B2(n_6080),
    .Y(n_6999));
 AOI222xp33_ASAP7_75t_L g213410 (.A1(n_5927),
    .A2(n_2200),
    .B1(n_3029),
    .B2(n_1581),
    .C1(n_5472),
    .C2(n_1451),
    .Y(n_6998));
 AOI32xp33_ASAP7_75t_L g213411 (.A1(n_6191),
    .A2(n_6011),
    .A3(n_4941),
    .B1(n_6316),
    .B2(n_1966),
    .Y(n_6997));
 AOI21xp5_ASAP7_75t_SL g213412 (.A1(n_6321),
    .A2(sa12[0]),
    .B(n_6829),
    .Y(n_6996));
 OAI222xp33_ASAP7_75t_SL g213413 (.A1(n_5954),
    .A2(n_2108),
    .B1(n_5477),
    .B2(n_1660),
    .C1(n_1344),
    .C2(n_2993),
    .Y(n_6995));
 AOI222xp33_ASAP7_75t_L g213414 (.A1(n_5476),
    .A2(n_2390),
    .B1(n_5898),
    .B2(n_2153),
    .C1(n_3054),
    .C2(n_1587),
    .Y(n_6994));
 AOI222xp33_ASAP7_75t_SL g213415 (.A1(n_5891),
    .A2(n_2136),
    .B1(n_1586),
    .B2(n_3105),
    .C1(n_5465),
    .C2(n_1436),
    .Y(n_6993));
 AOI32xp33_ASAP7_75t_SL g213416 (.A1(n_6338),
    .A2(n_8183),
    .A3(sa21[2]),
    .B1(n_6538),
    .B2(n_2682),
    .Y(n_6992));
 AOI22xp5_ASAP7_75t_SL g213417 (.A1(n_8196),
    .A2(n_6465),
    .B1(n_5938),
    .B2(n_6139),
    .Y(n_6991));
 OAI221xp5_ASAP7_75t_L g213418 (.A1(n_4284),
    .A2(n_2396),
    .B1(n_4324),
    .B2(n_2081),
    .C(n_6539),
    .Y(n_6990));
 AO21x1_ASAP7_75t_SL g213419 (.A1(n_6261),
    .A2(n_6176),
    .B(n_3226),
    .Y(n_6989));
 AOI332xp33_ASAP7_75t_SL g213420 (.A1(n_5987),
    .A2(n_5504),
    .A3(n_1870),
    .B1(n_1625),
    .B2(n_2552),
    .B3(sa30[0]),
    .C1(n_6235),
    .C2(sa30[0]),
    .Y(n_6988));
 AOI22xp5_ASAP7_75t_SL g213421 (.A1(n_1608),
    .A2(n_6400),
    .B1(n_2094),
    .B2(n_6425),
    .Y(n_6987));
 OAI221xp5_ASAP7_75t_SL g213422 (.A1(n_4308),
    .A2(n_1628),
    .B1(n_1355),
    .B2(n_3847),
    .C(n_6426),
    .Y(n_6986));
 OAI22xp5_ASAP7_75t_L g213423 (.A1(n_1509),
    .A2(n_6291),
    .B1(n_3596),
    .B2(n_4398),
    .Y(n_6985));
 AOI22xp5_ASAP7_75t_SL g213424 (.A1(n_2277),
    .A2(n_6387),
    .B1(n_2124),
    .B2(n_6427),
    .Y(n_6984));
 AOI221xp5_ASAP7_75t_L g213425 (.A1(n_6004),
    .A2(n_8182),
    .B1(n_5685),
    .B2(sa11[0]),
    .C(n_2937),
    .Y(n_6983));
 AOI332xp33_ASAP7_75t_SL g213426 (.A1(n_6231),
    .A2(n_4928),
    .A3(n_1877),
    .B1(n_2563),
    .B2(n_1668),
    .B3(sa01[0]),
    .C1(n_6269),
    .C2(sa01[0]),
    .Y(n_6982));
 AOI22xp5_ASAP7_75t_SL g213427 (.A1(n_2189),
    .A2(n_6364),
    .B1(n_2273),
    .B2(n_6423),
    .Y(n_6981));
 A2O1A1Ixp33_ASAP7_75t_L g213428 (.A1(n_1625),
    .A2(n_5466),
    .B(n_6279),
    .C(n_3353),
    .Y(n_6980));
 OAI31xp33_ASAP7_75t_SL g213429 (.A1(n_6005),
    .A2(n_3190),
    .A3(n_3038),
    .B(n_8213),
    .Y(n_6977));
 A2O1A1Ixp33_ASAP7_75t_SL g213430 (.A1(n_1498),
    .A2(n_5226),
    .B(n_6035),
    .C(n_2722),
    .Y(n_6976));
 OAI21xp33_ASAP7_75t_R g213431 (.A1(n_5124),
    .A2(n_6161),
    .B(n_2719),
    .Y(n_6975));
 OAI31xp33_ASAP7_75t_L g213432 (.A1(n_5214),
    .A2(n_5460),
    .A3(n_5331),
    .B(n_2707),
    .Y(n_6974));
 OAI21xp33_ASAP7_75t_L g213433 (.A1(n_5130),
    .A2(n_5873),
    .B(n_2693),
    .Y(n_6973));
 NAND3xp33_ASAP7_75t_SL g213434 (.A(n_5714),
    .B(n_5706),
    .C(n_2693),
    .Y(n_6972));
 A2O1A1Ixp33_ASAP7_75t_R g213435 (.A1(n_1500),
    .A2(n_5103),
    .B(n_5241),
    .C(sa21[0]),
    .Y(n_6971));
 AOI211xp5_ASAP7_75t_SL g213436 (.A1(n_5324),
    .A2(n_2077),
    .B(n_5846),
    .C(sa12[2]),
    .Y(n_6970));
 NAND2xp5_ASAP7_75t_L g213437 (.A(n_6529),
    .B(n_2026),
    .Y(n_6969));
 AOI21xp5_ASAP7_75t_R g213438 (.A1(n_5240),
    .A2(n_6120),
    .B(n_3508),
    .Y(n_6968));
 A2O1A1Ixp33_ASAP7_75t_L g213439 (.A1(n_3787),
    .A2(n_4277),
    .B(n_5695),
    .C(n_2191),
    .Y(n_6967));
 A2O1A1Ixp33_ASAP7_75t_L g213440 (.A1(n_3786),
    .A2(n_4294),
    .B(n_5683),
    .C(n_2163),
    .Y(n_6966));
 A2O1A1Ixp33_ASAP7_75t_SL g213441 (.A1(n_1395),
    .A2(n_4921),
    .B(n_5905),
    .C(n_2599),
    .Y(n_6965));
 AOI21xp5_ASAP7_75t_L g213442 (.A1(n_5664),
    .A2(n_5878),
    .B(n_1866),
    .Y(n_6964));
 O2A1O1Ixp33_ASAP7_75t_L g213443 (.A1(n_1560),
    .A2(n_5376),
    .B(n_5344),
    .C(n_1981),
    .Y(n_6963));
 A2O1A1Ixp33_ASAP7_75t_SL g213444 (.A1(n_1497),
    .A2(n_5359),
    .B(n_5906),
    .C(n_2601),
    .Y(n_6962));
 A2O1A1Ixp33_ASAP7_75t_SL g213445 (.A1(n_1547),
    .A2(n_5305),
    .B(n_5850),
    .C(n_2646),
    .Y(n_6961));
 NAND3xp33_ASAP7_75t_L g213446 (.A(n_6032),
    .B(n_1965),
    .C(n_5934),
    .Y(n_6960));
 A2O1A1Ixp33_ASAP7_75t_SL g213447 (.A1(sa31[6]),
    .A2(n_3830),
    .B(n_5586),
    .C(n_1866),
    .Y(n_6959));
 AOI211xp5_ASAP7_75t_L g213448 (.A1(n_5184),
    .A2(sa31[6]),
    .B(n_5025),
    .C(n_8213),
    .Y(n_6958));
 A2O1A1Ixp33_ASAP7_75t_R g213449 (.A1(n_1455),
    .A2(n_3823),
    .B(n_5590),
    .C(sa12[0]),
    .Y(n_6957));
 NAND2xp5_ASAP7_75t_L g213450 (.A(n_6223),
    .B(n_6490),
    .Y(n_6956));
 OAI21xp5_ASAP7_75t_L g213451 (.A1(n_4829),
    .A2(n_5939),
    .B(n_1697),
    .Y(n_6955));
 OAI31xp33_ASAP7_75t_L g213452 (.A1(n_4943),
    .A2(n_4762),
    .A3(n_3808),
    .B(n_2608),
    .Y(n_6954));
 A2O1A1Ixp33_ASAP7_75t_SL g213453 (.A1(n_1413),
    .A2(n_5272),
    .B(n_5560),
    .C(sa22[2]),
    .Y(n_6953));
 OAI211xp5_ASAP7_75t_L g213454 (.A1(n_2850),
    .A2(n_3061),
    .B(n_5588),
    .C(n_5525),
    .Y(n_6952));
 AOI22xp33_ASAP7_75t_SL g213455 (.A1(n_5576),
    .A2(n_5675),
    .B1(n_5541),
    .B2(n_5981),
    .Y(n_6951));
 A2O1A1Ixp33_ASAP7_75t_L g213456 (.A1(n_1405),
    .A2(n_5215),
    .B(n_5756),
    .C(n_1857),
    .Y(n_6950));
 A2O1A1Ixp33_ASAP7_75t_L g213457 (.A1(n_2421),
    .A2(n_5221),
    .B(n_5763),
    .C(n_8188),
    .Y(n_6949));
 NAND2xp5_ASAP7_75t_SL g213458 (.A(n_6263),
    .B(n_6180),
    .Y(n_6948));
 NAND2xp5_ASAP7_75t_SL g213459 (.A(n_6278),
    .B(n_1795),
    .Y(n_6947));
 NOR2xp33_ASAP7_75t_L g213460 (.A(n_6282),
    .B(n_6178),
    .Y(n_6946));
 O2A1O1Ixp33_ASAP7_75t_L g213461 (.A1(n_1491),
    .A2(n_2968),
    .B(n_5902),
    .C(n_2250),
    .Y(n_6945));
 NOR2xp33_ASAP7_75t_SL g213462 (.A(n_6255),
    .B(n_1794),
    .Y(n_6944));
 OAI21xp5_ASAP7_75t_SL g213463 (.A1(n_5236),
    .A2(n_5707),
    .B(n_1531),
    .Y(n_6979));
 A2O1A1O1Ixp25_ASAP7_75t_L g213464 (.A1(n_2456),
    .A2(n_3844),
    .B(n_1373),
    .C(n_5793),
    .D(n_3452),
    .Y(n_6943));
 AOI21xp5_ASAP7_75t_SL g213465 (.A1(n_5595),
    .A2(n_6054),
    .B(n_2260),
    .Y(n_6942));
 NOR2xp33_ASAP7_75t_SL g213466 (.A(n_6260),
    .B(n_6171),
    .Y(n_6941));
 OAI21xp33_ASAP7_75t_R g213467 (.A1(n_5607),
    .A2(n_6047),
    .B(n_2258),
    .Y(n_6940));
 AOI21xp33_ASAP7_75t_L g213468 (.A1(n_5246),
    .A2(n_6077),
    .B(n_3457),
    .Y(n_6939));
 A2O1A1O1Ixp25_ASAP7_75t_R g213469 (.A1(n_2439),
    .A2(n_4295),
    .B(n_2074),
    .C(n_5830),
    .D(n_3440),
    .Y(n_6938));
 NAND2xp5_ASAP7_75t_L g213470 (.A(n_5515),
    .B(n_6247),
    .Y(n_6937));
 OAI21xp33_ASAP7_75t_SL g213471 (.A1(n_5592),
    .A2(n_6000),
    .B(n_2632),
    .Y(n_6936));
 OAI21xp5_ASAP7_75t_SL g213472 (.A1(n_5913),
    .A2(n_5604),
    .B(n_2251),
    .Y(n_6935));
 OAI21xp33_ASAP7_75t_R g213473 (.A1(n_4903),
    .A2(n_5638),
    .B(n_2245),
    .Y(n_6934));
 A2O1A1O1Ixp25_ASAP7_75t_L g213474 (.A1(n_2450),
    .A2(n_4300),
    .B(n_1584),
    .C(n_5827),
    .D(n_3431),
    .Y(n_6933));
 A2O1A1O1Ixp25_ASAP7_75t_R g213475 (.A1(n_2481),
    .A2(n_4291),
    .B(n_1418),
    .C(n_5828),
    .D(n_3405),
    .Y(n_6932));
 AOI21xp5_ASAP7_75t_SL g213476 (.A1(n_5540),
    .A2(n_5919),
    .B(n_2204),
    .Y(n_6931));
 AOI22xp33_ASAP7_75t_SL g213477 (.A1(n_5728),
    .A2(n_5693),
    .B1(n_6053),
    .B2(n_5935),
    .Y(n_6930));
 A2O1A1Ixp33_ASAP7_75t_L g213478 (.A1(n_1935),
    .A2(n_5137),
    .B(n_5029),
    .C(n_1528),
    .Y(n_6978));
 OAI21xp33_ASAP7_75t_L g213479 (.A1(n_6122),
    .A2(n_5490),
    .B(n_2720),
    .Y(n_6929));
 AOI21xp33_ASAP7_75t_L g213480 (.A1(n_4944),
    .A2(n_5602),
    .B(n_1509),
    .Y(n_6928));
 A2O1A1Ixp33_ASAP7_75t_L g213481 (.A1(sa31[6]),
    .A2(n_5102),
    .B(n_5631),
    .C(n_1866),
    .Y(n_6927));
 A2O1A1Ixp33_ASAP7_75t_R g213482 (.A1(n_3748),
    .A2(n_5346),
    .B(n_1533),
    .C(n_5729),
    .Y(n_6926));
 A2O1A1Ixp33_ASAP7_75t_R g213483 (.A1(sa33[3]),
    .A2(n_2792),
    .B(n_5858),
    .C(n_2664),
    .Y(n_6925));
 AOI211xp5_ASAP7_75t_SL g213484 (.A1(n_4115),
    .A2(n_1587),
    .B(n_5625),
    .C(n_5520),
    .Y(n_6924));
 A2O1A1Ixp33_ASAP7_75t_L g213485 (.A1(n_1512),
    .A2(n_3275),
    .B(n_5859),
    .C(n_2679),
    .Y(n_6923));
 O2A1O1Ixp33_ASAP7_75t_L g213486 (.A1(n_1483),
    .A2(n_3081),
    .B(n_5822),
    .C(n_2183),
    .Y(n_6922));
 A2O1A1Ixp33_ASAP7_75t_R g213487 (.A1(n_1500),
    .A2(n_4463),
    .B(n_6089),
    .C(n_3559),
    .Y(n_6921));
 AOI33xp33_ASAP7_75t_SL g213488 (.A1(n_3928),
    .A2(n_5304),
    .A3(n_5354),
    .B1(n_6097),
    .B2(n_5229),
    .B3(n_3404),
    .Y(n_6920));
 A2O1A1Ixp33_ASAP7_75t_R g213489 (.A1(n_1497),
    .A2(n_4042),
    .B(n_6102),
    .C(n_2124),
    .Y(n_6919));
 O2A1O1Ixp33_ASAP7_75t_SL g213490 (.A1(n_1394),
    .A2(n_4740),
    .B(n_6096),
    .C(n_3359),
    .Y(n_6918));
 OAI211xp5_ASAP7_75t_SL g213491 (.A1(n_1417),
    .A2(n_5378),
    .B(n_5817),
    .C(sa00[2]),
    .Y(n_6917));
 OAI211xp5_ASAP7_75t_L g213492 (.A1(n_1722),
    .A2(n_2980),
    .B(n_6034),
    .C(n_4807),
    .Y(n_6916));
 O2A1O1Ixp33_ASAP7_75t_L g213493 (.A1(n_2351),
    .A2(n_4869),
    .B(n_5002),
    .C(sa31[2]),
    .Y(n_6915));
 A2O1A1Ixp33_ASAP7_75t_R g213494 (.A1(n_8702),
    .A2(n_4814),
    .B(n_1965),
    .C(n_2687),
    .Y(n_6914));
 OAI21xp5_ASAP7_75t_SL g213495 (.A1(n_5251),
    .A2(n_5821),
    .B(n_2678),
    .Y(n_6913));
 O2A1O1Ixp33_ASAP7_75t_SL g213496 (.A1(n_3476),
    .A2(n_4320),
    .B(n_2084),
    .C(n_6580),
    .Y(n_6912));
 O2A1O1Ixp33_ASAP7_75t_R g213497 (.A1(n_2353),
    .A2(n_4861),
    .B(n_5014),
    .C(sa22[2]),
    .Y(n_6911));
 A2O1A1Ixp33_ASAP7_75t_L g213498 (.A1(n_3767),
    .A2(n_3522),
    .B(n_5816),
    .C(n_2676),
    .Y(n_6910));
 A2O1A1Ixp33_ASAP7_75t_L g213499 (.A1(n_2364),
    .A2(n_4866),
    .B(n_5001),
    .C(n_8208),
    .Y(n_6909));
 A2O1A1Ixp33_ASAP7_75t_SL g213500 (.A1(n_2357),
    .A2(n_4931),
    .B(n_5006),
    .C(n_1531),
    .Y(n_6908));
 A2O1A1Ixp33_ASAP7_75t_R g213501 (.A1(n_2354),
    .A2(n_4855),
    .B(n_5010),
    .C(n_1540),
    .Y(n_6907));
 A2O1A1Ixp33_ASAP7_75t_R g213502 (.A1(n_2355),
    .A2(n_4893),
    .B(n_4988),
    .C(n_1494),
    .Y(n_6906));
 A2O1A1Ixp33_ASAP7_75t_L g213503 (.A1(n_2370),
    .A2(n_4889),
    .B(n_4992),
    .C(n_8199),
    .Y(n_6905));
 O2A1O1Ixp33_ASAP7_75t_SL g213504 (.A1(n_2368),
    .A2(n_4860),
    .B(n_5007),
    .C(sa11[2]),
    .Y(n_6904));
 OAI211xp5_ASAP7_75t_SL g213505 (.A1(n_2073),
    .A2(n_5356),
    .B(n_6155),
    .C(n_5443),
    .Y(n_6903));
 A2O1A1Ixp33_ASAP7_75t_L g213506 (.A1(n_2462),
    .A2(n_4022),
    .B(n_5839),
    .C(sa12[0]),
    .Y(n_6902));
 OAI21xp33_ASAP7_75t_SL g213507 (.A1(n_5734),
    .A2(n_6215),
    .B(n_3410),
    .Y(n_6901));
 O2A1O1Ixp33_ASAP7_75t_L g213508 (.A1(n_2302),
    .A2(n_3779),
    .B(n_5979),
    .C(sa32[2]),
    .Y(n_6900));
 O2A1O1Ixp33_ASAP7_75t_SL g213509 (.A1(n_3471),
    .A2(n_4303),
    .B(n_1586),
    .C(n_6579),
    .Y(n_6899));
 O2A1O1Ixp33_ASAP7_75t_L g213510 (.A1(n_1408),
    .A2(n_5378),
    .B(n_5825),
    .C(n_1698),
    .Y(n_6898));
 O2A1O1Ixp33_ASAP7_75t_R g213511 (.A1(n_3525),
    .A2(n_4282),
    .B(n_2075),
    .C(n_6578),
    .Y(n_6897));
 AOI21xp33_ASAP7_75t_R g213512 (.A1(n_6205),
    .A2(n_5824),
    .B(n_3510),
    .Y(n_6896));
 A2O1A1Ixp33_ASAP7_75t_SL g213513 (.A1(n_2142),
    .A2(n_2938),
    .B(n_5807),
    .C(n_2630),
    .Y(n_6895));
 O2A1O1Ixp33_ASAP7_75t_SL g213514 (.A1(n_2158),
    .A2(n_3108),
    .B(n_5810),
    .C(n_2609),
    .Y(n_6894));
 O2A1O1Ixp33_ASAP7_75t_L g213515 (.A1(sa02[7]),
    .A2(n_3059),
    .B(n_5601),
    .C(n_3561),
    .Y(n_6893));
 A2O1A1Ixp33_ASAP7_75t_L g213516 (.A1(n_1526),
    .A2(n_2981),
    .B(n_5600),
    .C(n_3575),
    .Y(n_6892));
 OAI211xp5_ASAP7_75t_SL g213517 (.A1(n_2078),
    .A2(n_5219),
    .B(n_6143),
    .C(n_5444),
    .Y(n_6891));
 O2A1O1Ixp33_ASAP7_75t_L g213518 (.A1(n_3407),
    .A2(n_4279),
    .B(n_1411),
    .C(n_6581),
    .Y(n_6890));
 A2O1A1Ixp33_ASAP7_75t_SL g213519 (.A1(n_1746),
    .A2(n_4301),
    .B(n_1418),
    .C(n_6582),
    .Y(n_6889));
 O2A1O1Ixp33_ASAP7_75t_SL g213520 (.A1(n_3345),
    .A2(n_4293),
    .B(n_1581),
    .C(n_6576),
    .Y(n_6888));
 OAI22xp5_ASAP7_75t_SL g213521 (.A1(n_1532),
    .A2(n_5855),
    .B1(n_3845),
    .B2(n_5306),
    .Y(n_6887));
 O2A1O1Ixp33_ASAP7_75t_SL g213522 (.A1(n_2170),
    .A2(n_3916),
    .B(n_5820),
    .C(n_1877),
    .Y(n_6886));
 OAI21xp33_ASAP7_75t_L g213523 (.A1(n_5835),
    .A2(n_6202),
    .B(n_2581),
    .Y(n_6885));
 OAI21xp33_ASAP7_75t_L g213524 (.A1(n_5064),
    .A2(n_5801),
    .B(n_3607),
    .Y(n_6884));
 O2A1O1Ixp33_ASAP7_75t_L g213525 (.A1(n_3333),
    .A2(n_3973),
    .B(n_6075),
    .C(n_2595),
    .Y(n_6883));
 OAI211xp5_ASAP7_75t_SL g213526 (.A1(n_2489),
    .A2(n_3078),
    .B(n_6173),
    .C(n_6069),
    .Y(n_6882));
 A2O1A1Ixp33_ASAP7_75t_SL g213527 (.A1(n_2458),
    .A2(n_4408),
    .B(n_2059),
    .C(n_6650),
    .Y(n_6881));
 O2A1O1Ixp33_ASAP7_75t_SL g213528 (.A1(n_3293),
    .A2(n_3971),
    .B(n_6066),
    .C(n_2565),
    .Y(n_6880));
 NAND3xp33_ASAP7_75t_L g213529 (.A(n_6067),
    .B(n_6225),
    .C(n_6037),
    .Y(n_6879));
 NAND3xp33_ASAP7_75t_L g213530 (.A(n_5738),
    .B(n_4557),
    .C(n_5484),
    .Y(n_6878));
 A2O1A1Ixp33_ASAP7_75t_L g213531 (.A1(n_2847),
    .A2(n_4126),
    .B(n_6087),
    .C(n_2124),
    .Y(n_6877));
 OAI21xp33_ASAP7_75t_L g213532 (.A1(n_5710),
    .A2(n_6226),
    .B(n_3548),
    .Y(n_6876));
 O2A1O1Ixp33_ASAP7_75t_L g213533 (.A1(sa13[7]),
    .A2(n_3060),
    .B(n_5597),
    .C(n_2201),
    .Y(n_6875));
 NOR2xp33_ASAP7_75t_L g213534 (.A(n_6211),
    .B(n_6406),
    .Y(n_6874));
 O2A1O1Ixp33_ASAP7_75t_SL g213535 (.A1(n_1602),
    .A2(n_3547),
    .B(n_5630),
    .C(n_2672),
    .Y(n_6873));
 AOI211xp5_ASAP7_75t_L g213536 (.A1(n_5209),
    .A2(n_2092),
    .B(n_6154),
    .C(n_5469),
    .Y(n_6872));
 NAND3xp33_ASAP7_75t_SL g213537 (.A(n_6177),
    .B(n_5736),
    .C(n_4650),
    .Y(n_6871));
 AOI211xp5_ASAP7_75t_R g213538 (.A1(n_4131),
    .A2(n_1625),
    .B(n_6048),
    .C(n_1870),
    .Y(n_6870));
 AO21x1_ASAP7_75t_L g213539 (.A1(n_5618),
    .A2(n_6228),
    .B(n_3558),
    .Y(n_6869));
 OAI211xp5_ASAP7_75t_R g213540 (.A1(n_3813),
    .A2(n_3995),
    .B(n_6200),
    .C(n_6033),
    .Y(n_6868));
 A2O1A1Ixp33_ASAP7_75t_L g213541 (.A1(n_3268),
    .A2(n_3380),
    .B(n_1850),
    .C(n_6602),
    .Y(n_6867));
 A2O1A1Ixp33_ASAP7_75t_L g213542 (.A1(n_1547),
    .A2(n_5414),
    .B(n_5723),
    .C(n_2615),
    .Y(n_6866));
 AOI22xp33_ASAP7_75t_SL g213543 (.A1(n_5579),
    .A2(n_5640),
    .B1(n_2542),
    .B2(n_5942),
    .Y(n_6865));
 AOI31xp33_ASAP7_75t_R g213544 (.A1(n_6026),
    .A2(n_4574),
    .A3(n_3188),
    .B(n_3595),
    .Y(n_6864));
 OAI21xp33_ASAP7_75t_L g213545 (.A1(n_5759),
    .A2(n_6182),
    .B(n_2239),
    .Y(n_6863));
 A2O1A1Ixp33_ASAP7_75t_L g213546 (.A1(n_2040),
    .A2(n_5379),
    .B(n_5769),
    .C(n_2627),
    .Y(n_6862));
 O2A1O1Ixp33_ASAP7_75t_SL g213547 (.A1(n_2066),
    .A2(n_4385),
    .B(n_5744),
    .C(n_1533),
    .Y(n_6861));
 OAI21xp33_ASAP7_75t_SL g213548 (.A1(n_5433),
    .A2(n_5808),
    .B(n_2267),
    .Y(n_6860));
 OAI21xp33_ASAP7_75t_R g213549 (.A1(n_5947),
    .A2(n_5623),
    .B(n_1540),
    .Y(n_6859));
 A2O1A1Ixp33_ASAP7_75t_SL g213550 (.A1(n_1545),
    .A2(n_4619),
    .B(n_6088),
    .C(n_2649),
    .Y(n_6858));
 OAI31xp33_ASAP7_75t_R g213551 (.A1(n_6016),
    .A2(n_4525),
    .A3(n_3203),
    .B(n_3557),
    .Y(n_6857));
 A2O1A1Ixp33_ASAP7_75t_R g213552 (.A1(n_2849),
    .A2(n_3960),
    .B(n_5754),
    .C(n_2264),
    .Y(n_6856));
 AOI211xp5_ASAP7_75t_SL g213553 (.A1(n_3913),
    .A2(n_1596),
    .B(n_6012),
    .C(n_1968),
    .Y(n_6855));
 NOR2xp33_ASAP7_75t_SL g213554 (.A(n_6654),
    .B(n_6184),
    .Y(n_6854));
 AOI21xp33_ASAP7_75t_R g213555 (.A1(n_4090),
    .A2(n_5783),
    .B(n_2179),
    .Y(n_6853));
 AOI21xp33_ASAP7_75t_R g213556 (.A1(n_5795),
    .A2(n_4067),
    .B(n_2125),
    .Y(n_6852));
 AOI21xp33_ASAP7_75t_R g213557 (.A1(n_5788),
    .A2(n_4066),
    .B(n_2265),
    .Y(n_6851));
 AOI21xp5_ASAP7_75t_R g213558 (.A1(n_4092),
    .A2(n_5791),
    .B(n_2221),
    .Y(n_6850));
 OAI21xp33_ASAP7_75t_R g213559 (.A1(n_4079),
    .A2(n_5792),
    .B(n_2624),
    .Y(n_6849));
 OAI21xp33_ASAP7_75t_L g213560 (.A1(n_4071),
    .A2(n_5799),
    .B(n_2258),
    .Y(n_6848));
 OAI21xp33_ASAP7_75t_R g213561 (.A1(n_4080),
    .A2(n_5780),
    .B(n_2239),
    .Y(n_6847));
 O2A1O1Ixp33_ASAP7_75t_SL g213562 (.A1(n_1567),
    .A2(n_5377),
    .B(n_5767),
    .C(n_1980),
    .Y(n_6846));
 A2O1A1Ixp33_ASAP7_75t_L g213563 (.A1(n_2523),
    .A2(n_2938),
    .B(n_5789),
    .C(n_3335),
    .Y(n_6845));
 A2O1A1Ixp33_ASAP7_75t_SL g213564 (.A1(n_2386),
    .A2(n_5380),
    .B(n_5768),
    .C(n_8213),
    .Y(n_6844));
 A2O1A1Ixp33_ASAP7_75t_L g213565 (.A1(n_1657),
    .A2(n_3057),
    .B(n_6090),
    .C(n_3410),
    .Y(n_6843));
 NAND3xp33_ASAP7_75t_SL g213566 (.A(n_6174),
    .B(n_5697),
    .C(n_4606),
    .Y(n_6842));
 A2O1A1Ixp33_ASAP7_75t_L g213567 (.A1(n_2397),
    .A2(n_5527),
    .B(n_4782),
    .C(n_2259),
    .Y(n_6841));
 AO21x1_ASAP7_75t_L g213568 (.A1(n_4781),
    .A2(n_6175),
    .B(n_2266),
    .Y(n_6840));
 OAI21xp33_ASAP7_75t_SL g213569 (.A1(n_5797),
    .A2(n_6201),
    .B(n_3549),
    .Y(n_6839));
 OAI21xp33_ASAP7_75t_SL g213570 (.A1(n_5761),
    .A2(n_6111),
    .B(n_2601),
    .Y(n_6838));
 NAND4xp25_ASAP7_75t_SL g213571 (.A(n_6101),
    .B(n_5369),
    .C(n_4105),
    .D(n_3409),
    .Y(n_6837));
 OAI21xp33_ASAP7_75t_SL g213572 (.A1(n_5955),
    .A2(n_5598),
    .B(n_2005),
    .Y(n_6836));
 OAI211xp5_ASAP7_75t_L g213573 (.A1(n_1373),
    .A2(n_3849),
    .B(n_6038),
    .C(n_4166),
    .Y(n_6835));
 AOI21xp5_ASAP7_75t_SL g213574 (.A1(n_5474),
    .A2(n_1436),
    .B(n_6487),
    .Y(n_6834));
 OAI221xp5_ASAP7_75t_SL g213575 (.A1(n_6040),
    .A2(n_4279),
    .B1(n_4519),
    .B2(n_1565),
    .C(n_6147),
    .Y(n_6833));
 OAI21xp33_ASAP7_75t_SL g213576 (.A1(n_5882),
    .A2(n_5782),
    .B(n_2542),
    .Y(n_6832));
 OAI21xp33_ASAP7_75t_SL g213578 (.A1(n_5687),
    .A2(n_6219),
    .B(n_2624),
    .Y(n_6830));
 NOR4xp25_ASAP7_75t_SL g213579 (.A(n_6194),
    .B(n_4844),
    .C(n_4917),
    .D(sa12[0]),
    .Y(n_6829));
 OAI31xp33_ASAP7_75t_R g213580 (.A1(n_5928),
    .A2(n_3005),
    .A3(n_3201),
    .B(n_8217),
    .Y(n_6828));
 NOR5xp2_ASAP7_75t_SL g213581 (.A(n_5253),
    .B(n_4534),
    .C(n_5370),
    .D(n_4065),
    .E(n_3402),
    .Y(n_6827));
 OAI31xp33_ASAP7_75t_SL g213582 (.A1(n_6008),
    .A2(n_3186),
    .A3(n_3019),
    .B(n_1509),
    .Y(n_6826));
 OAI221xp5_ASAP7_75t_L g213583 (.A1(n_1460),
    .A2(n_5387),
    .B1(n_4993),
    .B2(n_3245),
    .C(n_6029),
    .Y(n_6825));
 AOI21xp5_ASAP7_75t_SL g213584 (.A1(n_6232),
    .A2(n_5111),
    .B(n_1877),
    .Y(n_6824));
 AOI211xp5_ASAP7_75t_SL g213585 (.A1(n_3952),
    .A2(n_2485),
    .B(n_5716),
    .C(n_3457),
    .Y(n_6822));
 OAI21xp33_ASAP7_75t_L g213586 (.A1(n_5764),
    .A2(n_5884),
    .B(n_3579),
    .Y(n_6821));
 OAI21xp5_ASAP7_75t_R g213587 (.A1(n_5777),
    .A2(n_6229),
    .B(n_3583),
    .Y(n_6820));
 OAI221xp5_ASAP7_75t_SL g213588 (.A1(n_4672),
    .A2(n_2423),
    .B1(n_3008),
    .B2(n_2177),
    .C(n_5924),
    .Y(n_6819));
 AOI221xp5_ASAP7_75t_L g213589 (.A1(n_5050),
    .A2(n_1585),
    .B1(n_4496),
    .B2(n_2392),
    .C(n_4952),
    .Y(n_6818));
 OAI21xp5_ASAP7_75t_SL g213590 (.A1(n_5648),
    .A2(n_5064),
    .B(n_2603),
    .Y(n_6817));
 A2O1A1Ixp33_ASAP7_75t_L g213591 (.A1(n_1433),
    .A2(n_5429),
    .B(n_5647),
    .C(n_2629),
    .Y(n_6816));
 AOI221xp5_ASAP7_75t_SL g213592 (.A1(n_5062),
    .A2(n_2084),
    .B1(n_4513),
    .B2(n_1643),
    .C(n_4963),
    .Y(n_6815));
 NAND5xp2_ASAP7_75t_L g213593 (.A(n_5312),
    .B(n_5320),
    .C(n_3905),
    .D(sa33[5]),
    .E(n_2163),
    .Y(n_6814));
 AOI221xp5_ASAP7_75t_SL g213594 (.A1(n_1391),
    .A2(n_5067),
    .B1(n_4494),
    .B2(n_1641),
    .C(n_4976),
    .Y(n_6813));
 OAI211xp5_ASAP7_75t_SL g213595 (.A1(n_5990),
    .A2(n_5591),
    .B(n_2220),
    .C(n_1878),
    .Y(n_6812));
 OAI21xp33_ASAP7_75t_L g213596 (.A1(n_6227),
    .A2(n_5770),
    .B(n_2094),
    .Y(n_6811));
 OAI221xp5_ASAP7_75t_SL g213597 (.A1(n_4283),
    .A2(n_3793),
    .B1(n_5055),
    .B2(n_2081),
    .C(n_5188),
    .Y(n_6810));
 OAI211xp5_ASAP7_75t_SL g213598 (.A1(n_1654),
    .A2(n_4311),
    .B(n_6236),
    .C(n_6213),
    .Y(n_6809));
 OAI21xp33_ASAP7_75t_L g213599 (.A1(n_6056),
    .A2(n_6206),
    .B(n_3430),
    .Y(n_6808));
 AOI221xp5_ASAP7_75t_L g213600 (.A1(n_5063),
    .A2(n_1589),
    .B1(n_4544),
    .B2(n_1638),
    .C(n_4967),
    .Y(n_6807));
 AOI221xp5_ASAP7_75t_SL g213601 (.A1(n_5071),
    .A2(n_1572),
    .B1(n_4487),
    .B2(n_1652),
    .C(n_4964),
    .Y(n_6806));
 A2O1A1Ixp33_ASAP7_75t_L g213602 (.A1(n_1413),
    .A2(n_4128),
    .B(n_5999),
    .C(sa22[0]),
    .Y(n_6805));
 O2A1O1Ixp33_ASAP7_75t_L g213603 (.A1(n_1647),
    .A2(n_5437),
    .B(n_5917),
    .C(n_1869),
    .Y(n_6804));
 AOI211xp5_ASAP7_75t_L g213604 (.A1(n_2976),
    .A2(n_3396),
    .B(n_6045),
    .C(n_5920),
    .Y(n_6803));
 AOI221xp5_ASAP7_75t_R g213605 (.A1(n_4345),
    .A2(n_1550),
    .B1(n_6044),
    .B2(n_3284),
    .C(n_4910),
    .Y(n_6802));
 A2O1A1Ixp33_ASAP7_75t_L g213606 (.A1(n_2421),
    .A2(n_4138),
    .B(n_6027),
    .C(n_1966),
    .Y(n_6801));
 O2A1O1Ixp33_ASAP7_75t_SL g213607 (.A1(n_1656),
    .A2(n_5417),
    .B(n_5929),
    .C(n_8182),
    .Y(n_6800));
 OAI22xp33_ASAP7_75t_R g213608 (.A1(n_3391),
    .A2(n_6042),
    .B1(n_3189),
    .B2(n_4427),
    .Y(n_6799));
 A2O1A1Ixp33_ASAP7_75t_L g213609 (.A1(n_1605),
    .A2(n_1766),
    .B(n_6007),
    .C(sa02[0]),
    .Y(n_6798));
 OAI322xp33_ASAP7_75t_R g213610 (.A1(n_5330),
    .A2(n_5329),
    .A3(n_1458),
    .B1(n_4393),
    .B2(n_1389),
    .C1(n_2074),
    .C2(n_3148),
    .Y(n_6797));
 A2O1A1Ixp33_ASAP7_75t_R g213611 (.A1(sa11[6]),
    .A2(n_5170),
    .B(n_3795),
    .C(sa11[0]),
    .Y(n_6796));
 A2O1A1Ixp33_ASAP7_75t_L g213612 (.A1(n_2560),
    .A2(n_1634),
    .B(n_5923),
    .C(n_5475),
    .Y(n_6795));
 OAI21xp5_ASAP7_75t_SL g213613 (.A1(n_2424),
    .A2(n_5394),
    .B(n_6259),
    .Y(n_6794));
 O2A1O1Ixp33_ASAP7_75t_L g213614 (.A1(n_1651),
    .A2(n_5445),
    .B(n_5921),
    .C(n_1965),
    .Y(n_6793));
 O2A1O1Ixp33_ASAP7_75t_L g213615 (.A1(n_3555),
    .A2(n_2412),
    .B(n_5948),
    .C(n_1965),
    .Y(n_6792));
 OAI21xp33_ASAP7_75t_R g213616 (.A1(n_5612),
    .A2(n_1794),
    .B(n_2258),
    .Y(n_6791));
 A2O1A1Ixp33_ASAP7_75t_L g213617 (.A1(n_1638),
    .A2(n_4315),
    .B(n_5556),
    .C(n_2152),
    .Y(n_6790));
 OAI21xp33_ASAP7_75t_R g213618 (.A1(n_5726),
    .A2(n_6202),
    .B(n_2581),
    .Y(n_6789));
 OAI221xp5_ASAP7_75t_SL g213619 (.A1(n_5252),
    .A2(n_1379),
    .B1(n_5107),
    .B2(n_1935),
    .C(n_4843),
    .Y(n_6788));
 OAI221xp5_ASAP7_75t_L g213620 (.A1(n_4407),
    .A2(n_2501),
    .B1(n_4926),
    .B2(n_3381),
    .C(n_5311),
    .Y(n_6787));
 AOI221xp5_ASAP7_75t_SL g213621 (.A1(n_4612),
    .A2(n_2094),
    .B1(n_2984),
    .B2(n_1754),
    .C(n_6448),
    .Y(n_6786));
 O2A1O1Ixp33_ASAP7_75t_L g213622 (.A1(n_2045),
    .A2(n_5418),
    .B(n_5650),
    .C(n_2541),
    .Y(n_6785));
 O2A1O1Ixp33_ASAP7_75t_L g213623 (.A1(n_1662),
    .A2(n_4287),
    .B(n_5557),
    .C(n_2190),
    .Y(n_6784));
 A2O1A1Ixp33_ASAP7_75t_SL g213624 (.A1(n_1572),
    .A2(n_3875),
    .B(n_6055),
    .C(n_3673),
    .Y(n_6783));
 AOI21xp5_ASAP7_75t_R g213625 (.A1(n_5718),
    .A2(n_6197),
    .B(n_1696),
    .Y(n_6782));
 NAND4xp25_ASAP7_75t_L g213626 (.A(n_5635),
    .B(n_5127),
    .C(n_5076),
    .D(n_2666),
    .Y(n_6781));
 AOI21xp5_ASAP7_75t_L g213627 (.A1(n_5671),
    .A2(n_1796),
    .B(n_2610),
    .Y(n_6780));
 OAI221xp5_ASAP7_75t_SL g213628 (.A1(n_5265),
    .A2(n_1568),
    .B1(n_1773),
    .B2(n_2855),
    .C(n_5711),
    .Y(n_6779));
 A2O1A1Ixp33_ASAP7_75t_SL g213629 (.A1(n_8690),
    .A2(n_4292),
    .B(n_5538),
    .C(n_1608),
    .Y(n_6778));
 OAI21xp33_ASAP7_75t_L g213630 (.A1(n_5691),
    .A2(n_6201),
    .B(n_2601),
    .Y(n_6777));
 OAI211xp5_ASAP7_75t_SL g213631 (.A1(n_2606),
    .A2(n_5510),
    .B(n_5596),
    .C(n_4956),
    .Y(n_6776));
 NAND5xp2_ASAP7_75t_SL g213632 (.A(n_5261),
    .B(n_5249),
    .C(n_4704),
    .D(n_4526),
    .E(n_3378),
    .Y(n_6775));
 OAI21xp33_ASAP7_75t_R g213633 (.A1(n_6207),
    .A2(n_5922),
    .B(n_2599),
    .Y(n_6774));
 OAI211xp5_ASAP7_75t_L g213634 (.A1(n_2068),
    .A2(n_5125),
    .B(n_6117),
    .C(n_5506),
    .Y(n_6773));
 OAI21xp5_ASAP7_75t_SL g213635 (.A1(n_5667),
    .A2(n_6186),
    .B(n_2245),
    .Y(n_6772));
 OAI211xp5_ASAP7_75t_L g213636 (.A1(n_1463),
    .A2(n_5086),
    .B(n_5989),
    .C(n_4847),
    .Y(n_6771));
 A2O1A1Ixp33_ASAP7_75t_L g213637 (.A1(n_2464),
    .A2(n_4209),
    .B(n_2068),
    .C(n_6344),
    .Y(n_6770));
 NAND4xp25_ASAP7_75t_L g213638 (.A(n_5493),
    .B(n_5118),
    .C(n_5177),
    .D(n_2673),
    .Y(n_6769));
 OAI211xp5_ASAP7_75t_L g213639 (.A1(n_1546),
    .A2(n_4678),
    .B(n_6200),
    .C(n_6160),
    .Y(n_6768));
 A2O1A1Ixp33_ASAP7_75t_L g213640 (.A1(n_1653),
    .A2(n_4327),
    .B(n_5551),
    .C(n_2184),
    .Y(n_6767));
 AOI221xp5_ASAP7_75t_SL g213641 (.A1(n_4922),
    .A2(n_3382),
    .B1(n_4498),
    .B2(n_2936),
    .C(n_5775),
    .Y(n_6766));
 A2O1A1Ixp33_ASAP7_75t_R g213642 (.A1(n_1566),
    .A2(n_4325),
    .B(n_5568),
    .C(n_2251),
    .Y(n_6765));
 A2O1A1Ixp33_ASAP7_75t_L g213643 (.A1(n_1453),
    .A2(n_4297),
    .B(n_5562),
    .C(n_2163),
    .Y(n_6764));
 A2O1A1Ixp33_ASAP7_75t_SL g213644 (.A1(n_2392),
    .A2(n_5474),
    .B(n_5606),
    .C(n_2220),
    .Y(n_6763));
 OAI211xp5_ASAP7_75t_L g213645 (.A1(n_2434),
    .A2(n_4395),
    .B(n_5550),
    .C(n_5524),
    .Y(n_6762));
 OAI211xp5_ASAP7_75t_R g213646 (.A1(n_2412),
    .A2(n_4465),
    .B(n_5548),
    .C(n_5438),
    .Y(n_6761));
 OAI311xp33_ASAP7_75t_R g213647 (.A1(n_4279),
    .A2(n_1560),
    .A3(n_2620),
    .B1(n_4948),
    .C1(n_5583),
    .Y(n_6760));
 OAI21xp33_ASAP7_75t_L g213648 (.A1(n_1395),
    .A2(n_5845),
    .B(n_5663),
    .Y(n_6759));
 OAI211xp5_ASAP7_75t_SL g213649 (.A1(n_2053),
    .A2(n_4634),
    .B(n_5505),
    .C(n_5871),
    .Y(n_6758));
 OAI211xp5_ASAP7_75t_R g213650 (.A1(n_2057),
    .A2(n_4698),
    .B(n_5503),
    .C(n_6124),
    .Y(n_6757));
 OAI211xp5_ASAP7_75t_L g213651 (.A1(n_1560),
    .A2(n_4639),
    .B(n_5502),
    .C(n_5870),
    .Y(n_6756));
 OAI221xp5_ASAP7_75t_SL g213652 (.A1(n_5186),
    .A2(n_1640),
    .B1(n_5105),
    .B2(n_1367),
    .C(n_5164),
    .Y(n_6755));
 OAI211xp5_ASAP7_75t_L g213653 (.A1(n_1378),
    .A2(n_4679),
    .B(n_5868),
    .C(n_5501),
    .Y(n_6754));
 OAI211xp5_ASAP7_75t_R g213654 (.A1(n_2482),
    .A2(n_3928),
    .B(n_5719),
    .C(n_1737),
    .Y(n_6753));
 OAI221xp5_ASAP7_75t_SL g213655 (.A1(n_5075),
    .A2(n_1455),
    .B1(n_4162),
    .B2(n_1418),
    .C(n_5977),
    .Y(n_6752));
 O2A1O1Ixp33_ASAP7_75t_R g213656 (.A1(n_2787),
    .A2(n_4297),
    .B(n_1453),
    .C(n_6301),
    .Y(n_6751));
 OAI211xp5_ASAP7_75t_L g213657 (.A1(n_1646),
    .A2(n_4404),
    .B(n_5545),
    .C(n_5525),
    .Y(n_6750));
 AOI222xp33_ASAP7_75t_SL g213658 (.A1(n_5134),
    .A2(n_1399),
    .B1(n_5106),
    .B2(n_1844),
    .C1(n_4127),
    .C2(n_1424),
    .Y(n_6749));
 OAI221xp5_ASAP7_75t_SL g213659 (.A1(n_5165),
    .A2(n_1642),
    .B1(n_5101),
    .B2(sa31[6]),
    .C(n_5167),
    .Y(n_6748));
 OAI211xp5_ASAP7_75t_SL g213660 (.A1(n_1376),
    .A2(n_4377),
    .B(n_5546),
    .C(n_5500),
    .Y(n_6747));
 AOI211xp5_ASAP7_75t_L g213661 (.A1(n_4456),
    .A2(n_1633),
    .B(n_5549),
    .C(n_5530),
    .Y(n_6746));
 O2A1O1Ixp33_ASAP7_75t_SL g213662 (.A1(n_1729),
    .A2(n_4325),
    .B(n_1566),
    .C(n_6289),
    .Y(n_6745));
 AOI21xp5_ASAP7_75t_SL g213663 (.A1(n_5844),
    .A2(n_1850),
    .B(n_5655),
    .Y(n_6744));
 OAI221xp5_ASAP7_75t_SL g213664 (.A1(n_5479),
    .A2(n_1383),
    .B1(n_4546),
    .B2(n_1459),
    .C(n_6113),
    .Y(n_6743));
 NAND4xp25_ASAP7_75t_SL g213665 (.A(n_5141),
    .B(n_5419),
    .C(n_5492),
    .D(n_2684),
    .Y(n_6742));
 OAI211xp5_ASAP7_75t_SL g213666 (.A1(n_1541),
    .A2(n_5129),
    .B(n_6119),
    .C(n_5484),
    .Y(n_6741));
 NAND5xp2_ASAP7_75t_SL g213667 (.A(n_5189),
    .B(n_5341),
    .C(n_4537),
    .D(n_4181),
    .E(n_3335),
    .Y(n_6740));
 NOR2xp33_ASAP7_75t_SL g213668 (.A(n_6311),
    .B(n_5751),
    .Y(n_6739));
 OAI221xp5_ASAP7_75t_L g213669 (.A1(n_5448),
    .A2(n_1407),
    .B1(n_4652),
    .B2(n_1460),
    .C(n_6135),
    .Y(n_6738));
 OAI21xp5_ASAP7_75t_SL g213670 (.A1(n_1461),
    .A2(n_5843),
    .B(n_5662),
    .Y(n_6737));
 AOI21xp5_ASAP7_75t_R g213671 (.A1(n_5478),
    .A2(n_1657),
    .B(n_6285),
    .Y(n_6736));
 AOI221xp5_ASAP7_75t_SL g213672 (.A1(n_5200),
    .A2(n_2082),
    .B1(n_4373),
    .B2(n_1413),
    .C(n_6092),
    .Y(n_6735));
 NAND5xp2_ASAP7_75t_SL g213673 (.A(n_5262),
    .B(n_4690),
    .C(n_5287),
    .D(n_4204),
    .E(n_3353),
    .Y(n_6734));
 AOI222xp33_ASAP7_75t_L g213674 (.A1(n_5851),
    .A2(n_1839),
    .B1(n_4410),
    .B2(n_1451),
    .C1(n_3171),
    .C2(n_1581),
    .Y(n_6733));
 AOI21xp5_ASAP7_75t_SL g213675 (.A1(n_5849),
    .A2(n_1464),
    .B(n_5660),
    .Y(n_6732));
 NAND4xp25_ASAP7_75t_L g213676 (.A(n_6212),
    .B(n_5570),
    .C(n_5450),
    .D(n_2664),
    .Y(n_6731));
 OAI21xp5_ASAP7_75t_SL g213677 (.A1(n_1498),
    .A2(n_5836),
    .B(n_5659),
    .Y(n_6730));
 AOI21xp33_ASAP7_75t_L g213678 (.A1(n_1341),
    .A2(n_1938),
    .B(n_5656),
    .Y(n_6729));
 OAI221xp5_ASAP7_75t_SL g213679 (.A1(n_4901),
    .A2(n_3338),
    .B1(n_4493),
    .B2(n_1753),
    .C(n_5753),
    .Y(n_6728));
 OAI221xp5_ASAP7_75t_SL g213680 (.A1(n_5464),
    .A2(n_2423),
    .B1(n_4193),
    .B2(n_1404),
    .C(n_6151),
    .Y(n_6727));
 AOI221xp5_ASAP7_75t_R g213681 (.A1(n_5472),
    .A2(n_2404),
    .B1(n_4516),
    .B2(n_1346),
    .C(n_6152),
    .Y(n_6726));
 AOI222xp33_ASAP7_75t_SL g213682 (.A1(n_4503),
    .A2(n_1554),
    .B1(n_3698),
    .B2(n_2089),
    .C1(n_5852),
    .C2(n_1496),
    .Y(n_6725));
 AOI221xp5_ASAP7_75t_SL g213683 (.A1(n_4919),
    .A2(n_3358),
    .B1(n_4442),
    .B2(n_2926),
    .C(n_5748),
    .Y(n_6724));
 AOI222xp33_ASAP7_75t_SL g213684 (.A1(n_5841),
    .A2(n_1456),
    .B1(n_4488),
    .B2(n_8703),
    .C1(n_1370),
    .C2(n_3138),
    .Y(n_6723));
 OAI221xp5_ASAP7_75t_SL g213685 (.A1(n_1590),
    .A2(n_5151),
    .B1(n_4492),
    .B2(n_1666),
    .C(n_6091),
    .Y(n_6722));
 AOI211xp5_ASAP7_75t_SL g213686 (.A1(n_4831),
    .A2(n_1456),
    .B(n_5670),
    .C(sa12[0]),
    .Y(n_6721));
 AOI221xp5_ASAP7_75t_SL g213687 (.A1(n_4486),
    .A2(n_2918),
    .B1(n_4421),
    .B2(n_3211),
    .C(n_6318),
    .Y(n_6720));
 AOI211xp5_ASAP7_75t_L g213688 (.A1(n_4996),
    .A2(n_3268),
    .B(n_4852),
    .C(sa11[0]),
    .Y(n_6719));
 OAI21xp5_ASAP7_75t_L g213689 (.A1(n_1656),
    .A2(n_4450),
    .B(n_6547),
    .Y(n_6718));
 AOI221xp5_ASAP7_75t_SL g213690 (.A1(n_5461),
    .A2(n_1664),
    .B1(n_4396),
    .B2(n_1935),
    .C(n_5875),
    .Y(n_6717));
 AO21x1_ASAP7_75t_SL g213691 (.A1(n_1440),
    .A2(n_5527),
    .B(n_6470),
    .Y(n_6716));
 NAND4xp25_ASAP7_75t_L g213692 (.A(n_5577),
    .B(n_6214),
    .C(n_5117),
    .D(n_2646),
    .Y(n_6715));
 NAND4xp25_ASAP7_75t_SL g213693 (.A(n_5584),
    .B(n_5116),
    .C(n_5487),
    .D(n_2676),
    .Y(n_6714));
 AOI221xp5_ASAP7_75t_L g213694 (.A1(n_5065),
    .A2(n_1496),
    .B1(n_5175),
    .B2(n_1555),
    .C(n_4851),
    .Y(n_6713));
 AOI221xp5_ASAP7_75t_L g213695 (.A1(n_4918),
    .A2(n_3343),
    .B1(n_4438),
    .B2(n_3182),
    .C(n_5776),
    .Y(n_6712));
 OAI221xp5_ASAP7_75t_L g213696 (.A1(n_4484),
    .A2(n_2930),
    .B1(n_4467),
    .B2(sa02[1]),
    .C(n_6308),
    .Y(n_6711));
 OAI221xp5_ASAP7_75t_L g213697 (.A1(n_4455),
    .A2(n_1392),
    .B1(n_4478),
    .B2(n_1546),
    .C(n_5634),
    .Y(n_6710));
 AOI221xp5_ASAP7_75t_L g213698 (.A1(n_4376),
    .A2(n_1401),
    .B1(n_1781),
    .B2(n_1542),
    .C(n_5627),
    .Y(n_6709));
 OAI222xp33_ASAP7_75t_L g213699 (.A1(n_4495),
    .A2(n_3506),
    .B1(n_6073),
    .B2(n_3389),
    .C1(n_4448),
    .C2(n_1473),
    .Y(n_6708));
 OAI22xp33_ASAP7_75t_SL g213700 (.A1(sa31[6]),
    .A2(n_5856),
    .B1(n_1392),
    .B2(n_3726),
    .Y(n_6707));
 A2O1A1Ixp33_ASAP7_75t_SL g213701 (.A1(n_4828),
    .A2(n_5081),
    .B(sa01[0]),
    .C(n_4275),
    .Y(n_6706));
 OAI222xp33_ASAP7_75t_L g213702 (.A1(n_5953),
    .A2(n_2185),
    .B1(n_5456),
    .B2(n_1553),
    .C1(n_3117),
    .C2(n_1373),
    .Y(n_6705));
 AOI222xp33_ASAP7_75t_L g213703 (.A1(n_5941),
    .A2(n_2098),
    .B1(n_5447),
    .B2(n_1652),
    .C1(n_2987),
    .C2(n_1572),
    .Y(n_6704));
 OAI221xp5_ASAP7_75t_L g213704 (.A1(n_5937),
    .A2(n_2117),
    .B1(n_5458),
    .B2(n_1565),
    .C(n_4254),
    .Y(n_6703));
 OAI221xp5_ASAP7_75t_R g213705 (.A1(n_5930),
    .A2(n_2146),
    .B1(n_3033),
    .B2(n_2083),
    .C(n_6133),
    .Y(n_6702));
 O2A1O1Ixp33_ASAP7_75t_L g213706 (.A1(n_5416),
    .A2(n_4825),
    .B(n_8196),
    .C(n_4249),
    .Y(n_6701));
 OAI221xp5_ASAP7_75t_SL g213707 (.A1(n_3381),
    .A2(n_5637),
    .B1(n_4592),
    .B2(n_4407),
    .C(n_5239),
    .Y(n_6700));
 AO21x1_ASAP7_75t_SL g213708 (.A1(n_1737),
    .A2(n_5633),
    .B(n_5745),
    .Y(n_6699));
 AOI21xp33_ASAP7_75t_L g213709 (.A1(n_5553),
    .A2(n_3390),
    .B(n_5741),
    .Y(n_6698));
 AOI321xp33_ASAP7_75t_SL g213710 (.A1(n_4372),
    .A2(n_2386),
    .A3(n_3306),
    .B1(n_4059),
    .B2(n_2039),
    .C(n_6050),
    .Y(n_6697));
 OAI221xp5_ASAP7_75t_SL g213711 (.A1(n_3894),
    .A2(n_2053),
    .B1(n_3954),
    .B2(n_2141),
    .C(n_5730),
    .Y(n_6696));
 OAI21xp33_ASAP7_75t_L g213712 (.A1(n_2821),
    .A2(n_5614),
    .B(n_6121),
    .Y(n_6695));
 AOI221xp5_ASAP7_75t_SL g213713 (.A1(n_1609),
    .A2(n_3929),
    .B1(n_1765),
    .B2(n_2077),
    .C(n_5732),
    .Y(n_6694));
 OAI221xp5_ASAP7_75t_SL g213714 (.A1(n_5132),
    .A2(n_2047),
    .B1(n_4019),
    .B2(n_2580),
    .C(n_6051),
    .Y(n_6693));
 AOI22xp33_ASAP7_75t_R g213715 (.A1(n_3392),
    .A2(n_6041),
    .B1(n_2540),
    .B2(n_4425),
    .Y(n_6692));
 AOI221xp5_ASAP7_75t_L g213716 (.A1(n_5122),
    .A2(n_1447),
    .B1(n_1770),
    .B2(n_2564),
    .C(n_6049),
    .Y(n_6691));
 OAI211xp5_ASAP7_75t_L g213717 (.A1(n_1558),
    .A2(n_4570),
    .B(n_5682),
    .C(n_5271),
    .Y(n_6690));
 OAI321xp33_ASAP7_75t_SL g213718 (.A1(n_4344),
    .A2(n_3298),
    .A3(n_2411),
    .B1(n_1417),
    .B2(n_4030),
    .C(n_6030),
    .Y(n_6689));
 AOI321xp33_ASAP7_75t_L g213719 (.A1(n_4338),
    .A2(n_2824),
    .A3(n_2431),
    .B1(n_4115),
    .B2(n_1448),
    .C(n_6023),
    .Y(n_6688));
 OAI321xp33_ASAP7_75t_L g213720 (.A1(n_4379),
    .A2(n_2846),
    .A3(n_1567),
    .B1(n_1562),
    .B2(n_4167),
    .C(n_6014),
    .Y(n_6687));
 OAI221xp5_ASAP7_75t_SL g213721 (.A1(n_1791),
    .A2(n_1634),
    .B1(n_3032),
    .B2(n_2104),
    .C(n_5658),
    .Y(n_6686));
 OAI221xp5_ASAP7_75t_SL g213722 (.A1(n_5613),
    .A2(n_3269),
    .B1(n_3865),
    .B2(n_1450),
    .C(n_4950),
    .Y(n_6685));
 AOI21xp5_ASAP7_75t_SL g213723 (.A1(n_5621),
    .A2(n_3392),
    .B(n_5681),
    .Y(n_6684));
 AOI221xp5_ASAP7_75t_SL g213724 (.A1(n_3875),
    .A2(n_2055),
    .B1(n_1572),
    .B2(n_5391),
    .C(n_5653),
    .Y(n_6683));
 OAI221xp5_ASAP7_75t_SL g213725 (.A1(n_5389),
    .A2(n_2063),
    .B1(n_1765),
    .B2(n_1582),
    .C(n_5677),
    .Y(n_6682));
 OAI321xp33_ASAP7_75t_SL g213726 (.A1(n_4279),
    .A2(n_2091),
    .A3(n_2620),
    .B1(n_1562),
    .B2(n_3893),
    .C(n_5649),
    .Y(n_6681));
 OAI321xp33_ASAP7_75t_SL g213727 (.A1(n_4278),
    .A2(n_1344),
    .A3(n_2634),
    .B1(n_1450),
    .B2(n_3876),
    .C(n_5652),
    .Y(n_6680));
 OAI321xp33_ASAP7_75t_SL g213728 (.A1(n_4303),
    .A2(n_1584),
    .A3(n_2650),
    .B1(n_2059),
    .B2(n_3877),
    .C(n_5676),
    .Y(n_6679));
 OAI221xp5_ASAP7_75t_SL g213729 (.A1(n_5402),
    .A2(n_2083),
    .B1(n_3896),
    .B2(n_1546),
    .C(n_5669),
    .Y(n_6678));
 OR3x1_ASAP7_75t_SL g213730 (.A(n_5874),
    .B(n_4268),
    .C(n_3668),
    .Y(n_6677));
 AOI321xp33_ASAP7_75t_L g213731 (.A1(n_4284),
    .A2(n_1424),
    .A3(n_1704),
    .B1(n_3894),
    .B2(n_1440),
    .C(n_5603),
    .Y(n_6676));
 OAI221xp5_ASAP7_75t_L g213732 (.A1(n_5119),
    .A2(n_1381),
    .B1(n_3903),
    .B2(n_1434),
    .C(n_5666),
    .Y(n_6675));
 AOI221xp5_ASAP7_75t_L g213733 (.A1(n_5394),
    .A2(n_1356),
    .B1(n_3907),
    .B2(n_1545),
    .C(n_5678),
    .Y(n_6674));
 NOR3xp33_ASAP7_75t_SL g213734 (.A(n_4970),
    .B(n_5326),
    .C(n_5698),
    .Y(n_6673));
 OAI221xp5_ASAP7_75t_SL g213735 (.A1(n_4121),
    .A2(n_2868),
    .B1(n_3054),
    .B2(n_1588),
    .C(n_5957),
    .Y(n_6672));
 AOI221xp5_ASAP7_75t_R g213736 (.A1(n_4119),
    .A2(n_2867),
    .B1(n_3117),
    .B2(n_1366),
    .C(n_5945),
    .Y(n_6671));
 OAI22xp33_ASAP7_75t_L g213737 (.A1(n_2123),
    .A2(n_5959),
    .B1(n_2074),
    .B2(n_3163),
    .Y(n_6670));
 AOI211xp5_ASAP7_75t_SL g213738 (.A1(n_3955),
    .A2(n_2440),
    .B(n_5709),
    .C(n_3381),
    .Y(n_6669));
 OAI211xp5_ASAP7_75t_L g213739 (.A1(sa11[6]),
    .A2(n_5098),
    .B(n_5969),
    .C(n_4840),
    .Y(n_6823));
 NOR2xp33_ASAP7_75t_L g213740 (.A(n_6450),
    .B(n_6233),
    .Y(n_6668));
 OAI221xp5_ASAP7_75t_L g213741 (.A1(n_4546),
    .A2(n_2399),
    .B1(n_2803),
    .B2(n_2074),
    .C(n_5643),
    .Y(n_6667));
 OAI211xp5_ASAP7_75t_L g213742 (.A1(n_1669),
    .A2(n_4370),
    .B(n_6084),
    .C(n_5358),
    .Y(n_6666));
 AND5x1_ASAP7_75t_SL g213743 (.A(n_5298),
    .B(n_5269),
    .C(n_4680),
    .D(n_4194),
    .E(n_3360),
    .Y(n_6665));
 NOR5xp2_ASAP7_75t_L g213744 (.A(n_5254),
    .B(n_4095),
    .C(n_5355),
    .D(n_4530),
    .E(n_3452),
    .Y(n_6664));
 NAND2xp5_ASAP7_75t_R g213745 (.A(n_5519),
    .B(n_5809),
    .Y(n_6663));
 OA211x2_ASAP7_75t_SL g213746 (.A1(n_1418),
    .A2(n_1765),
    .B(n_1796),
    .C(n_5238),
    .Y(n_6662));
 A2O1A1Ixp33_ASAP7_75t_R g213747 (.A1(n_1683),
    .A2(n_3824),
    .B(n_4798),
    .C(n_2203),
    .Y(n_6661));
 NAND2xp33_ASAP7_75t_L g213748 (.A(n_6214),
    .B(n_5733),
    .Y(n_6660));
 NAND2xp33_ASAP7_75t_L g213749 (.A(n_5052),
    .B(n_5722),
    .Y(n_6659));
 NAND2xp5_ASAP7_75t_L g213750 (.A(n_5752),
    .B(n_6203),
    .Y(n_6658));
 NOR2xp33_ASAP7_75t_SL g213751 (.A(n_5051),
    .B(n_5762),
    .Y(n_6657));
 NAND2xp5_ASAP7_75t_L g213752 (.A(n_5493),
    .B(n_5804),
    .Y(n_6656));
 AOI211xp5_ASAP7_75t_L g213753 (.A1(n_4491),
    .A2(n_1500),
    .B(n_5488),
    .C(n_4766),
    .Y(n_6655));
 NAND2xp5_ASAP7_75t_L g213754 (.A(n_4213),
    .B(n_5720),
    .Y(n_6654));
 NOR5xp2_ASAP7_75t_SL g213755 (.A(n_5282),
    .B(n_4053),
    .C(n_4673),
    .D(n_5192),
    .E(n_3440),
    .Y(n_6653));
 OAI21xp33_ASAP7_75t_R g213756 (.A1(n_4895),
    .A2(n_4890),
    .B(n_3456),
    .Y(n_6652));
 NAND2xp33_ASAP7_75t_L g213757 (.A(n_4565),
    .B(n_5717),
    .Y(n_6651));
 AOI211xp5_ASAP7_75t_L g213758 (.A1(n_4196),
    .A2(n_1586),
    .B(n_4780),
    .C(n_1495),
    .Y(n_6650));
 O2A1O1Ixp33_ASAP7_75t_L g213759 (.A1(n_1669),
    .A2(n_3873),
    .B(n_4884),
    .C(n_1915),
    .Y(n_6649));
 A2O1A1Ixp33_ASAP7_75t_L g213760 (.A1(n_2192),
    .A2(n_1762),
    .B(n_4816),
    .C(sa00[0]),
    .Y(n_6648));
 NAND2xp33_ASAP7_75t_L g213761 (.A(n_5069),
    .B(n_5661),
    .Y(n_6647));
 AOI21xp5_ASAP7_75t_R g213762 (.A1(n_5468),
    .A2(n_4835),
    .B(n_1528),
    .Y(n_6646));
 NAND2xp5_ASAP7_75t_L g213763 (.A(n_5510),
    .B(n_6018),
    .Y(n_6645));
 OAI21xp33_ASAP7_75t_SL g213764 (.A1(n_4725),
    .A2(n_4874),
    .B(n_2684),
    .Y(n_6644));
 OAI221xp5_ASAP7_75t_L g213765 (.A1(n_5383),
    .A2(n_1376),
    .B1(n_4309),
    .B2(n_1544),
    .C(n_4863),
    .Y(n_6643));
 NAND2xp5_ASAP7_75t_L g213766 (.A(n_5508),
    .B(n_6057),
    .Y(n_6642));
 NOR2xp33_ASAP7_75t_SL g213767 (.A(n_5784),
    .B(n_6193),
    .Y(n_6641));
 A2O1A1Ixp33_ASAP7_75t_SL g213768 (.A1(sa03[3]),
    .A2(n_3811),
    .B(n_4808),
    .C(n_2601),
    .Y(n_6640));
 AOI211xp5_ASAP7_75t_L g213769 (.A1(n_3114),
    .A2(n_1683),
    .B(n_5041),
    .C(n_4627),
    .Y(n_6639));
 NAND2xp33_ASAP7_75t_L g213770 (.A(n_1797),
    .B(n_5773),
    .Y(n_6638));
 NAND2xp33_ASAP7_75t_L g213771 (.A(n_6197),
    .B(n_5766),
    .Y(n_6637));
 NOR2xp33_ASAP7_75t_L g213772 (.A(n_4960),
    .B(n_6189),
    .Y(n_6636));
 AOI221xp5_ASAP7_75t_SL g213773 (.A1(n_5535),
    .A2(n_2055),
    .B1(n_4449),
    .B2(n_1572),
    .C(n_5352),
    .Y(n_6635));
 AOI221xp5_ASAP7_75t_SL g213774 (.A1(n_3904),
    .A2(n_1391),
    .B1(n_5429),
    .B2(n_2042),
    .C(n_5367),
    .Y(n_6634));
 NAND2xp33_ASAP7_75t_R g213775 (.A(n_6216),
    .B(n_5679),
    .Y(n_6633));
 A2O1A1Ixp33_ASAP7_75t_SL g213776 (.A1(n_1343),
    .A2(n_3828),
    .B(n_4790),
    .C(n_3401),
    .Y(n_6632));
 NAND2xp33_ASAP7_75t_R g213777 (.A(n_4560),
    .B(n_5689),
    .Y(n_6631));
 NOR2xp33_ASAP7_75t_L g213778 (.A(n_3359),
    .B(n_6104),
    .Y(n_6630));
 OAI211xp5_ASAP7_75t_L g213779 (.A1(n_1678),
    .A2(n_3009),
    .B(n_5045),
    .C(n_4557),
    .Y(n_6629));
 OAI211xp5_ASAP7_75t_R g213780 (.A1(n_1679),
    .A2(n_3122),
    .B(n_5046),
    .C(n_4609),
    .Y(n_6628));
 OAI21xp33_ASAP7_75t_R g213781 (.A1(n_4769),
    .A2(n_5011),
    .B(n_1697),
    .Y(n_6627));
 OR3x1_ASAP7_75t_L g213782 (.A(n_4770),
    .B(n_4641),
    .C(n_2937),
    .Y(n_6626));
 NAND2xp5_ASAP7_75t_R g213783 (.A(n_5619),
    .B(n_1795),
    .Y(n_6625));
 NOR2xp33_ASAP7_75t_SL g213784 (.A(n_5665),
    .B(n_6224),
    .Y(n_6624));
 NAND2xp5_ASAP7_75t_L g213785 (.A(n_6164),
    .B(n_1795),
    .Y(n_6623));
 AOI21xp33_ASAP7_75t_R g213786 (.A1(n_4775),
    .A2(n_4991),
    .B(n_2541),
    .Y(n_6622));
 OAI21xp33_ASAP7_75t_R g213787 (.A1(n_2059),
    .A2(n_5534),
    .B(n_5651),
    .Y(n_6621));
 NOR2xp33_ASAP7_75t_L g213788 (.A(n_5642),
    .B(n_6196),
    .Y(n_6620));
 NAND2xp5_ASAP7_75t_L g213789 (.A(n_5646),
    .B(n_6230),
    .Y(n_6619));
 AOI211xp5_ASAP7_75t_L g213790 (.A1(n_4589),
    .A2(n_1585),
    .B(n_6193),
    .C(n_3784),
    .Y(n_6618));
 OR5x1_ASAP7_75t_SL g213791 (.A(n_3932),
    .B(n_1766),
    .C(n_4264),
    .D(n_4267),
    .E(n_3561),
    .Y(n_6617));
 OAI21xp33_ASAP7_75t_SL g213792 (.A1(n_1543),
    .A2(n_5430),
    .B(n_5713),
    .Y(n_6616));
 NAND2xp5_ASAP7_75t_L g213793 (.A(n_5755),
    .B(n_6187),
    .Y(n_6615));
 NOR2xp33_ASAP7_75t_SL g213794 (.A(n_5757),
    .B(n_6171),
    .Y(n_6614));
 AOI21xp33_ASAP7_75t_L g213795 (.A1(n_1643),
    .A2(n_5521),
    .B(n_5758),
    .Y(n_6613));
 A2O1A1Ixp33_ASAP7_75t_L g213796 (.A1(n_1411),
    .A2(n_4471),
    .B(n_4778),
    .C(n_1981),
    .Y(n_6612));
 NAND2xp5_ASAP7_75t_L g213797 (.A(n_4771),
    .B(n_6180),
    .Y(n_6611));
 A2O1A1Ixp33_ASAP7_75t_R g213798 (.A1(n_2756),
    .A2(n_4181),
    .B(n_2347),
    .C(n_5015),
    .Y(n_6610));
 NOR2xp33_ASAP7_75t_L g213799 (.A(n_4792),
    .B(n_6178),
    .Y(n_6609));
 AOI21xp33_ASAP7_75t_L g213800 (.A1(n_4862),
    .A2(n_2350),
    .B(n_5026),
    .Y(n_6608));
 A2O1A1Ixp33_ASAP7_75t_L g213801 (.A1(n_2754),
    .A2(n_4191),
    .B(n_2358),
    .C(n_5018),
    .Y(n_6607));
 NAND2xp5_ASAP7_75t_R g213802 (.A(n_4772),
    .B(n_6183),
    .Y(n_6606));
 NAND2xp5_ASAP7_75t_R g213803 (.A(n_6195),
    .B(n_5731),
    .Y(n_6605));
 A2O1A1Ixp33_ASAP7_75t_SL g213804 (.A1(n_2755),
    .A2(n_4094),
    .B(n_2365),
    .C(n_5016),
    .Y(n_6604));
 OAI211xp5_ASAP7_75t_L g213805 (.A1(n_4147),
    .A2(n_4285),
    .B(n_5512),
    .C(n_4715),
    .Y(n_6603));
 AOI211xp5_ASAP7_75t_L g213806 (.A1(n_2044),
    .A2(n_2592),
    .B(n_4757),
    .C(n_2937),
    .Y(n_6602));
 NAND2xp5_ASAP7_75t_R g213807 (.A(n_5823),
    .B(n_6208),
    .Y(n_6601));
 OA211x2_ASAP7_75t_SL g213808 (.A1(n_2047),
    .A2(n_4332),
    .B(n_5463),
    .C(n_4719),
    .Y(n_6600));
 A2O1A1Ixp33_ASAP7_75t_SL g213809 (.A1(n_2059),
    .A2(n_4354),
    .B(n_5222),
    .C(n_5263),
    .Y(n_6599));
 O2A1O1Ixp33_ASAP7_75t_SL g213810 (.A1(n_2413),
    .A2(n_4355),
    .B(n_5195),
    .C(n_5270),
    .Y(n_6598));
 A2O1A1Ixp33_ASAP7_75t_L g213811 (.A1(n_1548),
    .A2(n_4360),
    .B(n_5218),
    .C(n_5279),
    .Y(n_6597));
 A2O1A1Ixp33_ASAP7_75t_SL g213812 (.A1(n_2057),
    .A2(n_3863),
    .B(n_5217),
    .C(n_5274),
    .Y(n_6596));
 A2O1A1Ixp33_ASAP7_75t_SL g213813 (.A1(n_2045),
    .A2(n_3880),
    .B(n_5213),
    .C(n_5285),
    .Y(n_6595));
 O2A1O1Ixp33_ASAP7_75t_L g213814 (.A1(n_2404),
    .A2(n_3885),
    .B(n_5181),
    .C(n_5297),
    .Y(n_6594));
 A2O1A1Ixp33_ASAP7_75t_SL g213815 (.A1(n_2043),
    .A2(n_3897),
    .B(n_5211),
    .C(n_5281),
    .Y(n_6593));
 OAI211xp5_ASAP7_75t_L g213816 (.A1(n_3861),
    .A2(n_4270),
    .B(n_5721),
    .C(n_2646),
    .Y(n_6592));
 A2O1A1Ixp33_ASAP7_75t_L g213817 (.A1(n_1934),
    .A2(n_4403),
    .B(n_5208),
    .C(n_2220),
    .Y(n_6591));
 AOI221xp5_ASAP7_75t_SL g213818 (.A1(n_3727),
    .A2(n_1566),
    .B1(n_1559),
    .B2(n_2530),
    .C(n_5805),
    .Y(n_6590));
 AOI211xp5_ASAP7_75t_L g213819 (.A1(n_4013),
    .A2(n_1673),
    .B(n_5227),
    .C(n_4803),
    .Y(n_6589));
 A2O1A1Ixp33_ASAP7_75t_SL g213820 (.A1(sa22[3]),
    .A2(n_2781),
    .B(n_4813),
    .C(n_2671),
    .Y(n_6588));
 AOI211xp5_ASAP7_75t_SL g213821 (.A1(n_4011),
    .A2(n_2471),
    .B(n_5231),
    .C(n_4805),
    .Y(n_6587));
 A2O1A1Ixp33_ASAP7_75t_SL g213822 (.A1(n_1343),
    .A2(n_2784),
    .B(n_4815),
    .C(n_2684),
    .Y(n_6586));
 NAND2xp33_ASAP7_75t_SL g213823 (.A(n_4812),
    .B(n_5786),
    .Y(n_6585));
 O2A1O1Ixp33_ASAP7_75t_L g213824 (.A1(n_1859),
    .A2(n_4044),
    .B(n_4810),
    .C(n_3398),
    .Y(n_6584));
 AOI211xp5_ASAP7_75t_SL g213825 (.A1(n_1549),
    .A2(n_2506),
    .B(n_5781),
    .C(n_5256),
    .Y(n_6583));
 AOI211xp5_ASAP7_75t_SL g213826 (.A1(n_4488),
    .A2(n_2413),
    .B(n_5409),
    .C(n_3744),
    .Y(n_6582));
 OAI211xp5_ASAP7_75t_SL g213827 (.A1(n_1568),
    .A2(n_4436),
    .B(n_5421),
    .C(n_3747),
    .Y(n_6581));
 OAI211xp5_ASAP7_75t_SL g213828 (.A1(n_1632),
    .A2(n_4478),
    .B(n_5439),
    .C(n_3745),
    .Y(n_6580));
 OAI211xp5_ASAP7_75t_SL g213829 (.A1(n_2422),
    .A2(n_4466),
    .B(n_5427),
    .C(n_3741),
    .Y(n_6579));
 OAI211xp5_ASAP7_75t_L g213830 (.A1(n_1383),
    .A2(n_4393),
    .B(n_5424),
    .C(n_3742),
    .Y(n_6578));
 NOR3xp33_ASAP7_75t_SL g213831 (.A(n_5899),
    .B(n_4949),
    .C(n_1510),
    .Y(n_6577));
 NAND2xp33_ASAP7_75t_SL g213832 (.A(n_5451),
    .B(n_6134),
    .Y(n_6576));
 OAI211xp5_ASAP7_75t_SL g213833 (.A1(n_1458),
    .A2(n_4821),
    .B(n_5224),
    .C(n_3439),
    .Y(n_6575));
 OAI221xp5_ASAP7_75t_L g213834 (.A1(n_5388),
    .A2(n_4981),
    .B1(n_4476),
    .B2(n_1632),
    .C(n_2646),
    .Y(n_6574));
 A2O1A1Ixp33_ASAP7_75t_R g213835 (.A1(n_1458),
    .A2(n_4381),
    .B(n_5371),
    .C(n_2180),
    .Y(n_6573));
 AOI211xp5_ASAP7_75t_L g213836 (.A1(n_3571),
    .A2(n_2103),
    .B(n_5280),
    .C(n_3923),
    .Y(n_6572));
 O2A1O1Ixp33_ASAP7_75t_SL g213837 (.A1(n_8210),
    .A2(n_4218),
    .B(n_4795),
    .C(n_2595),
    .Y(n_6571));
 O2A1O1Ixp33_ASAP7_75t_L g213838 (.A1(n_1518),
    .A2(n_4589),
    .B(n_4787),
    .C(n_2565),
    .Y(n_6570));
 AOI221xp5_ASAP7_75t_L g213839 (.A1(n_3087),
    .A2(n_2023),
    .B1(n_2952),
    .B2(n_1439),
    .C(n_4867),
    .Y(n_6569));
 OAI221xp5_ASAP7_75t_SL g213840 (.A1(n_5264),
    .A2(n_1656),
    .B1(n_4129),
    .B2(n_2844),
    .C(n_5315),
    .Y(n_6568));
 OAI221xp5_ASAP7_75t_R g213841 (.A1(n_2424),
    .A2(n_2922),
    .B1(n_1544),
    .B2(n_1522),
    .C(n_6071),
    .Y(n_6567));
 OAI221xp5_ASAP7_75t_L g213842 (.A1(n_5302),
    .A2(n_2057),
    .B1(n_4117),
    .B2(n_1590),
    .C(n_4806),
    .Y(n_6566));
 AOI21xp33_ASAP7_75t_L g213843 (.A1(n_5410),
    .A2(n_4870),
    .B(sa12[0]),
    .Y(n_6565));
 AOI21xp33_ASAP7_75t_L g213844 (.A1(n_5399),
    .A2(n_4985),
    .B(n_6061),
    .Y(n_6564));
 OAI221xp5_ASAP7_75t_R g213845 (.A1(n_3060),
    .A2(n_3492),
    .B1(n_1769),
    .B2(n_1674),
    .C(n_5694),
    .Y(n_6563));
 AOI211xp5_ASAP7_75t_SL g213846 (.A1(n_3893),
    .A2(n_1559),
    .B(n_5725),
    .C(n_5183),
    .Y(n_6562));
 NOR3xp33_ASAP7_75t_L g213847 (.A(n_6079),
    .B(n_4575),
    .C(n_3934),
    .Y(n_6561));
 OAI211xp5_ASAP7_75t_L g213848 (.A1(n_1933),
    .A2(n_4477),
    .B(n_5232),
    .C(n_3572),
    .Y(n_6560));
 OAI211xp5_ASAP7_75t_L g213849 (.A1(n_1850),
    .A2(n_4046),
    .B(n_5234),
    .C(n_3551),
    .Y(n_6559));
 OAI211xp5_ASAP7_75t_SL g213850 (.A1(n_1632),
    .A2(n_4082),
    .B(n_4796),
    .C(n_4210),
    .Y(n_6558));
 OAI211xp5_ASAP7_75t_SL g213851 (.A1(n_5004),
    .A2(n_5351),
    .B(n_4897),
    .C(n_2673),
    .Y(n_6557));
 A2O1A1Ixp33_ASAP7_75t_SL g213852 (.A1(n_2473),
    .A2(n_4287),
    .B(n_2070),
    .C(n_5832),
    .Y(n_6556));
 OAI211xp5_ASAP7_75t_SL g213853 (.A1(n_1544),
    .A2(n_4252),
    .B(n_5498),
    .C(n_6115),
    .Y(n_6555));
 OAI211xp5_ASAP7_75t_L g213854 (.A1(n_1568),
    .A2(n_4103),
    .B(n_4788),
    .C(n_4161),
    .Y(n_6554));
 A2O1A1Ixp33_ASAP7_75t_L g213855 (.A1(n_1984),
    .A2(n_4576),
    .B(n_4801),
    .C(n_2615),
    .Y(n_6553));
 A2O1A1Ixp33_ASAP7_75t_SL g213856 (.A1(n_1680),
    .A2(n_4216),
    .B(n_2061),
    .C(n_5853),
    .Y(n_6552));
 AOI211xp5_ASAP7_75t_R g213857 (.A1(n_5336),
    .A2(n_4999),
    .B(n_4872),
    .C(n_2672),
    .Y(n_6551));
 OAI311xp33_ASAP7_75t_SL g213858 (.A1(n_3285),
    .A2(n_3313),
    .A3(n_2430),
    .B1(n_4155),
    .C1(n_4784),
    .Y(n_6550));
 A2O1A1Ixp33_ASAP7_75t_L g213859 (.A1(n_2471),
    .A2(n_4219),
    .B(n_1450),
    .C(n_5848),
    .Y(n_6549));
 NAND2xp5_ASAP7_75t_SL g213860 (.A(n_5984),
    .B(n_5702),
    .Y(n_6548));
 AOI221xp5_ASAP7_75t_SL g213861 (.A1(n_4205),
    .A2(n_2069),
    .B1(n_2804),
    .B2(n_2044),
    .C(n_5523),
    .Y(n_6547));
 AOI211xp5_ASAP7_75t_SL g213862 (.A1(n_3985),
    .A2(n_1432),
    .B(n_5290),
    .C(n_5452),
    .Y(n_6546));
 OAI211xp5_ASAP7_75t_L g213863 (.A1(n_1651),
    .A2(n_4141),
    .B(n_6068),
    .C(n_2679),
    .Y(n_6545));
 OAI211xp5_ASAP7_75t_L g213864 (.A1(n_2447),
    .A2(n_3135),
    .B(n_5366),
    .C(n_4520),
    .Y(n_6544));
 O2A1O1Ixp33_ASAP7_75t_SL g213865 (.A1(n_1975),
    .A2(n_3857),
    .B(n_4989),
    .C(n_6083),
    .Y(n_6543));
 O2A1O1Ixp33_ASAP7_75t_R g213866 (.A1(n_1671),
    .A2(n_4382),
    .B(n_1435),
    .C(n_5847),
    .Y(n_6542));
 AOI211xp5_ASAP7_75t_SL g213867 (.A1(n_3944),
    .A2(n_1657),
    .B(n_5319),
    .C(n_5485),
    .Y(n_6541));
 OAI221xp5_ASAP7_75t_L g213868 (.A1(n_5268),
    .A2(n_1417),
    .B1(n_4146),
    .B2(n_1571),
    .C(n_4786),
    .Y(n_6540));
 NOR3xp33_ASAP7_75t_L g213869 (.A(n_5128),
    .B(n_5074),
    .C(n_2672),
    .Y(n_6539));
 OAI221xp5_ASAP7_75t_L g213870 (.A1(n_5286),
    .A2(n_1544),
    .B1(n_4136),
    .B2(n_2073),
    .C(n_4774),
    .Y(n_6538));
 OAI211xp5_ASAP7_75t_L g213871 (.A1(n_1383),
    .A2(n_4048),
    .B(n_5506),
    .C(n_5322),
    .Y(n_6537));
 OAI211xp5_ASAP7_75t_L g213872 (.A1(n_2412),
    .A2(n_4040),
    .B(n_5481),
    .C(n_5337),
    .Y(n_6536));
 OAI321xp33_ASAP7_75t_L g213873 (.A1(n_4290),
    .A2(n_1590),
    .A3(n_2606),
    .B1(n_2057),
    .B2(n_3872),
    .C(n_5555),
    .Y(n_6535));
 OAI211xp5_ASAP7_75t_L g213874 (.A1(n_2422),
    .A2(n_3962),
    .B(n_5494),
    .C(n_5233),
    .Y(n_6534));
 AOI22xp33_ASAP7_75t_L g213875 (.A1(n_4982),
    .A2(n_5387),
    .B1(n_1406),
    .B2(n_3803),
    .Y(n_6533));
 OAI211xp5_ASAP7_75t_R g213876 (.A1(n_1407),
    .A2(n_3965),
    .B(n_5482),
    .C(n_5340),
    .Y(n_6532));
 OAI211xp5_ASAP7_75t_SL g213877 (.A1(n_1656),
    .A2(n_4047),
    .B(n_6074),
    .C(n_2670),
    .Y(n_6531));
 AOI322xp5_ASAP7_75t_SL g213878 (.A1(n_4651),
    .A2(n_2064),
    .A3(n_1603),
    .B1(n_8703),
    .B2(n_4500),
    .C1(n_3788),
    .C2(n_4301),
    .Y(n_6530));
 O2A1O1Ixp33_ASAP7_75t_SL g213879 (.A1(n_2492),
    .A2(n_4402),
    .B(n_1440),
    .C(n_5840),
    .Y(n_6529));
 AOI21xp5_ASAP7_75t_R g213880 (.A1(n_4303),
    .A2(n_2392),
    .B(n_6206),
    .Y(n_6528));
 AOI21xp5_ASAP7_75t_L g213881 (.A1(n_4282),
    .A2(n_2400),
    .B(n_6204),
    .Y(n_6527));
 A2O1A1Ixp33_ASAP7_75t_R g213882 (.A1(n_1595),
    .A2(n_3918),
    .B(n_4750),
    .C(n_1510),
    .Y(n_6526));
 AOI211xp5_ASAP7_75t_SL g213883 (.A1(n_4072),
    .A2(n_1465),
    .B(n_4730),
    .C(n_3843),
    .Y(n_6525));
 A2O1A1Ixp33_ASAP7_75t_L g213884 (.A1(n_2483),
    .A2(n_4298),
    .B(n_1578),
    .C(n_5837),
    .Y(n_6524));
 AO21x1_ASAP7_75t_SL g213885 (.A1(n_8703),
    .A2(n_5462),
    .B(sa12[2]),
    .Y(n_6523));
 A2O1A1Ixp33_ASAP7_75t_SL g213886 (.A1(n_2477),
    .A2(n_4286),
    .B(n_1381),
    .C(n_5834),
    .Y(n_6522));
 NOR4xp25_ASAP7_75t_L g213887 (.A(n_3955),
    .B(n_4182),
    .C(n_5299),
    .D(n_3921),
    .Y(n_6521));
 AOI21xp5_ASAP7_75t_SL g213888 (.A1(n_5378),
    .A2(n_1400),
    .B(n_5771),
    .Y(n_6520));
 AOI221xp5_ASAP7_75t_L g213889 (.A1(n_3815),
    .A2(n_4064),
    .B1(n_3817),
    .B2(n_1581),
    .C(sa33[0]),
    .Y(n_6519));
 OAI211xp5_ASAP7_75t_L g213890 (.A1(n_1634),
    .A2(n_3950),
    .B(n_5313),
    .C(n_5475),
    .Y(n_6518));
 A2O1A1Ixp33_ASAP7_75t_SL g213891 (.A1(n_2485),
    .A2(n_1777),
    .B(n_2083),
    .C(n_5829),
    .Y(n_6517));
 O2A1O1Ixp33_ASAP7_75t_L g213892 (.A1(n_2476),
    .A2(n_3846),
    .B(n_1401),
    .C(n_5838),
    .Y(n_6516));
 AOI222xp33_ASAP7_75t_L g213893 (.A1(n_4403),
    .A2(n_1436),
    .B1(n_3215),
    .B2(n_2450),
    .C1(n_4833),
    .C2(n_1404),
    .Y(n_6515));
 NAND3xp33_ASAP7_75t_L g213894 (.A(n_4819),
    .B(n_4745),
    .C(n_2957),
    .Y(n_6514));
 OAI21xp33_ASAP7_75t_L g213895 (.A1(n_2428),
    .A2(n_5392),
    .B(n_5765),
    .Y(n_6513));
 AO21x1_ASAP7_75t_L g213896 (.A1(n_1655),
    .A2(n_3876),
    .B(n_5620),
    .Y(n_6512));
 OAI211xp5_ASAP7_75t_L g213897 (.A1(n_1344),
    .A2(n_4287),
    .B(n_5441),
    .C(n_2670),
    .Y(n_6511));
 AOI211xp5_ASAP7_75t_L g213898 (.A1(n_3853),
    .A2(n_1412),
    .B(n_5578),
    .C(n_5420),
    .Y(n_6510));
 OAI221xp5_ASAP7_75t_SL g213899 (.A1(n_3045),
    .A2(n_1522),
    .B1(n_2424),
    .B2(n_3064),
    .C(n_4820),
    .Y(n_6509));
 AOI221xp5_ASAP7_75t_SL g213900 (.A1(n_4383),
    .A2(n_1545),
    .B1(n_5383),
    .B2(n_1446),
    .C(n_5328),
    .Y(n_6508));
 OAI221xp5_ASAP7_75t_SL g213901 (.A1(n_4003),
    .A2(n_1501),
    .B1(n_1629),
    .B2(n_2574),
    .C(n_6009),
    .Y(n_6507));
 O2A1O1Ixp33_ASAP7_75t_L g213902 (.A1(n_2468),
    .A2(n_4327),
    .B(n_1570),
    .C(n_5831),
    .Y(n_6506));
 AOI221xp5_ASAP7_75t_R g213903 (.A1(n_4676),
    .A2(n_1643),
    .B1(n_2889),
    .B2(n_1397),
    .C(n_4746),
    .Y(n_6505));
 OAI221xp5_ASAP7_75t_L g213904 (.A1(n_3987),
    .A2(sa11[6]),
    .B1(n_1450),
    .B2(n_2519),
    .C(n_5237),
    .Y(n_6504));
 AOI221xp5_ASAP7_75t_R g213905 (.A1(n_4063),
    .A2(n_1410),
    .B1(n_1451),
    .B2(n_2570),
    .C(n_5995),
    .Y(n_6503));
 AOI221xp5_ASAP7_75t_SL g213906 (.A1(n_3073),
    .A2(n_1754),
    .B1(n_2984),
    .B2(n_2282),
    .C(n_5774),
    .Y(n_6502));
 AOI221xp5_ASAP7_75t_L g213907 (.A1(n_2978),
    .A2(n_1982),
    .B1(n_3040),
    .B2(n_1405),
    .C(n_4824),
    .Y(n_6501));
 AOI211xp5_ASAP7_75t_L g213908 (.A1(n_3517),
    .A2(sa21[3]),
    .B(n_5704),
    .C(n_3467),
    .Y(n_6500));
 OAI22xp33_ASAP7_75t_R g213909 (.A1(n_4986),
    .A2(n_5397),
    .B1(n_2423),
    .B2(n_4403),
    .Y(n_6499));
 A2O1A1Ixp33_ASAP7_75t_SL g213910 (.A1(n_2448),
    .A2(n_4326),
    .B(n_2091),
    .C(n_5798),
    .Y(n_6498));
 AOI222xp33_ASAP7_75t_SL g213911 (.A1(n_4856),
    .A2(n_1938),
    .B1(n_4100),
    .B2(n_1748),
    .C1(n_2991),
    .C2(n_2079),
    .Y(n_6497));
 A2O1A1Ixp33_ASAP7_75t_R g213912 (.A1(n_1496),
    .A2(n_3996),
    .B(n_1438),
    .C(n_4331),
    .Y(n_6496));
 OAI211xp5_ASAP7_75t_L g213913 (.A1(n_1669),
    .A2(n_4043),
    .B(n_6125),
    .C(n_2666),
    .Y(n_6495));
 AOI211xp5_ASAP7_75t_L g213914 (.A1(n_4058),
    .A2(n_1401),
    .B(n_5499),
    .C(n_4975),
    .Y(n_6494));
 AOI211xp5_ASAP7_75t_L g213915 (.A1(n_2795),
    .A2(n_2055),
    .B(n_5572),
    .C(n_5415),
    .Y(n_6493));
 A2O1A1Ixp33_ASAP7_75t_L g213916 (.A1(n_2442),
    .A2(n_4314),
    .B(n_1590),
    .C(n_5779),
    .Y(n_6492));
 O2A1O1Ixp33_ASAP7_75t_L g213917 (.A1(n_2441),
    .A2(n_1776),
    .B(n_1424),
    .C(n_5796),
    .Y(n_6491));
 AOI221xp5_ASAP7_75t_L g213918 (.A1(n_3737),
    .A2(n_1349),
    .B1(n_5296),
    .B2(n_4983),
    .C(n_2683),
    .Y(n_6490));
 AOI221xp5_ASAP7_75t_L g213919 (.A1(n_3879),
    .A2(n_2062),
    .B1(n_4523),
    .B2(n_2416),
    .C(n_3769),
    .Y(n_6489));
 OAI211xp5_ASAP7_75t_SL g213920 (.A1(n_2591),
    .A2(n_4010),
    .B(n_5486),
    .C(n_4896),
    .Y(n_6488));
 OAI211xp5_ASAP7_75t_L g213921 (.A1(n_1676),
    .A2(n_3069),
    .B(n_4875),
    .C(n_4214),
    .Y(n_6487));
 OAI221xp5_ASAP7_75t_R g213922 (.A1(n_4168),
    .A2(n_1744),
    .B1(n_2961),
    .B2(n_2099),
    .C(n_5986),
    .Y(n_6486));
 OAI22xp33_ASAP7_75t_L g213923 (.A1(n_4727),
    .A2(n_1465),
    .B1(n_5363),
    .B2(n_1464),
    .Y(n_6485));
 OAI221xp5_ASAP7_75t_L g213924 (.A1(n_4404),
    .A2(n_2415),
    .B1(n_4016),
    .B2(n_2570),
    .C(n_4898),
    .Y(n_6484));
 OAI221xp5_ASAP7_75t_L g213925 (.A1(n_4167),
    .A2(n_2091),
    .B1(n_1730),
    .B2(n_1560),
    .C(n_5434),
    .Y(n_6483));
 AOI222xp33_ASAP7_75t_SL g213926 (.A1(n_4836),
    .A2(n_1501),
    .B1(n_4463),
    .B2(n_1350),
    .C1(n_3097),
    .C2(n_1401),
    .Y(n_6482));
 AOI211xp5_ASAP7_75t_L g213927 (.A1(n_3734),
    .A2(n_1633),
    .B(n_4759),
    .C(n_2398),
    .Y(n_6481));
 AOI22xp5_ASAP7_75t_SL g213928 (.A1(n_1499),
    .A2(n_4722),
    .B1(n_1498),
    .B2(n_5362),
    .Y(n_6480));
 AOI211xp5_ASAP7_75t_SL g213929 (.A1(n_4005),
    .A2(n_2589),
    .B(n_4904),
    .C(n_5483),
    .Y(n_6479));
 AOI22xp5_ASAP7_75t_SL g213930 (.A1(n_1496),
    .A2(n_4720),
    .B1(n_1497),
    .B2(n_5361),
    .Y(n_6478));
 AOI221xp5_ASAP7_75t_SL g213931 (.A1(n_4839),
    .A2(n_1499),
    .B1(n_2732),
    .B2(n_2090),
    .C(n_5204),
    .Y(n_6477));
 OAI211xp5_ASAP7_75t_L g213932 (.A1(n_1346),
    .A2(n_2899),
    .B(n_4718),
    .C(n_5191),
    .Y(n_6476));
 OAI31xp33_ASAP7_75t_R g213933 (.A1(n_4768),
    .A2(n_4086),
    .A3(n_4548),
    .B(n_2267),
    .Y(n_6475));
 OAI221xp5_ASAP7_75t_L g213934 (.A1(n_4502),
    .A2(n_4439),
    .B1(n_4497),
    .B2(n_2445),
    .C(n_5673),
    .Y(n_6474));
 AOI31xp33_ASAP7_75t_R g213935 (.A1(n_4749),
    .A2(n_4528),
    .A3(n_4074),
    .B(n_2244),
    .Y(n_6473));
 OAI221xp5_ASAP7_75t_R g213936 (.A1(n_4030),
    .A2(n_1573),
    .B1(n_2779),
    .B2(n_1417),
    .C(n_5407),
    .Y(n_6472));
 AOI21xp5_ASAP7_75t_SL g213937 (.A1(n_4188),
    .A2(n_1431),
    .B(n_6046),
    .Y(n_6471));
 OAI221xp5_ASAP7_75t_SL g213938 (.A1(n_4375),
    .A2(n_1442),
    .B1(n_4009),
    .B2(n_2548),
    .C(n_4881),
    .Y(n_6470));
 OAI211xp5_ASAP7_75t_L g213939 (.A1(n_2546),
    .A2(n_4014),
    .B(n_5489),
    .C(n_4878),
    .Y(n_6469));
 OAI211xp5_ASAP7_75t_L g213940 (.A1(n_2550),
    .A2(n_1769),
    .B(n_5494),
    .C(n_4883),
    .Y(n_6468));
 AOI21xp5_ASAP7_75t_L g213941 (.A1(n_5384),
    .A2(n_1664),
    .B(n_5628),
    .Y(n_6467));
 NAND2xp5_ASAP7_75t_L g213942 (.A(n_5481),
    .B(n_6158),
    .Y(n_6466));
 OAI221xp5_ASAP7_75t_SL g213943 (.A1(n_4110),
    .A2(n_1716),
    .B1(n_2987),
    .B2(n_1342),
    .C(n_5956),
    .Y(n_6465));
 NAND4xp25_ASAP7_75t_L g213944 (.A(n_4663),
    .B(n_4854),
    .C(n_3220),
    .D(n_3183),
    .Y(n_6464));
 OAI211xp5_ASAP7_75t_SL g213945 (.A1(n_2059),
    .A2(n_4303),
    .B(n_5517),
    .C(n_4714),
    .Y(n_6463));
 OAI211xp5_ASAP7_75t_SL g213946 (.A1(n_1938),
    .A2(n_4069),
    .B(n_4751),
    .C(n_3800),
    .Y(n_6462));
 OAI211xp5_ASAP7_75t_SL g213947 (.A1(n_1933),
    .A2(n_3994),
    .B(n_4753),
    .C(n_3799),
    .Y(n_6461));
 AOI221xp5_ASAP7_75t_SL g213948 (.A1(n_1762),
    .A2(n_2241),
    .B1(n_4363),
    .B2(n_1570),
    .C(n_5248),
    .Y(n_6460));
 OAI221xp5_ASAP7_75t_L g213949 (.A1(n_1571),
    .A2(n_2795),
    .B1(n_1417),
    .B2(n_8200),
    .C(n_5547),
    .Y(n_6459));
 OAI21xp33_ASAP7_75t_SL g213950 (.A1(n_2053),
    .A2(n_4195),
    .B(n_6031),
    .Y(n_6458));
 OAI221xp5_ASAP7_75t_SL g213951 (.A1(n_2948),
    .A2(n_2015),
    .B1(n_3025),
    .B2(n_1450),
    .C(n_4710),
    .Y(n_6457));
 OAI211xp5_ASAP7_75t_SL g213952 (.A1(n_1496),
    .A2(n_3998),
    .B(n_4755),
    .C(n_3798),
    .Y(n_6456));
 A2O1A1Ixp33_ASAP7_75t_SL g213953 (.A1(n_2820),
    .A2(n_4286),
    .B(n_1623),
    .C(n_5639),
    .Y(n_6455));
 OAI221xp5_ASAP7_75t_SL g213954 (.A1(n_4113),
    .A2(n_1381),
    .B1(n_2777),
    .B2(n_2043),
    .C(n_5120),
    .Y(n_6454));
 AOI211xp5_ASAP7_75t_SL g213955 (.A1(n_2933),
    .A2(n_2490),
    .B(n_1762),
    .C(n_5952),
    .Y(n_6453));
 OAI311xp33_ASAP7_75t_R g213956 (.A1(n_3320),
    .A2(n_2074),
    .A3(n_3433),
    .B1(n_1740),
    .C1(n_4726),
    .Y(n_6452));
 NAND2xp5_ASAP7_75t_L g213957 (.A(n_6213),
    .B(n_5877),
    .Y(n_6451));
 OAI322xp33_ASAP7_75t_R g213958 (.A1(n_1355),
    .A2(n_2832),
    .A3(n_2573),
    .B1(n_4349),
    .B2(n_1541),
    .C1(n_4262),
    .C2(n_1628),
    .Y(n_6449));
 AOI221xp5_ASAP7_75t_SL g213959 (.A1(n_4169),
    .A2(n_8703),
    .B1(n_2064),
    .B2(n_3274),
    .C(n_5645),
    .Y(n_6448));
 OAI221xp5_ASAP7_75t_L g213960 (.A1(n_4062),
    .A2(n_1363),
    .B1(n_3260),
    .B2(n_1551),
    .C(n_5531),
    .Y(n_6447));
 AOI221xp5_ASAP7_75t_SL g213961 (.A1(n_4474),
    .A2(n_4597),
    .B1(n_4442),
    .B2(n_2494),
    .C(n_5674),
    .Y(n_6446));
 AOI222xp33_ASAP7_75t_L g213962 (.A1(n_4832),
    .A2(n_1459),
    .B1(n_4381),
    .B2(n_1421),
    .C1(n_3163),
    .C2(n_1423),
    .Y(n_6445));
 OAI211xp5_ASAP7_75t_SL g213963 (.A1(n_4125),
    .A2(n_1404),
    .B(n_4756),
    .C(n_3801),
    .Y(n_6444));
 OAI211xp5_ASAP7_75t_L g213964 (.A1(n_3288),
    .A2(n_3129),
    .B(n_4885),
    .C(n_5496),
    .Y(n_6443));
 A2O1A1Ixp33_ASAP7_75t_R g213965 (.A1(n_2819),
    .A2(n_4298),
    .B(n_1647),
    .C(n_5609),
    .Y(n_6442));
 OAI211xp5_ASAP7_75t_L g213966 (.A1(n_1568),
    .A2(n_4122),
    .B(n_4748),
    .C(n_1565),
    .Y(n_6441));
 AOI211xp5_ASAP7_75t_R g213967 (.A1(n_4003),
    .A2(n_1446),
    .B(n_5997),
    .C(n_3785),
    .Y(n_6440));
 AOI211xp5_ASAP7_75t_L g213968 (.A1(n_4114),
    .A2(n_1458),
    .B(n_4760),
    .C(n_3809),
    .Y(n_6439));
 OAI311xp33_ASAP7_75t_L g213969 (.A1(n_3421),
    .A2(n_3386),
    .A3(n_2091),
    .B1(n_3358),
    .C1(n_4728),
    .Y(n_6438));
 OAI221xp5_ASAP7_75t_L g213970 (.A1(n_3997),
    .A2(n_1565),
    .B1(n_3145),
    .B2(n_1562),
    .C(n_5573),
    .Y(n_6437));
 OAI211xp5_ASAP7_75t_L g213971 (.A1(n_1456),
    .A2(n_3957),
    .B(n_4758),
    .C(n_3802),
    .Y(n_6436));
 A2O1A1Ixp33_ASAP7_75t_SL g213972 (.A1(n_1671),
    .A2(n_1623),
    .B(n_5043),
    .C(n_5372),
    .Y(n_6435));
 OAI211xp5_ASAP7_75t_L g213973 (.A1(n_2081),
    .A2(n_1761),
    .B(n_5585),
    .C(n_5073),
    .Y(n_6434));
 OAI221xp5_ASAP7_75t_SL g213974 (.A1(n_3866),
    .A2(n_1373),
    .B1(n_1763),
    .B2(n_2047),
    .C(n_5543),
    .Y(n_6433));
 OAI221xp5_ASAP7_75t_L g213975 (.A1(n_4102),
    .A2(n_2428),
    .B1(n_3547),
    .B2(n_2501),
    .C(n_4913),
    .Y(n_6432));
 OAI221xp5_ASAP7_75t_SL g213976 (.A1(n_1790),
    .A2(n_1651),
    .B1(n_4124),
    .B2(n_3290),
    .C(n_5020),
    .Y(n_6431));
 OAI211xp5_ASAP7_75t_SL g213977 (.A1(n_1541),
    .A2(n_2817),
    .B(n_5965),
    .C(n_4154),
    .Y(n_6430));
 AOI221xp5_ASAP7_75t_SL g213978 (.A1(n_3972),
    .A2(n_3297),
    .B1(n_3037),
    .B2(n_1982),
    .C(n_4880),
    .Y(n_6429));
 NOR2xp33_ASAP7_75t_SL g213979 (.A(n_5207),
    .B(n_5636),
    .Y(n_6428));
 OAI221xp5_ASAP7_75t_SL g213980 (.A1(n_4508),
    .A2(n_2066),
    .B1(n_2444),
    .B2(n_2088),
    .C(n_6064),
    .Y(n_6427));
 NOR3xp33_ASAP7_75t_SL g213981 (.A(n_5488),
    .B(n_5442),
    .C(n_2667),
    .Y(n_6426));
 OAI211xp5_ASAP7_75t_SL g213982 (.A1(n_3290),
    .A2(n_3089),
    .B(n_5594),
    .C(n_5438),
    .Y(n_6425));
 OAI221xp5_ASAP7_75t_L g213983 (.A1(n_4189),
    .A2(n_1584),
    .B1(n_3258),
    .B2(n_2059),
    .C(n_5522),
    .Y(n_6424));
 OAI221xp5_ASAP7_75t_L g213984 (.A1(n_4494),
    .A2(n_1624),
    .B1(n_2078),
    .B2(n_1673),
    .C(n_6013),
    .Y(n_6423));
 AOI211xp5_ASAP7_75t_L g213985 (.A1(n_1416),
    .A2(n_2316),
    .B(n_6025),
    .C(n_4626),
    .Y(n_6422));
 AOI221xp5_ASAP7_75t_L g213986 (.A1(n_4419),
    .A2(n_4452),
    .B1(n_4486),
    .B2(n_2471),
    .C(n_5611),
    .Y(n_6421));
 AOI322xp5_ASAP7_75t_L g213987 (.A1(n_2813),
    .A2(n_1667),
    .A3(n_2328),
    .B1(n_1447),
    .B2(n_3856),
    .C1(n_4892),
    .C2(n_1465),
    .Y(n_6420));
 OAI211xp5_ASAP7_75t_L g213988 (.A1(n_2068),
    .A2(n_4282),
    .B(n_5515),
    .C(n_4871),
    .Y(n_6419));
 AOI221xp5_ASAP7_75t_SL g213989 (.A1(n_4458),
    .A2(n_1405),
    .B1(n_1423),
    .B2(n_2465),
    .C(n_5960),
    .Y(n_6418));
 NAND3xp33_ASAP7_75t_L g213990 (.A(n_5616),
    .B(n_5348),
    .C(n_1495),
    .Y(n_6417));
 AOI211xp5_ASAP7_75t_L g213991 (.A1(n_1765),
    .A2(n_2414),
    .B(n_5622),
    .C(n_8199),
    .Y(n_6416));
 OAI322xp33_ASAP7_75t_SL g213992 (.A1(n_3252),
    .A2(n_1442),
    .A3(n_3342),
    .B1(n_5139),
    .B2(n_1395),
    .C1(n_3103),
    .C2(n_2081),
    .Y(n_6415));
 OAI221xp5_ASAP7_75t_SL g213993 (.A1(n_3965),
    .A2(n_1654),
    .B1(n_1756),
    .B2(n_1571),
    .C(n_5974),
    .Y(n_6414));
 O2A1O1Ixp33_ASAP7_75t_SL g213994 (.A1(sa30[3]),
    .A2(n_3197),
    .B(n_5533),
    .C(n_3804),
    .Y(n_6413));
 OAI211xp5_ASAP7_75t_L g213995 (.A1(n_2388),
    .A2(n_4667),
    .B(n_4717),
    .C(n_4848),
    .Y(n_6412));
 AOI221xp5_ASAP7_75t_L g213996 (.A1(n_4973),
    .A2(n_1737),
    .B1(n_1783),
    .B2(n_3127),
    .C(n_5310),
    .Y(n_6411));
 AND4x1_ASAP7_75t_SL g213997 (.A(n_5444),
    .B(n_4902),
    .C(n_3193),
    .D(n_1870),
    .Y(n_6410));
 AOI321xp33_ASAP7_75t_SL g213998 (.A1(n_2785),
    .A2(n_2827),
    .A3(n_2072),
    .B1(n_3846),
    .B2(n_1350),
    .C(n_4834),
    .Y(n_6409));
 OAI221xp5_ASAP7_75t_SL g213999 (.A1(n_4295),
    .A2(n_1389),
    .B1(n_4090),
    .B2(n_3248),
    .C(n_4845),
    .Y(n_6408));
 OAI21xp33_ASAP7_75t_L g214000 (.A1(n_1429),
    .A2(n_4300),
    .B(n_5563),
    .Y(n_6407));
 OAI32xp33_ASAP7_75t_L g214001 (.A1(n_3261),
    .A2(n_2430),
    .A3(n_2300),
    .B1(n_1371),
    .B2(n_4938),
    .Y(n_6406));
 OAI211xp5_ASAP7_75t_L g214002 (.A1(n_1556),
    .A2(n_4693),
    .B(n_4716),
    .C(n_4849),
    .Y(n_6405));
 OAI221xp5_ASAP7_75t_SL g214003 (.A1(n_4968),
    .A2(n_3389),
    .B1(n_4448),
    .B2(n_3046),
    .C(n_5321),
    .Y(n_6404));
 OAI221xp5_ASAP7_75t_L g214004 (.A1(n_3844),
    .A2(n_1558),
    .B1(n_4067),
    .B2(n_2801),
    .C(n_4858),
    .Y(n_6403));
 OAI221xp5_ASAP7_75t_L g214005 (.A1(n_1711),
    .A2(n_1467),
    .B1(n_1461),
    .B2(n_3464),
    .C(n_4794),
    .Y(n_6402));
 OAI221xp5_ASAP7_75t_SL g214006 (.A1(n_4084),
    .A2(n_2088),
    .B1(n_2800),
    .B2(n_2047),
    .C(n_6058),
    .Y(n_6401));
 OAI211xp5_ASAP7_75t_SL g214007 (.A1(n_1651),
    .A2(n_4604),
    .B(n_4707),
    .C(n_4887),
    .Y(n_6400));
 OAI211xp5_ASAP7_75t_R g214008 (.A1(n_2061),
    .A2(n_4174),
    .B(n_4972),
    .C(n_3935),
    .Y(n_6399));
 AND4x1_ASAP7_75t_L g214009 (.A(n_5443),
    .B(n_4894),
    .C(n_3196),
    .D(n_1968),
    .Y(n_6398));
 OAI211xp5_ASAP7_75t_SL g214010 (.A1(n_1543),
    .A2(n_4049),
    .B(n_4987),
    .C(n_3945),
    .Y(n_6397));
 AOI221xp5_ASAP7_75t_SL g214011 (.A1(n_4187),
    .A2(n_1622),
    .B1(n_1445),
    .B2(n_2555),
    .C(n_4969),
    .Y(n_6396));
 AOI221xp5_ASAP7_75t_R g214012 (.A1(n_4176),
    .A2(n_2402),
    .B1(n_1451),
    .B2(n_2539),
    .C(n_4945),
    .Y(n_6395));
 OAI221xp5_ASAP7_75t_L g214013 (.A1(n_2814),
    .A2(n_1986),
    .B1(n_2918),
    .B2(n_1377),
    .C(n_4791),
    .Y(n_6394));
 OAI21xp33_ASAP7_75t_L g214014 (.A1(n_1644),
    .A2(n_1777),
    .B(n_5565),
    .Y(n_6393));
 A2O1A1Ixp33_ASAP7_75t_L g214015 (.A1(n_2377),
    .A2(n_2835),
    .B(n_1501),
    .C(n_5567),
    .Y(n_6392));
 AOI211xp5_ASAP7_75t_L g214016 (.A1(n_2803),
    .A2(n_2075),
    .B(n_6149),
    .C(n_2737),
    .Y(n_6391));
 OAI211xp5_ASAP7_75t_SL g214017 (.A1(n_1582),
    .A2(n_4302),
    .B(n_5072),
    .C(n_4712),
    .Y(n_6390));
 AOI21xp33_ASAP7_75t_R g214018 (.A1(n_5096),
    .A2(n_1845),
    .B(n_4830),
    .Y(n_6389));
 OAI211xp5_ASAP7_75t_SL g214019 (.A1(n_1628),
    .A2(n_4034),
    .B(n_4936),
    .C(n_5009),
    .Y(n_6388));
 OAI321xp33_ASAP7_75t_L g214020 (.A1(n_1732),
    .A2(n_1558),
    .A3(n_2457),
    .B1(n_2066),
    .B2(n_4570),
    .C(n_5912),
    .Y(n_6387));
 OAI221xp5_ASAP7_75t_R g214021 (.A1(n_4660),
    .A2(n_1665),
    .B1(n_2395),
    .B2(n_2505),
    .C(n_4955),
    .Y(n_6386));
 NAND3xp33_ASAP7_75t_SL g214022 (.A(n_5421),
    .B(n_4826),
    .C(n_2994),
    .Y(n_6385));
 AOI221xp5_ASAP7_75t_L g214023 (.A1(n_2921),
    .A2(n_1464),
    .B1(n_1712),
    .B2(sa01[3]),
    .C(n_4793),
    .Y(n_6384));
 OAI21xp33_ASAP7_75t_L g214024 (.A1(n_1639),
    .A2(n_4286),
    .B(n_5552),
    .Y(n_6383));
 AOI221xp5_ASAP7_75t_L g214025 (.A1(n_4538),
    .A2(n_2427),
    .B1(n_2397),
    .B2(n_2501),
    .C(n_4954),
    .Y(n_6382));
 AOI221xp5_ASAP7_75t_SL g214026 (.A1(n_4581),
    .A2(n_1657),
    .B1(n_2815),
    .B2(n_3166),
    .C(n_5908),
    .Y(n_6381));
 AOI222xp33_ASAP7_75t_L g214027 (.A1(n_5172),
    .A2(n_1346),
    .B1(n_2954),
    .B2(n_2404),
    .C1(n_1419),
    .C2(n_2850),
    .Y(n_6380));
 NAND4xp25_ASAP7_75t_L g214028 (.A(n_4823),
    .B(n_4016),
    .C(n_2931),
    .D(n_3636),
    .Y(n_6379));
 OAI221xp5_ASAP7_75t_L g214029 (.A1(n_3071),
    .A2(n_1476),
    .B1(n_1639),
    .B2(n_3053),
    .C(n_5109),
    .Y(n_6378));
 AOI221xp5_ASAP7_75t_SL g214030 (.A1(n_4553),
    .A2(n_2387),
    .B1(n_3159),
    .B2(n_3241),
    .C(n_5909),
    .Y(n_6377));
 OAI221xp5_ASAP7_75t_L g214031 (.A1(n_4467),
    .A2(n_4393),
    .B1(n_4061),
    .B2(n_4468),
    .C(n_5561),
    .Y(n_6376));
 OAI221xp5_ASAP7_75t_SL g214032 (.A1(n_4467),
    .A2(n_3044),
    .B1(n_4468),
    .B2(n_2522),
    .C(n_6114),
    .Y(n_6375));
 OAI21xp33_ASAP7_75t_R g214033 (.A1(n_2068),
    .A2(n_1786),
    .B(n_6116),
    .Y(n_6374));
 O2A1O1Ixp33_ASAP7_75t_SL g214034 (.A1(n_2477),
    .A2(n_1622),
    .B(n_5350),
    .C(n_6065),
    .Y(n_6373));
 AOI211xp5_ASAP7_75t_L g214035 (.A1(n_1768),
    .A2(n_3358),
    .B(n_5668),
    .C(n_5323),
    .Y(n_6372));
 NAND4xp25_ASAP7_75t_L g214036 (.A(n_5267),
    .B(n_4549),
    .C(n_3181),
    .D(n_3676),
    .Y(n_6371));
 NOR4xp25_ASAP7_75t_SL g214037 (.A(n_6024),
    .B(n_5273),
    .C(n_4179),
    .D(n_4681),
    .Y(n_6370));
 OAI21xp33_ASAP7_75t_L g214038 (.A1(n_1417),
    .A2(n_4656),
    .B(n_6132),
    .Y(n_6369));
 OAI221xp5_ASAP7_75t_L g214039 (.A1(n_4088),
    .A2(n_1623),
    .B1(n_3075),
    .B2(n_1476),
    .C(n_4888),
    .Y(n_6368));
 OAI221xp5_ASAP7_75t_L g214040 (.A1(n_4424),
    .A2(n_2964),
    .B1(n_4422),
    .B2(n_2586),
    .C(n_6136),
    .Y(n_6367));
 AOI211xp5_ASAP7_75t_SL g214041 (.A1(n_2917),
    .A2(n_2843),
    .B(n_5523),
    .C(n_5575),
    .Y(n_6366));
 AOI211xp5_ASAP7_75t_SL g214042 (.A1(n_3930),
    .A2(n_1739),
    .B(n_5690),
    .C(n_5327),
    .Y(n_6365));
 OAI211xp5_ASAP7_75t_SL g214043 (.A1(n_1624),
    .A2(n_4563),
    .B(n_5024),
    .C(n_5514),
    .Y(n_6364));
 AOI321xp33_ASAP7_75t_L g214044 (.A1(n_2792),
    .A2(n_2416),
    .A3(n_2483),
    .B1(n_4523),
    .B2(n_2401),
    .C(n_5918),
    .Y(n_6363));
 AND3x1_ASAP7_75t_SL g214045 (.A(n_5451),
    .B(n_4827),
    .C(n_3011),
    .Y(n_6362));
 AOI211xp5_ASAP7_75t_L g214046 (.A1(n_3991),
    .A2(n_2058),
    .B(n_5539),
    .C(n_5082),
    .Y(n_6361));
 O2A1O1Ixp33_ASAP7_75t_SL g214047 (.A1(n_2353),
    .A2(n_3881),
    .B(n_1395),
    .C(n_5039),
    .Y(n_6360));
 NOR3xp33_ASAP7_75t_L g214048 (.A(n_6015),
    .B(n_3205),
    .C(n_1723),
    .Y(n_6359));
 OAI21xp5_ASAP7_75t_R g214049 (.A1(n_2059),
    .A2(n_1787),
    .B(n_6153),
    .Y(n_6358));
 AOI22xp33_ASAP7_75t_R g214050 (.A1(n_1497),
    .A2(n_5178),
    .B1(n_1432),
    .B2(n_3556),
    .Y(n_6357));
 OAI21xp33_ASAP7_75t_R g214051 (.A1(n_1582),
    .A2(n_4647),
    .B(n_6156),
    .Y(n_6356));
 A2O1A1Ixp33_ASAP7_75t_L g214052 (.A1(n_2350),
    .A2(n_3897),
    .B(n_1938),
    .C(n_5033),
    .Y(n_6355));
 NOR4xp25_ASAP7_75t_L g214053 (.A(n_6022),
    .B(n_4686),
    .C(n_4607),
    .D(n_3405),
    .Y(n_6354));
 NOR4xp25_ASAP7_75t_SL g214054 (.A(n_5413),
    .B(n_5542),
    .C(n_4177),
    .D(n_1965),
    .Y(n_6353));
 OAI21xp33_ASAP7_75t_SL g214055 (.A1(n_1450),
    .A2(n_4659),
    .B(n_6167),
    .Y(n_6352));
 NOR3xp33_ASAP7_75t_SL g214056 (.A(n_5599),
    .B(n_5530),
    .C(n_4224),
    .Y(n_6351));
 NAND4xp25_ASAP7_75t_R g214057 (.A(n_5266),
    .B(n_4529),
    .C(n_3648),
    .D(n_3202),
    .Y(n_6350));
 AOI22xp5_ASAP7_75t_SL g214058 (.A1(n_3257),
    .A2(n_4998),
    .B1(n_2082),
    .B2(n_3816),
    .Y(n_6349));
 AOI211xp5_ASAP7_75t_L g214059 (.A1(n_3951),
    .A2(n_3343),
    .B(n_5739),
    .C(n_5307),
    .Y(n_6348));
 OAI21xp33_ASAP7_75t_L g214060 (.A1(n_2061),
    .A2(n_4682),
    .B(n_5864),
    .Y(n_6347));
 OAI221xp5_ASAP7_75t_L g214061 (.A1(n_3059),
    .A2(n_3500),
    .B1(n_4007),
    .B2(n_2465),
    .C(n_6081),
    .Y(n_6346));
 AOI211xp5_ASAP7_75t_SL g214062 (.A1(n_4621),
    .A2(n_1405),
    .B(n_5023),
    .C(n_5095),
    .Y(n_6345));
 AOI211xp5_ASAP7_75t_L g214063 (.A1(n_4637),
    .A2(n_2075),
    .B(n_3738),
    .C(n_3740),
    .Y(n_6344));
 OAI221xp5_ASAP7_75t_R g214064 (.A1(n_1629),
    .A2(n_3218),
    .B1(n_3009),
    .B2(n_1522),
    .C(n_5980),
    .Y(n_6343));
 OAI21xp33_ASAP7_75t_L g214065 (.A1(n_1518),
    .A2(n_1727),
    .B(n_5860),
    .Y(n_6342));
 OAI21xp33_ASAP7_75t_L g214066 (.A1(n_8210),
    .A2(n_2802),
    .B(n_5857),
    .Y(n_6341));
 OAI221xp5_ASAP7_75t_L g214067 (.A1(n_3048),
    .A2(sa12[1]),
    .B1(n_3063),
    .B2(n_8691),
    .C(n_4857),
    .Y(n_6340));
 OAI221xp5_ASAP7_75t_SL g214068 (.A1(n_3273),
    .A2(n_8178),
    .B1(n_3593),
    .B2(n_1935),
    .C(n_4783),
    .Y(n_6339));
 OAI221xp5_ASAP7_75t_L g214069 (.A1(n_5383),
    .A2(n_1544),
    .B1(n_3907),
    .B2(n_1376),
    .C(n_3834),
    .Y(n_6338));
 OAI321xp33_ASAP7_75t_R g214070 (.A1(n_4297),
    .A2(n_2818),
    .A3(n_2061),
    .B1(n_2403),
    .B2(n_3879),
    .C(n_3835),
    .Y(n_6337));
 AOI321xp33_ASAP7_75t_L g214071 (.A1(n_4286),
    .A2(n_2042),
    .A3(n_2820),
    .B1(n_3903),
    .B2(n_1625),
    .C(n_3833),
    .Y(n_6336));
 OAI221xp5_ASAP7_75t_L g214072 (.A1(n_3545),
    .A2(n_2170),
    .B1(n_3084),
    .B2(n_1637),
    .C(n_4799),
    .Y(n_6335));
 OAI221xp5_ASAP7_75t_R g214073 (.A1(n_3477),
    .A2(n_2102),
    .B1(n_3020),
    .B2(n_2415),
    .C(n_4850),
    .Y(n_6334));
 OAI21xp33_ASAP7_75t_L g214074 (.A1(n_1450),
    .A2(n_4278),
    .B(n_5818),
    .Y(n_6333));
 OAI221xp5_ASAP7_75t_SL g214075 (.A1(n_3024),
    .A2(n_2141),
    .B1(n_2983),
    .B2(n_1442),
    .C(n_4777),
    .Y(n_6332));
 AOI221xp5_ASAP7_75t_SL g214076 (.A1(n_3098),
    .A2(n_2128),
    .B1(n_3040),
    .B2(n_2400),
    .C(n_4776),
    .Y(n_6331));
 OAI221xp5_ASAP7_75t_R g214077 (.A1(n_3116),
    .A2(n_2131),
    .B1(n_2950),
    .B2(n_1553),
    .C(n_4797),
    .Y(n_6330));
 OAI221xp5_ASAP7_75t_SL g214078 (.A1(n_2047),
    .A2(n_2130),
    .B1(n_3522),
    .B2(n_1497),
    .C(n_4773),
    .Y(n_6329));
 OAI32xp33_ASAP7_75t_L g214079 (.A1(n_3869),
    .A2(n_3758),
    .A3(n_1839),
    .B1(n_1410),
    .B2(n_3979),
    .Y(n_6328));
 OAI211xp5_ASAP7_75t_L g214080 (.A1(n_1658),
    .A2(n_4451),
    .B(n_5440),
    .C(n_5210),
    .Y(n_6327));
 OAI222xp33_ASAP7_75t_L g214081 (.A1(n_4432),
    .A2(n_2045),
    .B1(n_5098),
    .B2(n_1850),
    .C1(n_1656),
    .C2(n_2592),
    .Y(n_6326));
 OAI321xp33_ASAP7_75t_L g214082 (.A1(n_4296),
    .A2(n_3282),
    .A3(n_2068),
    .B1(n_2434),
    .B2(n_3886),
    .C(n_4804),
    .Y(n_6325));
 AOI222xp33_ASAP7_75t_R g214083 (.A1(n_5096),
    .A2(n_1461),
    .B1(n_4449),
    .B2(n_2055),
    .C1(n_1406),
    .C2(n_2590),
    .Y(n_6324));
 AOI21xp33_ASAP7_75t_L g214084 (.A1(n_3876),
    .A2(n_2044),
    .B(n_5790),
    .Y(n_6323));
 OAI222xp33_ASAP7_75t_L g214085 (.A1(n_3907),
    .A2(n_1541),
    .B1(n_3908),
    .B2(n_2073),
    .C1(n_1629),
    .C2(n_3718),
    .Y(n_6322));
 OAI222xp33_ASAP7_75t_R g214086 (.A1(n_4613),
    .A2(n_3394),
    .B1(n_5075),
    .B2(n_1456),
    .C1(n_1651),
    .C2(n_2543),
    .Y(n_6321));
 AOI221xp5_ASAP7_75t_L g214087 (.A1(n_3884),
    .A2(n_2067),
    .B1(n_3883),
    .B2(n_2435),
    .C(n_5292),
    .Y(n_6320));
 OAI211xp5_ASAP7_75t_L g214088 (.A1(n_1382),
    .A2(n_3882),
    .B(n_5163),
    .C(n_5291),
    .Y(n_6319));
 OAI22xp33_ASAP7_75t_SL g214089 (.A1(n_4907),
    .A2(n_1738),
    .B1(n_4418),
    .B2(n_1479),
    .Y(n_6318));
 AOI221xp5_ASAP7_75t_L g214090 (.A1(n_4107),
    .A2(n_1975),
    .B1(n_4108),
    .B2(sa21[3]),
    .C(n_1336),
    .Y(n_6317));
 OAI221xp5_ASAP7_75t_L g214091 (.A1(n_5097),
    .A2(n_1404),
    .B1(n_4703),
    .B2(n_3293),
    .C(n_2744),
    .Y(n_6316));
 OAI221xp5_ASAP7_75t_R g214092 (.A1(n_3022),
    .A2(n_2014),
    .B1(n_2415),
    .B2(n_2102),
    .C(n_4995),
    .Y(n_6315));
 OAI221xp5_ASAP7_75t_L g214093 (.A1(n_3085),
    .A2(n_1484),
    .B1(n_1639),
    .B2(n_2214),
    .C(n_4994),
    .Y(n_6314));
 AOI21xp33_ASAP7_75t_L g214094 (.A1(n_3956),
    .A2(n_2169),
    .B(n_5785),
    .Y(n_6313));
 OAI221xp5_ASAP7_75t_SL g214095 (.A1(n_2953),
    .A2(sa21[7]),
    .B1(n_1629),
    .B2(n_2120),
    .C(n_4980),
    .Y(n_6312));
 OAI22xp5_ASAP7_75t_R g214096 (.A1(n_3375),
    .A2(n_5110),
    .B1(n_3212),
    .B2(n_4422),
    .Y(n_6311));
 OAI221xp5_ASAP7_75t_SL g214097 (.A1(n_4738),
    .A2(sa31[6]),
    .B1(n_1397),
    .B2(n_4678),
    .C(n_3157),
    .Y(n_6310));
 OAI322xp33_ASAP7_75t_L g214098 (.A1(n_4349),
    .A2(n_3757),
    .A3(n_1501),
    .B1(n_3858),
    .B2(n_1336),
    .C1(n_1544),
    .C2(n_2536),
    .Y(n_6309));
 AOI22xp33_ASAP7_75t_R g214099 (.A1(n_1740),
    .A2(n_4891),
    .B1(n_3728),
    .B2(n_4469),
    .Y(n_6308));
 OAI221xp5_ASAP7_75t_L g214100 (.A1(n_3884),
    .A2(n_2074),
    .B1(n_3630),
    .B2(n_2497),
    .C(n_5168),
    .Y(n_6307));
 OAI222xp33_ASAP7_75t_R g214101 (.A1(n_3885),
    .A2(n_1578),
    .B1(n_3905),
    .B2(n_2126),
    .C1(n_3636),
    .C2(n_2572),
    .Y(n_6306));
 AOI221xp5_ASAP7_75t_L g214102 (.A1(n_4559),
    .A2(n_2390),
    .B1(n_1667),
    .B2(n_1670),
    .C(n_5244),
    .Y(n_6305));
 OAI221xp5_ASAP7_75t_R g214103 (.A1(n_5384),
    .A2(n_1665),
    .B1(n_3012),
    .B2(n_3328),
    .C(n_5294),
    .Y(n_6304));
 AOI221xp5_ASAP7_75t_L g214104 (.A1(n_3021),
    .A2(n_2929),
    .B1(n_4017),
    .B2(n_1680),
    .C(n_1869),
    .Y(n_6303));
 OAI221xp5_ASAP7_75t_L g214105 (.A1(n_5107),
    .A2(n_1371),
    .B1(n_1665),
    .B2(n_2593),
    .C(n_5185),
    .Y(n_6302));
 OAI22xp33_ASAP7_75t_R g214106 (.A1(n_1346),
    .A2(n_5104),
    .B1(n_1580),
    .B2(n_4104),
    .Y(n_6301));
 OAI322xp33_ASAP7_75t_L g214107 (.A1(n_2818),
    .A2(n_2570),
    .A3(n_1580),
    .B1(n_4240),
    .B2(n_2415),
    .C1(n_3869),
    .C2(n_2061),
    .Y(n_6300));
 OAI322xp33_ASAP7_75t_L g214108 (.A1(n_4347),
    .A2(n_3759),
    .A3(n_1404),
    .B1(n_4023),
    .B2(n_1934),
    .C1(n_2059),
    .C2(n_2503),
    .Y(n_6299));
 AOI211xp5_ASAP7_75t_R g214109 (.A1(n_5113),
    .A2(n_1413),
    .B(n_5277),
    .C(n_5088),
    .Y(n_6298));
 OAI322xp33_ASAP7_75t_R g214110 (.A1(n_4342),
    .A2(n_3762),
    .A3(n_1457),
    .B1(n_3986),
    .B2(n_1458),
    .C1(n_2068),
    .C2(n_2496),
    .Y(n_6297));
 OAI211xp5_ASAP7_75t_SL g214111 (.A1(n_1634),
    .A2(n_5414),
    .B(n_4761),
    .C(n_5083),
    .Y(n_6296));
 OAI322xp33_ASAP7_75t_R g214112 (.A1(n_1590),
    .A2(n_2822),
    .A3(n_2563),
    .B1(n_4370),
    .B2(n_2057),
    .C1(n_4231),
    .C2(n_1637),
    .Y(n_6295));
 OAI211xp5_ASAP7_75t_L g214113 (.A1(n_2066),
    .A2(n_5423),
    .B(n_4752),
    .C(n_5087),
    .Y(n_6294));
 OAI21xp33_ASAP7_75t_R g214114 (.A1(n_2434),
    .A2(n_5406),
    .B(n_6126),
    .Y(n_6293));
 OAI21xp33_ASAP7_75t_L g214115 (.A1(n_2422),
    .A2(n_5115),
    .B(n_6123),
    .Y(n_6292));
 AOI22xp33_ASAP7_75t_R g214116 (.A1(n_1497),
    .A2(n_5065),
    .B1(n_1432),
    .B2(n_2580),
    .Y(n_6291));
 OAI322xp33_ASAP7_75t_SL g214117 (.A1(n_1844),
    .A2(n_3755),
    .A3(n_4359),
    .B1(n_1761),
    .B2(n_1395),
    .C1(n_2053),
    .C2(n_2534),
    .Y(n_6290));
 OAI22xp33_ASAP7_75t_L g214118 (.A1(n_1498),
    .A2(n_5108),
    .B1(n_2091),
    .B2(n_4123),
    .Y(n_6289));
 OAI22xp33_ASAP7_75t_R g214119 (.A1(n_1839),
    .A2(n_5104),
    .B1(n_2061),
    .B2(n_4483),
    .Y(n_6288));
 AOI221xp5_ASAP7_75t_L g214120 (.A1(n_5068),
    .A2(n_1401),
    .B1(n_4533),
    .B2(n_1627),
    .C(n_4962),
    .Y(n_6287));
 OAI221xp5_ASAP7_75t_R g214121 (.A1(n_4667),
    .A2(n_1464),
    .B1(n_1637),
    .B2(n_2563),
    .C(n_4930),
    .Y(n_6286));
 OAI221xp5_ASAP7_75t_R g214122 (.A1(n_4550),
    .A2(n_1850),
    .B1(n_1660),
    .B2(n_2591),
    .C(n_4920),
    .Y(n_6285));
 AOI221xp5_ASAP7_75t_R g214123 (.A1(n_2046),
    .A2(n_2579),
    .B1(n_4692),
    .B2(n_1497),
    .C(n_4929),
    .Y(n_6284));
 OAI221xp5_ASAP7_75t_L g214124 (.A1(n_4677),
    .A2(n_1933),
    .B1(n_1642),
    .B2(n_2560),
    .C(n_4924),
    .Y(n_6283));
 AO332x1_ASAP7_75t_SL g214125 (.A1(n_4608),
    .A2(n_2065),
    .A3(n_1595),
    .B1(n_2800),
    .B2(n_3374),
    .B3(n_1439),
    .C1(n_4587),
    .C2(n_2089),
    .Y(n_6282));
 OAI332xp33_ASAP7_75t_L g214126 (.A1(n_4582),
    .A2(n_2403),
    .A3(n_2102),
    .B1(n_2061),
    .B2(n_2787),
    .B3(n_3357),
    .C1(n_4545),
    .C2(n_1580),
    .Y(n_6281));
 OAI221xp5_ASAP7_75t_R g214127 (.A1(n_4170),
    .A2(n_1456),
    .B1(n_8702),
    .B2(n_2544),
    .C(n_4916),
    .Y(n_6280));
 OAI221xp5_ASAP7_75t_SL g214128 (.A1(n_4561),
    .A2(n_1938),
    .B1(n_1640),
    .B2(n_2552),
    .C(n_4909),
    .Y(n_6279));
 AOI332xp33_ASAP7_75t_L g214129 (.A1(n_1603),
    .A2(n_2413),
    .A3(n_4651),
    .B1(n_3243),
    .B2(n_2077),
    .B3(n_1735),
    .C1(n_4696),
    .C2(n_2064),
    .Y(n_6278));
 OAI322xp33_ASAP7_75t_L g214130 (.A1(n_4370),
    .A2(n_3761),
    .A3(n_1464),
    .B1(n_3856),
    .B2(n_1463),
    .C1(n_1691),
    .C2(n_2057),
    .Y(n_6277));
 AOI221xp5_ASAP7_75t_L g214131 (.A1(n_4638),
    .A2(n_1498),
    .B1(n_2050),
    .B2(n_2545),
    .C(n_4906),
    .Y(n_6276));
 AOI221xp5_ASAP7_75t_R g214132 (.A1(n_4150),
    .A2(n_1500),
    .B1(n_1627),
    .B2(n_2574),
    .C(n_4905),
    .Y(n_6275));
 AOI22xp5_ASAP7_75t_R g214133 (.A1(n_1458),
    .A2(n_1789),
    .B1(n_2558),
    .B2(n_1405),
    .Y(n_6274));
 AOI322xp5_ASAP7_75t_L g214134 (.A1(n_3763),
    .A2(n_4368),
    .A3(n_1497),
    .B1(n_3848),
    .B2(n_1496),
    .C1(n_1439),
    .C2(n_2511),
    .Y(n_6273));
 AOI332xp33_ASAP7_75t_L g214135 (.A1(n_4617),
    .A2(n_1655),
    .A3(n_2095),
    .B1(n_2805),
    .B2(n_2044),
    .B3(n_1736),
    .C1(n_4635),
    .C2(n_1576),
    .Y(n_6272));
 OAI22xp33_ASAP7_75t_R g214136 (.A1(n_2053),
    .A2(n_5393),
    .B1(n_2428),
    .B2(n_3894),
    .Y(n_6271));
 OAI211xp5_ASAP7_75t_SL g214137 (.A1(n_1623),
    .A2(n_5429),
    .B(n_5514),
    .C(n_4763),
    .Y(n_6270));
 OAI21xp33_ASAP7_75t_L g214138 (.A1(n_1464),
    .A2(n_5086),
    .B(n_5212),
    .Y(n_6269));
 OAI211xp5_ASAP7_75t_L g214139 (.A1(n_2424),
    .A2(n_5431),
    .B(n_5300),
    .C(n_5509),
    .Y(n_6268));
 AOI322xp5_ASAP7_75t_SL g214140 (.A1(n_1713),
    .A2(n_1734),
    .A3(n_2058),
    .B1(n_1589),
    .B2(n_4558),
    .C1(n_5063),
    .C2(n_1667),
    .Y(n_6267));
 OAI322xp33_ASAP7_75t_R g214141 (.A1(n_3347),
    .A2(n_1548),
    .A3(n_2806),
    .B1(n_2083),
    .B2(n_4554),
    .C1(n_1634),
    .C2(n_5061),
    .Y(n_6266));
 AOI221xp5_ASAP7_75t_L g214142 (.A1(n_4148),
    .A2(n_2873),
    .B1(n_4088),
    .B2(n_2042),
    .C(n_4915),
    .Y(n_6265));
 OAI321xp33_ASAP7_75t_L g214143 (.A1(n_2059),
    .A2(n_3330),
    .A3(n_3259),
    .B1(n_5049),
    .B2(n_2422),
    .C(n_4846),
    .Y(n_6264));
 AOI21xp33_ASAP7_75t_L g214144 (.A1(n_5068),
    .A2(n_2425),
    .B(n_5605),
    .Y(n_6263));
 OAI322xp33_ASAP7_75t_L g214145 (.A1(n_3248),
    .A2(n_2068),
    .A3(n_3320),
    .B1(n_4060),
    .B2(n_2074),
    .C1(n_5057),
    .C2(n_2434),
    .Y(n_6262));
 AOI322xp5_ASAP7_75t_L g214146 (.A1(n_3253),
    .A2(n_3370),
    .A3(n_2054),
    .B1(n_2082),
    .B2(n_4592),
    .C1(n_5056),
    .C2(n_1413),
    .Y(n_6261));
 OAI322xp33_ASAP7_75t_SL g214147 (.A1(n_2778),
    .A2(n_3368),
    .A3(n_1390),
    .B1(n_4640),
    .B2(n_1381),
    .C1(n_1623),
    .C2(n_5066),
    .Y(n_6260));
 AOI311xp33_ASAP7_75t_SL g214148 (.A1(n_2785),
    .A2(n_2827),
    .A3(n_1350),
    .B(n_4248),
    .C(n_4536),
    .Y(n_6259));
 AOI322xp5_ASAP7_75t_L g214149 (.A1(n_1728),
    .A2(n_3385),
    .A3(n_1559),
    .B1(n_1412),
    .B2(n_4596),
    .C1(n_1788),
    .C2(n_1348),
    .Y(n_6258));
 AOI22xp33_ASAP7_75t_L g214150 (.A1(n_2075),
    .A2(n_5058),
    .B1(n_1422),
    .B2(n_4457),
    .Y(n_6257));
 OAI22xp5_ASAP7_75t_SL g214151 (.A1(n_1934),
    .A2(n_5097),
    .B1(n_2080),
    .B2(n_4138),
    .Y(n_6450));
 OAI322xp33_ASAP7_75t_R g214152 (.A1(n_3256),
    .A2(n_2081),
    .A3(n_2548),
    .B1(n_4359),
    .B2(n_2053),
    .C1(n_4266),
    .C2(n_1443),
    .Y(n_6256));
 OAI322xp33_ASAP7_75t_SL g214153 (.A1(n_2780),
    .A2(n_1742),
    .A3(n_2056),
    .B1(n_4674),
    .B2(n_1342),
    .C1(n_5070),
    .C2(n_1408),
    .Y(n_6255));
 OAI321xp33_ASAP7_75t_L g214154 (.A1(n_3277),
    .A2(n_2080),
    .A3(n_2550),
    .B1(n_2059),
    .B2(n_4347),
    .C(n_4935),
    .Y(n_6254));
 AOI322xp5_ASAP7_75t_L g214155 (.A1(n_4345),
    .A2(n_3764),
    .A3(n_1935),
    .B1(n_3141),
    .B2(n_3371),
    .C1(n_1552),
    .C2(n_2526),
    .Y(n_6253));
 OAI322xp33_ASAP7_75t_SL g214156 (.A1(n_3245),
    .A2(n_1571),
    .A3(n_2590),
    .B1(n_1654),
    .B2(n_4246),
    .C1(n_4366),
    .C2(n_1417),
    .Y(n_6252));
 AO22x1_ASAP7_75t_L g214157 (.A1(n_1395),
    .A2(n_5106),
    .B1(n_3281),
    .B2(n_4182),
    .Y(n_6251));
 AOI322xp5_ASAP7_75t_R g214158 (.A1(n_3260),
    .A2(n_3321),
    .A3(n_1552),
    .B1(n_2092),
    .B2(n_4593),
    .C1(n_4661),
    .C2(n_3184),
    .Y(n_6250));
 OAI221xp5_ASAP7_75t_SL g214159 (.A1(n_4081),
    .A2(n_1546),
    .B1(n_3995),
    .B2(n_1634),
    .C(n_4900),
    .Y(n_6249));
 OAI221xp5_ASAP7_75t_R g214160 (.A1(n_3958),
    .A2(n_1651),
    .B1(n_4101),
    .B2(n_1582),
    .C(n_4927),
    .Y(n_6248));
 AOI322xp5_ASAP7_75t_L g214161 (.A1(n_3283),
    .A2(n_2557),
    .A3(n_2075),
    .B1(n_1444),
    .B2(n_1780),
    .C1(n_2400),
    .C2(n_4265),
    .Y(n_6247));
 OAI211xp5_ASAP7_75t_L g214162 (.A1(n_2063),
    .A2(n_4291),
    .B(n_5412),
    .C(n_2679),
    .Y(n_6246));
 OAI22xp5_ASAP7_75t_SL g214163 (.A1(n_1499),
    .A2(n_5108),
    .B1(n_3286),
    .B2(n_4158),
    .Y(n_6245));
 AOI321xp33_ASAP7_75t_L g214164 (.A1(n_3257),
    .A2(n_3281),
    .A3(n_1415),
    .B1(n_4102),
    .B2(n_1440),
    .C(n_4958),
    .Y(n_6244));
 OAI32xp33_ASAP7_75t_SL g214165 (.A1(n_4732),
    .A2(n_3336),
    .A3(n_1336),
    .B1(n_2073),
    .B2(n_4236),
    .Y(n_6243));
 AOI321xp33_ASAP7_75t_SL g214166 (.A1(n_3254),
    .A2(n_3287),
    .A3(n_1349),
    .B1(n_4103),
    .B2(n_1561),
    .C(n_4932),
    .Y(n_6242));
 OAI221xp5_ASAP7_75t_R g214167 (.A1(n_3061),
    .A2(n_2102),
    .B1(n_4098),
    .B2(n_2850),
    .C(n_4531),
    .Y(n_6241));
 AOI211xp5_ASAP7_75t_L g214168 (.A1(n_4299),
    .A2(n_1586),
    .B(n_5428),
    .C(n_2661),
    .Y(n_6240));
 AOI211xp5_ASAP7_75t_L g214169 (.A1(n_4296),
    .A2(n_1423),
    .B(n_5114),
    .C(n_2652),
    .Y(n_6239));
 OAI22xp33_ASAP7_75t_R g214170 (.A1(n_1628),
    .A2(n_5471),
    .B1(n_1355),
    .B2(n_3097),
    .Y(n_6238));
 OAI311xp33_ASAP7_75t_SL g214171 (.A1(n_3296),
    .A2(n_3248),
    .A3(n_1389),
    .B1(n_3842),
    .C1(n_4522),
    .Y(n_6237));
 AOI211xp5_ASAP7_75t_SL g214172 (.A1(n_4327),
    .A2(n_1572),
    .B(n_5415),
    .C(n_2677),
    .Y(n_6236));
 OAI22xp33_ASAP7_75t_R g214173 (.A1(n_1938),
    .A2(n_5105),
    .B1(n_3413),
    .B2(n_4055),
    .Y(n_6235));
 OAI221xp5_ASAP7_75t_L g214174 (.A1(n_4193),
    .A2(n_1429),
    .B1(n_1726),
    .B2(n_1584),
    .C(n_5644),
    .Y(n_6234));
 INVxp67_ASAP7_75t_R g214175 (.A(n_5901),
    .Y(n_6231));
 INVxp67_ASAP7_75t_R g214176 (.A(n_6225),
    .Y(n_6226));
 INVxp67_ASAP7_75t_L g214177 (.A(n_6220),
    .Y(n_6221));
 INVxp67_ASAP7_75t_R g214178 (.A(n_6217),
    .Y(n_6218));
 INVxp67_ASAP7_75t_R g214179 (.A(n_6210),
    .Y(n_6211));
 INVxp67_ASAP7_75t_L g214180 (.A(n_6203),
    .Y(n_6204));
 INVxp67_ASAP7_75t_L g214182 (.A(n_6198),
    .Y(n_6199));
 INVxp67_ASAP7_75t_L g214184 (.A(n_6195),
    .Y(n_6196));
 INVxp67_ASAP7_75t_R g214185 (.A(n_6191),
    .Y(n_6192));
 INVxp67_ASAP7_75t_L g214186 (.A(n_6187),
    .Y(n_6188));
 INVx1_ASAP7_75t_L g214187 (.A(n_6185),
    .Y(n_6186));
 INVxp67_ASAP7_75t_R g214189 (.A(n_6183),
    .Y(n_6184));
 INVxp67_ASAP7_75t_L g214190 (.A(n_6182),
    .Y(n_6181));
 INVxp67_ASAP7_75t_L g214191 (.A(n_6180),
    .Y(n_6179));
 INVxp67_ASAP7_75t_R g214192 (.A(n_6177),
    .Y(n_6178));
 HB1xp67_ASAP7_75t_SL g214193 (.A(n_6174),
    .Y(n_6175));
 INVx1_ASAP7_75t_R g214195 (.A(n_6173),
    .Y(n_1794));
 NAND2xp5_ASAP7_75t_L g214196 (.A(sa12[2]),
    .B(n_5072),
    .Y(n_6169));
 NAND2xp33_ASAP7_75t_R g214197 (.A(n_1501),
    .B(n_5103),
    .Y(n_6168));
 OAI21xp33_ASAP7_75t_SL g214198 (.A1(n_2473),
    .A2(n_1655),
    .B(n_5338),
    .Y(n_6167));
 AOI221xp5_ASAP7_75t_L g214199 (.A1(n_2404),
    .A2(n_4104),
    .B1(n_2878),
    .B2(sa33[3]),
    .C(n_3814),
    .Y(n_6166));
 AOI211xp5_ASAP7_75t_L g214200 (.A1(n_3118),
    .A2(n_2077),
    .B(n_4709),
    .C(n_2610),
    .Y(n_6165));
 AOI211xp5_ASAP7_75t_L g214201 (.A1(n_3134),
    .A2(n_2462),
    .B(n_4879),
    .C(n_4691),
    .Y(n_6164));
 NOR3xp33_ASAP7_75t_L g214202 (.A(n_1768),
    .B(n_5301),
    .C(n_4159),
    .Y(n_6163));
 O2A1O1Ixp33_ASAP7_75t_R g214203 (.A1(n_2173),
    .A2(n_2904),
    .B(n_1984),
    .C(n_3739),
    .Y(n_6162));
 OAI211xp5_ASAP7_75t_L g214204 (.A1(n_1647),
    .A2(n_3920),
    .B(n_3775),
    .C(n_4609),
    .Y(n_6161));
 OAI21xp33_ASAP7_75t_R g214205 (.A1(n_2485),
    .A2(n_1633),
    .B(n_5333),
    .Y(n_6160));
 AOI211xp5_ASAP7_75t_SL g214206 (.A1(n_3236),
    .A2(n_2378),
    .B(n_4361),
    .C(n_1938),
    .Y(n_6159));
 AOI22xp33_ASAP7_75t_R g214207 (.A1(n_2543),
    .A2(n_4022),
    .B1(n_2414),
    .B2(n_4239),
    .Y(n_6158));
 OAI31xp33_ASAP7_75t_R g214208 (.A1(n_3263),
    .A2(n_2544),
    .A3(n_1512),
    .B(n_5036),
    .Y(n_6157));
 OAI22xp33_ASAP7_75t_R g214209 (.A1(n_2482),
    .A2(n_4232),
    .B1(n_2414),
    .B2(n_2481),
    .Y(n_6156));
 AOI22xp33_ASAP7_75t_L g214210 (.A1(n_1781),
    .A2(n_1446),
    .B1(n_1627),
    .B2(n_3238),
    .Y(n_6155));
 OAI21xp33_ASAP7_75t_R g214211 (.A1(n_1665),
    .A2(n_4414),
    .B(n_3750),
    .Y(n_6154));
 OAI21xp33_ASAP7_75t_R g214212 (.A1(n_2450),
    .A2(n_2421),
    .B(n_5339),
    .Y(n_6153));
 OAI22xp33_ASAP7_75t_R g214213 (.A1(n_2061),
    .A2(n_4237),
    .B1(n_2570),
    .B2(n_2415),
    .Y(n_6152));
 O2A1O1Ixp33_ASAP7_75t_R g214214 (.A1(n_2550),
    .A2(n_3311),
    .B(n_1352),
    .C(n_2745),
    .Y(n_6151));
 NAND2xp33_ASAP7_75t_R g214215 (.A(n_3712),
    .B(n_1790),
    .Y(n_6150));
 NAND2xp5_ASAP7_75t_R g214216 (.A(n_2962),
    .B(n_5424),
    .Y(n_6149));
 NAND2xp33_ASAP7_75t_R g214217 (.A(n_1459),
    .B(n_1789),
    .Y(n_6148));
 NAND2xp5_ASAP7_75t_L g214218 (.A(n_2090),
    .B(n_1788),
    .Y(n_6147));
 OAI211xp5_ASAP7_75t_L g214219 (.A1(n_1559),
    .A2(n_2746),
    .B(n_3254),
    .C(n_3287),
    .Y(n_6146));
 NAND2xp33_ASAP7_75t_R g214220 (.A(n_2410),
    .B(n_5390),
    .Y(n_6145));
 NOR2xp33_ASAP7_75t_R g214221 (.A(n_4765),
    .B(n_5082),
    .Y(n_6144));
 AOI21xp33_ASAP7_75t_L g214222 (.A1(n_4445),
    .A2(n_1622),
    .B(n_3743),
    .Y(n_6143));
 A2O1A1Ixp33_ASAP7_75t_L g214223 (.A1(n_1914),
    .A2(n_1691),
    .B(n_1637),
    .C(n_4822),
    .Y(n_6142));
 AOI211xp5_ASAP7_75t_R g214224 (.A1(n_3093),
    .A2(n_1447),
    .B(n_4908),
    .C(n_3934),
    .Y(n_6141));
 NOR2xp33_ASAP7_75t_L g214225 (.A(n_1363),
    .B(n_5400),
    .Y(n_6140));
 NOR3xp33_ASAP7_75t_SL g214226 (.A(n_5092),
    .B(n_3245),
    .C(n_3766),
    .Y(n_6139));
 OAI221xp5_ASAP7_75t_SL g214227 (.A1(n_3013),
    .A2(n_1658),
    .B1(n_3057),
    .B2(n_1662),
    .C(n_4739),
    .Y(n_6138));
 OAI21xp33_ASAP7_75t_R g214228 (.A1(n_1408),
    .A2(n_4506),
    .B(n_3746),
    .Y(n_6137));
 AOI22xp33_ASAP7_75t_R g214229 (.A1(n_3376),
    .A2(n_3938),
    .B1(n_2748),
    .B2(n_4480),
    .Y(n_6136));
 O2A1O1Ixp33_ASAP7_75t_R g214230 (.A1(n_2590),
    .A2(n_3298),
    .B(n_2055),
    .C(n_2741),
    .Y(n_6135));
 AOI22xp33_ASAP7_75t_R g214231 (.A1(n_2401),
    .A2(n_4410),
    .B1(n_1451),
    .B2(n_3239),
    .Y(n_6134));
 NAND2xp5_ASAP7_75t_L g214232 (.A(n_2398),
    .B(n_5455),
    .Y(n_6133));
 OAI22xp5_ASAP7_75t_R g214233 (.A1(n_2468),
    .A2(n_4235),
    .B1(n_2410),
    .B2(n_2467),
    .Y(n_6132));
 NOR2xp33_ASAP7_75t_R g214234 (.A(n_1568),
    .B(n_5112),
    .Y(n_6131));
 AOI211xp5_ASAP7_75t_R g214235 (.A1(n_3115),
    .A2(n_1433),
    .B(n_4971),
    .C(n_3797),
    .Y(n_6130));
 AOI21xp33_ASAP7_75t_R g214236 (.A1(n_4307),
    .A2(n_1699),
    .B(n_1624),
    .Y(n_6129));
 AOI221xp5_ASAP7_75t_SL g214237 (.A1(n_2416),
    .A2(n_2946),
    .B1(n_2062),
    .B2(n_2304),
    .C(n_4742),
    .Y(n_6128));
 OAI221xp5_ASAP7_75t_L g214238 (.A1(n_3035),
    .A2(n_1639),
    .B1(n_1390),
    .B2(n_2324),
    .C(n_4736),
    .Y(n_6127));
 NOR2xp33_ASAP7_75t_R g214239 (.A(n_5095),
    .B(n_5295),
    .Y(n_6126));
 OAI21xp33_ASAP7_75t_L g214240 (.A1(n_1859),
    .A2(n_3855),
    .B(n_4984),
    .Y(n_6125));
 OAI21xp33_ASAP7_75t_R g214241 (.A1(n_1668),
    .A2(n_2442),
    .B(n_5335),
    .Y(n_6124));
 NOR3xp33_ASAP7_75t_L g214242 (.A(n_5094),
    .B(n_3770),
    .C(n_3277),
    .Y(n_6123));
 OAI211xp5_ASAP7_75t_L g214243 (.A1(n_1568),
    .A2(n_3997),
    .B(n_4606),
    .C(n_3777),
    .Y(n_6122));
 AOI22xp33_ASAP7_75t_R g214244 (.A1(n_1435),
    .A2(n_4362),
    .B1(n_1641),
    .B2(n_4250),
    .Y(n_6121));
 O2A1O1Ixp33_ASAP7_75t_R g214245 (.A1(n_2443),
    .A2(n_3001),
    .B(n_2389),
    .C(n_3792),
    .Y(n_6120));
 AOI22xp33_ASAP7_75t_L g214246 (.A1(n_2574),
    .A2(n_4021),
    .B1(n_1446),
    .B2(n_4244),
    .Y(n_6119));
 OAI221xp5_ASAP7_75t_R g214247 (.A1(n_1628),
    .A2(n_2915),
    .B1(n_1541),
    .B2(n_1705),
    .C(n_5003),
    .Y(n_6118));
 O2A1O1Ixp33_ASAP7_75t_R g214248 (.A1(n_2558),
    .A2(n_3248),
    .B(n_2435),
    .C(n_5228),
    .Y(n_6117));
 OAI22xp33_ASAP7_75t_R g214249 (.A1(n_2438),
    .A2(n_4228),
    .B1(n_2435),
    .B2(n_2439),
    .Y(n_6116));
 OAI21xp33_ASAP7_75t_R g214250 (.A1(n_2475),
    .A2(n_2425),
    .B(n_5373),
    .Y(n_6115));
 AOI21xp5_ASAP7_75t_L g214251 (.A1(n_3932),
    .A2(n_1740),
    .B(n_5317),
    .Y(n_6114));
 AOI22xp33_ASAP7_75t_R g214252 (.A1(n_2067),
    .A2(n_4241),
    .B1(n_2557),
    .B2(n_1422),
    .Y(n_6113));
 OAI211xp5_ASAP7_75t_L g214253 (.A1(n_1541),
    .A2(n_3143),
    .B(n_4933),
    .C(n_3791),
    .Y(n_6112));
 A2O1A1Ixp33_ASAP7_75t_L g214254 (.A1(n_2847),
    .A2(n_2796),
    .B(n_2047),
    .C(n_4019),
    .Y(n_6111));
 OAI221xp5_ASAP7_75t_SL g214255 (.A1(n_2950),
    .A2(n_2066),
    .B1(n_2960),
    .B2(n_1558),
    .C(n_4743),
    .Y(n_6110));
 AOI221xp5_ASAP7_75t_SL g214256 (.A1(n_3531),
    .A2(n_2386),
    .B1(n_3160),
    .B2(n_1547),
    .C(n_5037),
    .Y(n_6109));
 AOI221xp5_ASAP7_75t_R g214257 (.A1(n_2921),
    .A2(n_1667),
    .B1(n_3170),
    .B2(n_2058),
    .C(n_4979),
    .Y(n_6108));
 NAND2xp33_ASAP7_75t_R g214258 (.A(n_1416),
    .B(n_1793),
    .Y(n_6107));
 O2A1O1Ixp33_ASAP7_75t_L g214259 (.A1(sa11[3]),
    .A2(n_2842),
    .B(n_4259),
    .C(sa11[6]),
    .Y(n_6106));
 O2A1O1Ixp33_ASAP7_75t_R g214260 (.A1(sa00[3]),
    .A2(n_3298),
    .B(n_4260),
    .C(n_1461),
    .Y(n_6105));
 O2A1O1Ixp33_ASAP7_75t_L g214261 (.A1(n_3342),
    .A2(n_3256),
    .B(sa22[3]),
    .C(n_4817),
    .Y(n_6104));
 A2O1A1Ixp33_ASAP7_75t_L g214262 (.A1(n_3284),
    .A2(n_1745),
    .B(n_8178),
    .C(n_4818),
    .Y(n_6103));
 OAI211xp5_ASAP7_75t_R g214263 (.A1(n_2306),
    .A2(n_2047),
    .B(n_4542),
    .C(n_3667),
    .Y(n_6102));
 O2A1O1Ixp33_ASAP7_75t_L g214264 (.A1(n_3357),
    .A2(n_3490),
    .B(n_1577),
    .C(n_4212),
    .Y(n_6101));
 O2A1O1Ixp33_ASAP7_75t_R g214265 (.A1(n_3345),
    .A2(n_2818),
    .B(sa33[3]),
    .C(n_4779),
    .Y(n_6100));
 OAI221xp5_ASAP7_75t_R g214266 (.A1(n_2992),
    .A2(sa01[7]),
    .B1(n_2388),
    .B2(n_2170),
    .C(n_4997),
    .Y(n_6099));
 A2O1A1Ixp33_ASAP7_75t_L g214267 (.A1(n_1979),
    .A2(n_2840),
    .B(n_3771),
    .C(n_1839),
    .Y(n_6098));
 A2O1A1Ixp33_ASAP7_75t_R g214268 (.A1(n_1971),
    .A2(n_3308),
    .B(n_3772),
    .C(n_1456),
    .Y(n_6097));
 OAI21xp33_ASAP7_75t_L g214269 (.A1(n_2725),
    .A2(n_4633),
    .B(n_1395),
    .Y(n_6096));
 OAI21xp5_ASAP7_75t_R g214270 (.A1(n_2727),
    .A2(n_4611),
    .B(n_1935),
    .Y(n_6095));
 O2A1O1Ixp33_ASAP7_75t_R g214271 (.A1(n_1716),
    .A2(n_3245),
    .B(sa00[3]),
    .C(n_4802),
    .Y(n_6094));
 O2A1O1Ixp33_ASAP7_75t_L g214272 (.A1(n_1747),
    .A2(n_3263),
    .B(n_1512),
    .C(n_4809),
    .Y(n_6093));
 NAND2xp33_ASAP7_75t_R g214273 (.A(n_5077),
    .B(n_3749),
    .Y(n_6092));
 O2A1O1Ixp33_ASAP7_75t_L g214274 (.A1(sa01[7]),
    .A2(n_2563),
    .B(n_2390),
    .C(n_5080),
    .Y(n_6091));
 AOI22xp33_ASAP7_75t_R g214275 (.A1(n_3765),
    .A2(n_4051),
    .B1(n_3206),
    .B2(n_1986),
    .Y(n_6090));
 NAND3xp33_ASAP7_75t_R g214276 (.A(n_4699),
    .B(n_3191),
    .C(n_3657),
    .Y(n_6089));
 OAI211xp5_ASAP7_75t_SL g214277 (.A1(sa21[3]),
    .A2(n_1677),
    .B(n_5500),
    .C(n_4211),
    .Y(n_6088));
 OAI221xp5_ASAP7_75t_L g214278 (.A1(n_3153),
    .A2(n_1556),
    .B1(n_2047),
    .B2(n_3540),
    .C(n_4644),
    .Y(n_6087));
 O2A1O1Ixp33_ASAP7_75t_R g214279 (.A1(n_3330),
    .A2(n_3497),
    .B(n_1586),
    .C(n_4601),
    .Y(n_6086));
 OAI21xp33_ASAP7_75t_R g214280 (.A1(n_3596),
    .A2(n_4386),
    .B(n_2712),
    .Y(n_6085));
 O2A1O1Ixp33_ASAP7_75t_R g214281 (.A1(n_3317),
    .A2(n_3475),
    .B(n_1589),
    .C(n_4190),
    .Y(n_6084));
 OAI21xp5_ASAP7_75t_SL g214282 (.A1(n_2424),
    .A2(n_4463),
    .B(n_2668),
    .Y(n_6083));
 AOI211xp5_ASAP7_75t_SL g214283 (.A1(n_3754),
    .A2(n_3435),
    .B(n_3336),
    .C(n_1501),
    .Y(n_6082));
 AOI221xp5_ASAP7_75t_R g214284 (.A1(n_1444),
    .A2(n_2522),
    .B1(n_1421),
    .B2(n_3237),
    .C(n_1857),
    .Y(n_6081));
 A2O1A1Ixp33_ASAP7_75t_R g214285 (.A1(n_1736),
    .A2(n_1755),
    .B(n_1344),
    .C(n_4200),
    .Y(n_6080));
 OAI211xp5_ASAP7_75t_R g214286 (.A1(n_1760),
    .A2(n_1637),
    .B(n_3916),
    .C(n_2152),
    .Y(n_6079));
 O2A1O1Ixp33_ASAP7_75t_L g214287 (.A1(n_1534),
    .A2(n_2580),
    .B(n_1554),
    .C(n_5436),
    .Y(n_6078));
 AOI211xp5_ASAP7_75t_R g214288 (.A1(n_3210),
    .A2(n_1645),
    .B(n_3038),
    .C(n_3807),
    .Y(n_6077));
 NAND3xp33_ASAP7_75t_R g214289 (.A(n_5391),
    .B(n_1416),
    .C(sa00[0]),
    .Y(n_6076));
 O2A1O1Ixp33_ASAP7_75t_R g214290 (.A1(n_3296),
    .A2(n_3282),
    .B(n_2067),
    .C(n_5258),
    .Y(n_6075));
 A2O1A1Ixp33_ASAP7_75t_R g214291 (.A1(sa11[6]),
    .A2(n_2844),
    .B(n_2429),
    .C(n_5405),
    .Y(n_6074));
 AOI211xp5_ASAP7_75t_L g214292 (.A1(n_1436),
    .A2(n_3216),
    .B(n_1723),
    .C(n_3818),
    .Y(n_6073));
 NAND3xp33_ASAP7_75t_R g214293 (.A(n_1791),
    .B(n_2039),
    .C(n_1866),
    .Y(n_6072));
 AOI211xp5_ASAP7_75t_R g214294 (.A1(n_1627),
    .A2(n_3158),
    .B(n_3002),
    .C(n_3810),
    .Y(n_6071));
 A2O1A1Ixp33_ASAP7_75t_R g214295 (.A1(n_1935),
    .A2(n_3313),
    .B(n_1449),
    .C(n_5048),
    .Y(n_6070));
 AOI211xp5_ASAP7_75t_L g214296 (.A1(n_2963),
    .A2(n_2410),
    .B(n_4687),
    .C(n_3554),
    .Y(n_6069));
 A2O1A1Ixp33_ASAP7_75t_L g214297 (.A1(n_1455),
    .A2(n_3290),
    .B(n_8690),
    .C(n_5403),
    .Y(n_6068));
 A2O1A1Ixp33_ASAP7_75t_L g214298 (.A1(n_1346),
    .A2(n_2850),
    .B(n_1451),
    .C(n_5395),
    .Y(n_6067));
 O2A1O1Ixp33_ASAP7_75t_SL g214299 (.A1(n_2829),
    .A2(n_3277),
    .B(n_1431),
    .C(n_5275),
    .Y(n_6066));
 OAI21xp33_ASAP7_75t_SL g214300 (.A1(n_2043),
    .A2(n_4662),
    .B(n_5504),
    .Y(n_6065));
 AOI22xp33_ASAP7_75t_SL g214301 (.A1(n_2046),
    .A2(n_4368),
    .B1(n_2847),
    .B2(n_2976),
    .Y(n_6064));
 AOI21xp33_ASAP7_75t_R g214302 (.A1(n_4028),
    .A2(n_1374),
    .B(n_1528),
    .Y(n_6063));
 NAND3xp33_ASAP7_75t_R g214303 (.A(n_5394),
    .B(n_1542),
    .C(sa21[0]),
    .Y(n_6062));
 OAI21xp33_ASAP7_75t_R g214304 (.A1(n_1383),
    .A2(n_4381),
    .B(n_2653),
    .Y(n_6061));
 NOR3xp33_ASAP7_75t_L g214305 (.A(n_5278),
    .B(n_4666),
    .C(n_4076),
    .Y(n_6060));
 OAI221xp5_ASAP7_75t_R g214306 (.A1(n_1758),
    .A2(n_1986),
    .B1(n_1662),
    .B2(n_1387),
    .C(n_1739),
    .Y(n_6059));
 AOI21xp5_ASAP7_75t_R g214307 (.A1(n_4505),
    .A2(n_1432),
    .B(n_5133),
    .Y(n_6058));
 AOI221xp5_ASAP7_75t_SL g214308 (.A1(n_3020),
    .A2(n_1346),
    .B1(n_1451),
    .B2(n_2127),
    .C(n_5495),
    .Y(n_6057));
 OAI322xp33_ASAP7_75t_L g214309 (.A1(n_2280),
    .A2(n_2422),
    .A3(n_3259),
    .B1(n_2001),
    .B2(n_2080),
    .C1(n_1403),
    .C2(n_4233),
    .Y(n_6056));
 NAND3xp33_ASAP7_75t_L g214310 (.A(n_5069),
    .B(n_4625),
    .C(n_4178),
    .Y(n_6055));
 AOI21xp5_ASAP7_75t_SL g214311 (.A1(n_3017),
    .A2(n_3361),
    .B(n_5446),
    .Y(n_6054));
 AOI211xp5_ASAP7_75t_R g214312 (.A1(n_1712),
    .A2(n_1447),
    .B(n_4153),
    .C(n_1877),
    .Y(n_6053));
 OAI31xp33_ASAP7_75t_R g214313 (.A1(n_2868),
    .A2(n_3001),
    .A3(n_2822),
    .B(n_2431),
    .Y(n_6052));
 O2A1O1Ixp33_ASAP7_75t_R g214314 (.A1(n_2580),
    .A2(n_2801),
    .B(n_1432),
    .C(n_5452),
    .Y(n_6051));
 OAI211xp5_ASAP7_75t_SL g214315 (.A1(n_1644),
    .A2(n_3213),
    .B(n_3922),
    .C(n_2627),
    .Y(n_6050));
 A2O1A1Ixp33_ASAP7_75t_R g214316 (.A1(n_2564),
    .A2(n_2813),
    .B(n_1666),
    .C(n_5459),
    .Y(n_6049));
 OAI321xp33_ASAP7_75t_R g214317 (.A1(n_2168),
    .A2(n_1938),
    .A3(n_1484),
    .B1(n_8177),
    .B2(n_2884),
    .C(n_1640),
    .Y(n_6048));
 OAI211xp5_ASAP7_75t_L g214318 (.A1(n_2098),
    .A2(n_1654),
    .B(n_1721),
    .C(n_4646),
    .Y(n_6047));
 OAI211xp5_ASAP7_75t_SL g214319 (.A1(n_1429),
    .A2(n_3603),
    .B(n_3925),
    .C(n_2202),
    .Y(n_6046));
 OAI211xp5_ASAP7_75t_L g214320 (.A1(n_1496),
    .A2(n_3570),
    .B(n_3667),
    .C(n_1509),
    .Y(n_6045));
 OAI21xp33_ASAP7_75t_R g214321 (.A1(n_2430),
    .A2(n_4316),
    .B(n_3129),
    .Y(n_6044));
 AOI211xp5_ASAP7_75t_L g214322 (.A1(n_3067),
    .A2(n_8690),
    .B(n_3924),
    .C(n_2237),
    .Y(n_6043));
 AOI211xp5_ASAP7_75t_R g214323 (.A1(n_2925),
    .A2(n_2404),
    .B(n_4273),
    .C(n_3806),
    .Y(n_6042));
 OAI221xp5_ASAP7_75t_R g214324 (.A1(n_1646),
    .A2(n_2742),
    .B1(n_2061),
    .B2(n_3088),
    .C(n_3935),
    .Y(n_6041));
 AOI21xp5_ASAP7_75t_L g214325 (.A1(n_4470),
    .A2(n_1499),
    .B(n_1561),
    .Y(n_6040));
 OAI211xp5_ASAP7_75t_R g214326 (.A1(n_2399),
    .A2(n_3062),
    .B(n_3931),
    .C(n_2224),
    .Y(n_6039));
 AOI221xp5_ASAP7_75t_L g214327 (.A1(n_4584),
    .A2(n_1432),
    .B1(n_1731),
    .B2(n_1438),
    .C(n_1509),
    .Y(n_6038));
 O2A1O1Ixp33_ASAP7_75t_R g214328 (.A1(n_3345),
    .A2(n_2787),
    .B(n_2401),
    .C(n_2663),
    .Y(n_6037));
 OAI21xp33_ASAP7_75t_L g214329 (.A1(n_2041),
    .A2(n_3891),
    .B(n_5276),
    .Y(n_6036));
 OAI21xp33_ASAP7_75t_R g214330 (.A1(n_1498),
    .A2(n_3853),
    .B(n_1981),
    .Y(n_6035));
 AOI21xp33_ASAP7_75t_R g214331 (.A1(n_1682),
    .A2(n_4015),
    .B(n_8213),
    .Y(n_6034));
 O2A1O1Ixp33_ASAP7_75t_R g214332 (.A1(n_2486),
    .A2(n_3242),
    .B(n_2084),
    .C(n_1866),
    .Y(n_6033));
 OA21x2_ASAP7_75t_R g214333 (.A1(n_3394),
    .A2(n_3089),
    .B(n_5288),
    .Y(n_6032));
 AOI211xp5_ASAP7_75t_L g214334 (.A1(n_3729),
    .A2(n_2397),
    .B(n_3921),
    .C(n_2204),
    .Y(n_6031));
 AOI211xp5_ASAP7_75t_SL g214335 (.A1(n_2996),
    .A2(n_1653),
    .B(n_3938),
    .C(n_2183),
    .Y(n_6030));
 O2A1O1Ixp33_ASAP7_75t_R g214336 (.A1(n_2468),
    .A2(n_1711),
    .B(n_1572),
    .C(sa00[0]),
    .Y(n_6029));
 O2A1O1Ixp33_ASAP7_75t_R g214337 (.A1(n_2449),
    .A2(n_2783),
    .B(n_2090),
    .C(n_1980),
    .Y(n_6028));
 OAI321xp33_ASAP7_75t_L g214338 (.A1(n_2175),
    .A2(n_1403),
    .A3(sa13[7]),
    .B1(n_1518),
    .B2(n_2874),
    .C(n_1429),
    .Y(n_6027));
 AOI31xp33_ASAP7_75t_R g214339 (.A1(n_2777),
    .A2(n_1748),
    .A3(n_1367),
    .B(n_3613),
    .Y(n_6026));
 OAI31xp33_ASAP7_75t_R g214340 (.A1(n_2780),
    .A2(n_1716),
    .A3(n_1845),
    .B(n_3690),
    .Y(n_6025));
 OAI21xp33_ASAP7_75t_R g214341 (.A1(n_1567),
    .A2(n_4352),
    .B(n_3401),
    .Y(n_6024));
 OAI211xp5_ASAP7_75t_R g214342 (.A1(n_1637),
    .A2(n_3083),
    .B(n_3933),
    .C(n_2152),
    .Y(n_6023));
 A2O1A1Ixp33_ASAP7_75t_L g214343 (.A1(n_1735),
    .A2(n_3528),
    .B(n_1418),
    .C(n_5325),
    .Y(n_6022));
 AOI211xp5_ASAP7_75t_L g214344 (.A1(n_3176),
    .A2(n_1641),
    .B(n_3941),
    .C(n_2188),
    .Y(n_6021));
 OAI21xp33_ASAP7_75t_SL g214345 (.A1(n_2066),
    .A2(n_4042),
    .B(n_2676),
    .Y(n_6020));
 AOI211xp5_ASAP7_75t_L g214346 (.A1(n_2944),
    .A2(n_1554),
    .B(n_3951),
    .C(n_2276),
    .Y(n_6019));
 AOI221xp5_ASAP7_75t_L g214347 (.A1(n_3084),
    .A2(n_1463),
    .B1(n_1638),
    .B2(n_2223),
    .C(n_5513),
    .Y(n_6018));
 AOI211xp5_ASAP7_75t_L g214348 (.A1(n_3027),
    .A2(n_2429),
    .B(n_3930),
    .C(n_2190),
    .Y(n_6017));
 OAI31xp33_ASAP7_75t_R g214349 (.A1(n_3252),
    .A2(n_3342),
    .A3(n_1844),
    .B(n_3625),
    .Y(n_6016));
 OAI21xp33_ASAP7_75t_L g214350 (.A1(n_2080),
    .A2(n_3250),
    .B(n_5427),
    .Y(n_6015));
 AOI211xp5_ASAP7_75t_R g214351 (.A1(n_3198),
    .A2(n_2051),
    .B(n_1768),
    .C(n_2250),
    .Y(n_6014));
 AOI22xp5_ASAP7_75t_L g214352 (.A1(n_1641),
    .A2(n_4362),
    .B1(n_2042),
    .B2(n_4648),
    .Y(n_6013));
 OAI321xp33_ASAP7_75t_L g214353 (.A1(n_2143),
    .A2(n_1501),
    .A3(sa21[7]),
    .B1(n_1975),
    .B2(n_2885),
    .C(n_1629),
    .Y(n_6012));
 O2A1O1Ixp33_ASAP7_75t_R g214354 (.A1(n_2451),
    .A2(n_3250),
    .B(n_1586),
    .C(n_1966),
    .Y(n_6011));
 A2O1A1Ixp33_ASAP7_75t_R g214355 (.A1(n_2439),
    .A2(n_2803),
    .B(n_2074),
    .C(n_1857),
    .Y(n_6010));
 AOI221xp5_ASAP7_75t_L g214356 (.A1(n_2935),
    .A2(n_2425),
    .B1(n_1545),
    .B2(n_2574),
    .C(n_3002),
    .Y(n_6009));
 OAI21xp33_ASAP7_75t_R g214357 (.A1(n_1373),
    .A2(n_1732),
    .B(n_5435),
    .Y(n_6008));
 OAI321xp33_ASAP7_75t_L g214358 (.A1(n_2129),
    .A2(n_1457),
    .A3(sa02[7]),
    .B1(n_8210),
    .B2(n_3433),
    .C(n_1389),
    .Y(n_6007));
 AO21x1_ASAP7_75t_R g214359 (.A1(n_3141),
    .A2(n_4317),
    .B(n_1664),
    .Y(n_6006));
 OAI21xp33_ASAP7_75t_SL g214360 (.A1(n_1392),
    .A2(n_3242),
    .B(n_5439),
    .Y(n_6005));
 OAI211xp5_ASAP7_75t_L g214361 (.A1(n_2070),
    .A2(n_2814),
    .B(n_5440),
    .C(n_3195),
    .Y(n_6004));
 A2O1A1Ixp33_ASAP7_75t_R g214362 (.A1(n_1387),
    .A2(n_1657),
    .B(n_3859),
    .C(n_2841),
    .Y(n_6003));
 OAI22xp33_ASAP7_75t_R g214363 (.A1(n_1383),
    .A2(n_4622),
    .B1(n_2074),
    .B2(n_3986),
    .Y(n_6002));
 OAI31xp33_ASAP7_75t_R g214364 (.A1(n_2891),
    .A2(n_3373),
    .A3(n_2088),
    .B(n_3343),
    .Y(n_6001));
 OAI21xp33_ASAP7_75t_L g214365 (.A1(n_4058),
    .A2(n_1628),
    .B(n_5509),
    .Y(n_6000));
 OAI321xp33_ASAP7_75t_R g214366 (.A1(n_2141),
    .A2(n_1844),
    .A3(n_1536),
    .B1(n_1985),
    .B2(n_3424),
    .C(n_2396),
    .Y(n_5999));
 OA21x2_ASAP7_75t_R g214367 (.A1(n_2437),
    .A2(n_4356),
    .B(n_1664),
    .Y(n_5998));
 A2O1A1Ixp33_ASAP7_75t_R g214368 (.A1(n_2833),
    .A2(n_2827),
    .B(n_1543),
    .C(n_4020),
    .Y(n_5997));
 AOI21xp33_ASAP7_75t_R g214369 (.A1(n_4311),
    .A2(n_1717),
    .B(n_1571),
    .Y(n_5996));
 OAI221xp5_ASAP7_75t_R g214370 (.A1(n_2929),
    .A2(n_1646),
    .B1(n_2061),
    .B2(n_2570),
    .C(n_3011),
    .Y(n_5995));
 OAI31xp33_ASAP7_75t_R g214371 (.A1(n_1742),
    .A2(n_2879),
    .A3(n_1573),
    .B(n_3376),
    .Y(n_5994));
 AOI31xp33_ASAP7_75t_R g214372 (.A1(n_3331),
    .A2(n_2875),
    .A3(n_1586),
    .B(n_3389),
    .Y(n_5993));
 O2A1O1Ixp33_ASAP7_75t_R g214373 (.A1(n_2488),
    .A2(n_2430),
    .B(n_4075),
    .C(n_2372),
    .Y(n_5992));
 OAI31xp33_ASAP7_75t_L g214374 (.A1(n_3846),
    .A2(n_2476),
    .A3(n_1500),
    .B(n_1376),
    .Y(n_5991));
 OAI21xp33_ASAP7_75t_L g214375 (.A1(n_2829),
    .A2(n_3008),
    .B(n_5522),
    .Y(n_5990));
 OAI21xp33_ASAP7_75t_R g214376 (.A1(n_1714),
    .A2(n_4315),
    .B(n_2389),
    .Y(n_5989));
 AOI211xp5_ASAP7_75t_SL g214377 (.A1(n_2954),
    .A2(n_1581),
    .B(n_5021),
    .C(n_2582),
    .Y(n_5988));
 O2A1O1Ixp33_ASAP7_75t_L g214378 (.A1(n_2478),
    .A2(n_2789),
    .B(n_2079),
    .C(n_4978),
    .Y(n_5987));
 OAI31xp33_ASAP7_75t_R g214379 (.A1(n_3261),
    .A2(n_3313),
    .A3(n_2372),
    .B(n_8180),
    .Y(n_5986));
 AOI211xp5_ASAP7_75t_SL g214380 (.A1(n_3056),
    .A2(n_2079),
    .B(n_4966),
    .C(n_2628),
    .Y(n_5985));
 OAI21xp33_ASAP7_75t_R g214381 (.A1(n_2606),
    .A2(n_4290),
    .B(n_1667),
    .Y(n_5984));
 AOI31xp33_ASAP7_75t_R g214382 (.A1(n_2878),
    .A2(n_1577),
    .A3(n_1741),
    .B(n_3391),
    .Y(n_5983));
 AOI22xp33_ASAP7_75t_R g214383 (.A1(n_4573),
    .A2(n_1633),
    .B1(n_4006),
    .B2(n_2084),
    .Y(n_5982));
 NOR3xp33_ASAP7_75t_L g214384 (.A(n_5428),
    .B(n_4199),
    .C(n_8188),
    .Y(n_5981));
 AOI31xp33_ASAP7_75t_R g214385 (.A1(n_2827),
    .A2(n_2833),
    .A3(n_1446),
    .B(n_4536),
    .Y(n_5980));
 A2O1A1Ixp33_ASAP7_75t_R g214386 (.A1(n_2495),
    .A2(n_1348),
    .B(n_4179),
    .C(n_1621),
    .Y(n_5979));
 OAI221xp5_ASAP7_75t_L g214387 (.A1(n_3776),
    .A2(n_1551),
    .B1(n_1337),
    .B2(n_3288),
    .C(n_3781),
    .Y(n_5978));
 AOI21xp33_ASAP7_75t_R g214388 (.A1(n_3258),
    .A2(n_4300),
    .B(n_1429),
    .Y(n_6233));
 OAI21xp33_ASAP7_75t_R g214389 (.A1(n_3244),
    .A2(n_4292),
    .B(n_8690),
    .Y(n_5977));
 NOR2xp33_ASAP7_75t_L g214390 (.A(n_5309),
    .B(n_3926),
    .Y(n_5976));
 OA21x2_ASAP7_75t_SL g214391 (.A1(n_1344),
    .A2(n_3987),
    .B(n_5441),
    .Y(n_5975));
 AOI221xp5_ASAP7_75t_L g214392 (.A1(n_1406),
    .A2(n_3465),
    .B1(n_2757),
    .B2(n_2055),
    .C(n_1698),
    .Y(n_5974));
 AOI22xp33_ASAP7_75t_L g214393 (.A1(n_1622),
    .A2(n_4568),
    .B1(n_2079),
    .B2(n_3850),
    .Y(n_5973));
 OAI221xp5_ASAP7_75t_L g214394 (.A1(n_2936),
    .A2(n_1382),
    .B1(n_1354),
    .B2(n_3094),
    .C(n_4977),
    .Y(n_5972));
 OAI21xp33_ASAP7_75t_R g214395 (.A1(n_3248),
    .A2(n_4296),
    .B(n_1422),
    .Y(n_5971));
 OR3x1_ASAP7_75t_L g214396 (.A(n_3918),
    .B(n_4272),
    .C(n_3577),
    .Y(n_5970));
 OAI21xp33_ASAP7_75t_R g214397 (.A1(n_4288),
    .A2(n_2804),
    .B(n_1659),
    .Y(n_5969));
 OAI21xp33_ASAP7_75t_R g214398 (.A1(n_2866),
    .A2(n_4332),
    .B(n_2089),
    .Y(n_5968));
 OAI21xp33_ASAP7_75t_R g214399 (.A1(n_2780),
    .A2(n_4327),
    .B(n_1652),
    .Y(n_5967));
 OAI21xp33_ASAP7_75t_L g214400 (.A1(n_2347),
    .A2(n_3909),
    .B(n_1500),
    .Y(n_5966));
 AOI21xp5_ASAP7_75t_SL g214401 (.A1(n_3857),
    .A2(n_1356),
    .B(n_5442),
    .Y(n_5965));
 AOI21xp33_ASAP7_75t_R g214402 (.A1(n_4281),
    .A2(n_2618),
    .B(n_2434),
    .Y(n_5964));
 NAND2xp33_ASAP7_75t_L g214403 (.A(n_4837),
    .B(n_5017),
    .Y(n_5963));
 AO21x1_ASAP7_75t_R g214404 (.A1(n_2442),
    .A2(n_4338),
    .B(n_1669),
    .Y(n_5962));
 AOI21xp33_ASAP7_75t_R g214405 (.A1(n_4294),
    .A2(n_1693),
    .B(n_1647),
    .Y(n_5961));
 OAI21xp5_ASAP7_75t_L g214406 (.A1(n_3296),
    .A2(n_3146),
    .B(n_5524),
    .Y(n_5960));
 AOI31xp33_ASAP7_75t_R g214407 (.A1(n_4295),
    .A2(n_2439),
    .A3(n_1457),
    .B(n_2435),
    .Y(n_5959));
 O2A1O1Ixp33_ASAP7_75t_R g214408 (.A1(n_8189),
    .A2(n_1647),
    .B(n_3905),
    .C(n_2839),
    .Y(n_5958));
 OAI31xp33_ASAP7_75t_L g214409 (.A1(n_1714),
    .A2(n_2830),
    .A3(n_2358),
    .B(n_1464),
    .Y(n_5957));
 OAI31xp33_ASAP7_75t_R g214410 (.A1(n_2780),
    .A2(n_2838),
    .A3(n_2356),
    .B(n_1845),
    .Y(n_5956));
 OAI21xp5_ASAP7_75t_SL g214411 (.A1(n_2358),
    .A2(n_3862),
    .B(n_1463),
    .Y(n_6232));
 AOI31xp33_ASAP7_75t_R g214412 (.A1(n_2805),
    .A2(n_2843),
    .A3(n_2367),
    .B(sa11[6]),
    .Y(n_5955));
 AOI31xp33_ASAP7_75t_L g214413 (.A1(n_4287),
    .A2(n_2473),
    .A3(n_1850),
    .B(n_1655),
    .Y(n_5954));
 AOI31xp33_ASAP7_75t_L g214414 (.A1(n_3844),
    .A2(n_2456),
    .A3(n_1496),
    .B(n_2065),
    .Y(n_5953));
 OAI211xp5_ASAP7_75t_L g214415 (.A1(n_1654),
    .A2(n_3092),
    .B(n_3939),
    .C(n_2184),
    .Y(n_5952));
 O2A1O1Ixp33_ASAP7_75t_R g214416 (.A1(n_1502),
    .A2(n_2424),
    .B(n_3914),
    .C(n_2834),
    .Y(n_5951));
 AOI21xp33_ASAP7_75t_R g214417 (.A1(n_3884),
    .A2(n_2364),
    .B(n_1459),
    .Y(n_5950));
 OAI321xp33_ASAP7_75t_R g214418 (.A1(n_2550),
    .A2(n_1674),
    .A3(n_1518),
    .B1(n_1519),
    .B2(n_3310),
    .C(n_1403),
    .Y(n_5949));
 AO21x1_ASAP7_75t_R g214419 (.A1(n_2370),
    .A2(n_4355),
    .B(n_1456),
    .Y(n_5948));
 AOI31xp33_ASAP7_75t_R g214420 (.A1(n_2788),
    .A2(n_2849),
    .A3(n_2354),
    .B(n_1346),
    .Y(n_5947));
 AOI31xp33_ASAP7_75t_R g214421 (.A1(n_3287),
    .A2(n_3425),
    .A3(n_2360),
    .B(n_1499),
    .Y(n_5946));
 AOI31xp33_ASAP7_75t_R g214422 (.A1(n_2800),
    .A2(n_2847),
    .A3(n_2366),
    .B(n_1497),
    .Y(n_5945));
 OAI31xp33_ASAP7_75t_R g214423 (.A1(n_2806),
    .A2(n_2858),
    .A3(n_2351),
    .B(n_1397),
    .Y(n_5944));
 NOR3xp33_ASAP7_75t_L g214424 (.A(n_4868),
    .B(n_3819),
    .C(n_2541),
    .Y(n_5943));
 A2O1A1Ixp33_ASAP7_75t_SL g214425 (.A1(n_2843),
    .A2(n_3268),
    .B(n_1450),
    .C(n_4912),
    .Y(n_5942));
 OAI31xp33_ASAP7_75t_L g214426 (.A1(n_4327),
    .A2(n_2468),
    .A3(n_1461),
    .B(n_2411),
    .Y(n_5941));
 OAI31xp33_ASAP7_75t_R g214427 (.A1(n_1776),
    .A2(n_2441),
    .A3(n_1395),
    .B(n_2428),
    .Y(n_5940));
 OAI31xp33_ASAP7_75t_SL g214428 (.A1(n_3245),
    .A2(n_3366),
    .A3(n_1408),
    .B(n_4939),
    .Y(n_5939));
 OAI21xp5_ASAP7_75t_R g214429 (.A1(n_2468),
    .A2(n_4344),
    .B(n_2410),
    .Y(n_5938));
 AOI31xp33_ASAP7_75t_R g214430 (.A1(n_4326),
    .A2(n_2448),
    .A3(n_1499),
    .B(n_1348),
    .Y(n_5937));
 AOI221xp5_ASAP7_75t_L g214431 (.A1(n_3446),
    .A2(n_2427),
    .B1(n_2054),
    .B2(n_2547),
    .C(n_3005),
    .Y(n_5936));
 OA21x2_ASAP7_75t_L g214432 (.A1(n_1590),
    .A2(n_3856),
    .B(n_5076),
    .Y(n_5935));
 OAI21xp33_ASAP7_75t_R g214433 (.A1(n_3263),
    .A2(n_4292),
    .B(n_2414),
    .Y(n_5934));
 AOI31xp33_ASAP7_75t_R g214434 (.A1(n_4286),
    .A2(n_2477),
    .A3(n_1938),
    .B(n_1622),
    .Y(n_5933));
 AOI21xp33_ASAP7_75t_R g214435 (.A1(n_4287),
    .A2(n_3268),
    .B(n_1656),
    .Y(n_5932));
 AOI21xp33_ASAP7_75t_R g214436 (.A1(n_2488),
    .A2(n_4357),
    .B(n_2041),
    .Y(n_5931));
 AOI31xp33_ASAP7_75t_R g214437 (.A1(n_1777),
    .A2(n_2485),
    .A3(n_1397),
    .B(n_2387),
    .Y(n_5930));
 AOI211xp5_ASAP7_75t_L g214438 (.A1(n_2226),
    .A2(n_2429),
    .B(n_5090),
    .C(n_3269),
    .Y(n_5929));
 OAI21xp33_ASAP7_75t_R g214439 (.A1(n_2081),
    .A2(n_2782),
    .B(n_5077),
    .Y(n_5928));
 OAI31xp33_ASAP7_75t_R g214440 (.A1(n_4297),
    .A2(n_2484),
    .A3(n_1346),
    .B(n_1647),
    .Y(n_5927));
 A2O1A1Ixp33_ASAP7_75t_R g214441 (.A1(n_2551),
    .A2(n_2777),
    .B(n_1624),
    .C(n_4012),
    .Y(n_5926));
 AOI211xp5_ASAP7_75t_L g214442 (.A1(n_1445),
    .A2(n_3670),
    .B(n_3956),
    .C(n_3684),
    .Y(n_5925));
 AOI31xp33_ASAP7_75t_SL g214443 (.A1(n_3258),
    .A2(n_2828),
    .A3(n_2392),
    .B(n_4701),
    .Y(n_5924));
 O2A1O1Ixp33_ASAP7_75t_R g214444 (.A1(n_2560),
    .A2(n_2806),
    .B(n_2387),
    .C(n_4015),
    .Y(n_5923));
 OAI321xp33_ASAP7_75t_R g214445 (.A1(n_2441),
    .A2(n_2501),
    .A3(n_1844),
    .B1(n_2141),
    .B2(n_1443),
    .C(n_5511),
    .Y(n_5922));
 AOI221xp5_ASAP7_75t_R g214446 (.A1(n_8719),
    .A2(n_2196),
    .B1(n_4706),
    .B2(n_2064),
    .C(n_3263),
    .Y(n_5921));
 AOI21xp33_ASAP7_75t_R g214447 (.A1(n_2796),
    .A2(n_3844),
    .B(n_2066),
    .Y(n_5920));
 AOI21xp5_ASAP7_75t_SL g214448 (.A1(n_4026),
    .A2(n_1441),
    .B(n_5088),
    .Y(n_5919));
 OAI21xp33_ASAP7_75t_L g214449 (.A1(n_1380),
    .A2(n_1767),
    .B(n_5078),
    .Y(n_5918));
 AOI211xp5_ASAP7_75t_L g214450 (.A1(n_1451),
    .A2(n_2275),
    .B(n_5079),
    .C(n_2818),
    .Y(n_5917));
 OAI21xp33_ASAP7_75t_R g214451 (.A1(n_2495),
    .A2(n_4379),
    .B(n_1561),
    .Y(n_5916));
 AOI21xp33_ASAP7_75t_R g214452 (.A1(n_3370),
    .A2(n_4284),
    .B(n_1443),
    .Y(n_5915));
 OAI22xp33_ASAP7_75t_R g214453 (.A1(n_1845),
    .A2(n_3827),
    .B1(n_2585),
    .B2(n_2419),
    .Y(n_5914));
 AO21x1_ASAP7_75t_L g214454 (.A1(n_1561),
    .A2(n_3997),
    .B(n_5084),
    .Y(n_5913));
 OA21x2_ASAP7_75t_L g214455 (.A1(n_2047),
    .A2(n_3984),
    .B(n_5087),
    .Y(n_5912));
 AOI221xp5_ASAP7_75t_L g214456 (.A1(n_3077),
    .A2(n_2895),
    .B1(n_2984),
    .B2(n_1707),
    .C(n_4899),
    .Y(n_5911));
 OAI21xp33_ASAP7_75t_SL g214457 (.A1(n_1369),
    .A2(n_3961),
    .B(n_5093),
    .Y(n_5910));
 OAI21xp33_ASAP7_75t_L g214458 (.A1(n_1546),
    .A2(n_3949),
    .B(n_5083),
    .Y(n_5909));
 OAI21xp33_ASAP7_75t_L g214459 (.A1(n_2045),
    .A2(n_3944),
    .B(n_5089),
    .Y(n_5908));
 AO21x1_ASAP7_75t_L g214460 (.A1(n_1449),
    .A2(n_4027),
    .B(n_5085),
    .Y(n_5907));
 OAI31xp33_ASAP7_75t_L g214461 (.A1(n_2801),
    .A2(n_2066),
    .A3(n_2326),
    .B(n_5487),
    .Y(n_5906));
 OAI32xp33_ASAP7_75t_L g214462 (.A1(n_3252),
    .A2(n_2428),
    .A3(n_2294),
    .B1(n_1354),
    .B2(n_3852),
    .Y(n_5905));
 OAI21xp33_ASAP7_75t_R g214463 (.A1(n_3174),
    .A2(n_1711),
    .B(n_5091),
    .Y(n_5904));
 OAI221xp5_ASAP7_75t_SL g214464 (.A1(n_3054),
    .A2(n_1666),
    .B1(n_1637),
    .B2(n_2959),
    .C(n_4754),
    .Y(n_5903));
 AOI22xp33_ASAP7_75t_L g214465 (.A1(n_2494),
    .A2(n_3825),
    .B1(n_2205),
    .B2(n_1566),
    .Y(n_5902));
 A2O1A1Ixp33_ASAP7_75t_L g214466 (.A1(n_2442),
    .A2(n_1712),
    .B(n_1590),
    .C(n_5503),
    .Y(n_5901));
 AOI211xp5_ASAP7_75t_L g214467 (.A1(n_2042),
    .A2(n_2621),
    .B(n_4764),
    .C(n_4089),
    .Y(n_5900));
 A2O1A1Ixp33_ASAP7_75t_SL g214468 (.A1(n_2456),
    .A2(n_1731),
    .B(n_2088),
    .C(n_5501),
    .Y(n_5899));
 OAI31xp33_ASAP7_75t_R g214469 (.A1(n_4315),
    .A2(n_2443),
    .A3(n_1463),
    .B(n_1666),
    .Y(n_5898));
 OAI221xp5_ASAP7_75t_SL g214470 (.A1(n_1644),
    .A2(n_2955),
    .B1(n_1392),
    .B2(n_3214),
    .C(n_4877),
    .Y(n_5897));
 OAI21xp33_ASAP7_75t_R g214471 (.A1(n_3846),
    .A2(n_2786),
    .B(n_1350),
    .Y(n_5896));
 AOI21xp33_ASAP7_75t_R g214472 (.A1(n_2907),
    .A2(n_4277),
    .B(n_1344),
    .Y(n_5895));
 OAI31xp33_ASAP7_75t_R g214473 (.A1(n_4292),
    .A2(n_2482),
    .A3(n_1455),
    .B(n_1651),
    .Y(n_5894));
 OAI321xp33_ASAP7_75t_L g214474 (.A1(n_2059),
    .A2(n_2177),
    .A3(n_1473),
    .B1(n_2423),
    .B2(n_1725),
    .C(n_4990),
    .Y(n_5893));
 AOI221xp5_ASAP7_75t_L g214475 (.A1(n_2064),
    .A2(n_3068),
    .B1(n_2077),
    .B2(n_2281),
    .C(n_5008),
    .Y(n_5892));
 OAI31xp33_ASAP7_75t_R g214476 (.A1(n_4299),
    .A2(n_2451),
    .A3(n_1934),
    .B(n_2422),
    .Y(n_5891));
 OAI221xp5_ASAP7_75t_R g214477 (.A1(n_1725),
    .A2(n_2393),
    .B1(n_1584),
    .B2(n_3604),
    .C(n_5022),
    .Y(n_5890));
 OAI221xp5_ASAP7_75t_L g214478 (.A1(n_3058),
    .A2(n_2419),
    .B1(n_1571),
    .B2(n_1612),
    .C(n_4734),
    .Y(n_5889));
 OAI21xp33_ASAP7_75t_R g214479 (.A1(n_2465),
    .A2(n_4282),
    .B(n_2067),
    .Y(n_6230));
 AOI21xp5_ASAP7_75t_R g214480 (.A1(n_4277),
    .A2(n_2471),
    .B(n_1450),
    .Y(n_6229));
 OAI21xp5_ASAP7_75t_R g214481 (.A1(n_1678),
    .A2(n_4309),
    .B(n_1542),
    .Y(n_6228));
 NOR2xp33_ASAP7_75t_L g214482 (.A(n_2059),
    .B(n_5534),
    .Y(n_5888));
 AOI21xp5_ASAP7_75t_R g214483 (.A1(n_4301),
    .A2(n_2462),
    .B(n_1582),
    .Y(n_6227));
 OAI21xp5_ASAP7_75t_L g214484 (.A1(n_1679),
    .A2(n_4293),
    .B(n_2062),
    .Y(n_6225));
 AOI21xp33_ASAP7_75t_R g214485 (.A1(n_1673),
    .A2(n_4307),
    .B(n_2043),
    .Y(n_6224));
 OAI21xp5_ASAP7_75t_R g214486 (.A1(n_4279),
    .A2(n_2495),
    .B(n_1559),
    .Y(n_6223));
 AOI21xp5_ASAP7_75t_R g214487 (.A1(n_4289),
    .A2(n_1670),
    .B(n_2057),
    .Y(n_6222));
 AOI21xp5_ASAP7_75t_R g214488 (.A1(n_2444),
    .A2(n_4331),
    .B(n_2047),
    .Y(n_6220));
 AOI21xp33_ASAP7_75t_R g214489 (.A1(n_4319),
    .A2(n_1682),
    .B(n_1546),
    .Y(n_6219));
 OAI21xp33_ASAP7_75t_L g214490 (.A1(n_2492),
    .A2(n_4283),
    .B(n_1440),
    .Y(n_6217));
 AO21x1_ASAP7_75t_L g214491 (.A1(n_2488),
    .A2(n_4323),
    .B(n_2041),
    .Y(n_6216));
 NAND2xp33_ASAP7_75t_R g214492 (.A(n_1416),
    .B(n_5535),
    .Y(n_5887));
 AND3x1_ASAP7_75t_R g214493 (.A(n_3987),
    .B(n_1850),
    .C(sa11[3]),
    .Y(n_6215));
 NAND2xp5_ASAP7_75t_L g214494 (.A(n_1933),
    .B(n_5388),
    .Y(n_6214));
 NAND2xp5_ASAP7_75t_R g214495 (.A(n_1460),
    .B(n_5386),
    .Y(n_6213));
 NAND2xp5_ASAP7_75t_R g214496 (.A(n_1839),
    .B(n_5396),
    .Y(n_6212));
 NAND2xp5_ASAP7_75t_L g214497 (.A(n_8180),
    .B(n_5047),
    .Y(n_6210));
 NOR2xp33_ASAP7_75t_R g214498 (.A(n_1455),
    .B(n_5403),
    .Y(n_6209));
 NAND2xp5_ASAP7_75t_SL g214499 (.A(n_1348),
    .B(n_5377),
    .Y(n_6208));
 NOR2xp33_ASAP7_75t_R g214500 (.A(n_2428),
    .B(n_5393),
    .Y(n_6207));
 NOR2xp33_ASAP7_75t_R g214501 (.A(n_1408),
    .B(n_5378),
    .Y(n_5886));
 AND2x2_ASAP7_75t_SL g214502 (.A(n_1404),
    .B(n_5397),
    .Y(n_6206));
 NAND2xp33_ASAP7_75t_L g214503 (.A(n_2386),
    .B(n_5379),
    .Y(n_6205));
 NAND2xp5_ASAP7_75t_R g214504 (.A(n_1459),
    .B(n_5398),
    .Y(n_6203));
 AND2x2_ASAP7_75t_L g214505 (.A(n_1419),
    .B(n_5437),
    .Y(n_6202));
 NOR2xp33_ASAP7_75t_R g214506 (.A(n_2424),
    .B(n_5383),
    .Y(n_5885));
 NOR2xp33_ASAP7_75t_L g214507 (.A(n_1544),
    .B(n_5430),
    .Y(n_5884));
 NOR2xp33_ASAP7_75t_L g214508 (.A(n_2047),
    .B(n_5422),
    .Y(n_6201));
 NOR2xp33_ASAP7_75t_L g214510 (.A(n_1450),
    .B(n_5418),
    .Y(n_5882));
 NAND2xp5_ASAP7_75t_L g214511 (.A(sa31[6]),
    .B(n_5388),
    .Y(n_6200));
 OAI211xp5_ASAP7_75t_R g214512 (.A1(n_8899),
    .A2(n_2783),
    .B(n_1559),
    .C(n_2448),
    .Y(n_1797));
 NOR2xp33_ASAP7_75t_L g214513 (.A(n_1850),
    .B(n_5405),
    .Y(n_6198));
 OAI211xp5_ASAP7_75t_R g214514 (.A1(sa22[4]),
    .A2(n_2782),
    .B(n_2054),
    .C(n_2440),
    .Y(n_6197));
 NAND2xp33_ASAP7_75t_L g214515 (.A(n_2077),
    .B(n_5445),
    .Y(n_1796));
 NOR2xp33_ASAP7_75t_SL g214516 (.A(n_1845),
    .B(n_5387),
    .Y(n_5881));
 NAND2xp33_ASAP7_75t_R g214517 (.A(n_1346),
    .B(n_5396),
    .Y(n_5880));
 NAND2xp5_ASAP7_75t_L g214518 (.A(n_1444),
    .B(n_5406),
    .Y(n_6195));
 AND2x2_ASAP7_75t_SL g214519 (.A(n_1455),
    .B(n_5404),
    .Y(n_6194));
 AOI211xp5_ASAP7_75t_L g214520 (.A1(n_3251),
    .A2(n_1505),
    .B(n_2059),
    .C(n_2451),
    .Y(n_6193));
 NAND2xp5_ASAP7_75t_L g214521 (.A(n_5397),
    .B(n_1934),
    .Y(n_6191));
 NOR2xp67_ASAP7_75t_L g214522 (.A(n_1457),
    .B(n_5399),
    .Y(n_6190));
 NOR2xp33_ASAP7_75t_R g214523 (.A(n_1371),
    .B(n_5048),
    .Y(n_6189));
 NAND2xp5_ASAP7_75t_L g214524 (.A(n_5507),
    .B(n_1451),
    .Y(n_6187));
 OAI21xp5_ASAP7_75t_L g214525 (.A1(n_4315),
    .A2(n_4290),
    .B(n_2389),
    .Y(n_6185));
 OAI21xp5_ASAP7_75t_SL g214526 (.A1(n_4302),
    .A2(n_4292),
    .B(n_8690),
    .Y(n_1795));
 NOR2xp33_ASAP7_75t_L g214527 (.A(n_1429),
    .B(n_5473),
    .Y(n_5879));
 OAI21xp5_ASAP7_75t_SL g214528 (.A1(n_4296),
    .A2(n_4282),
    .B(n_2400),
    .Y(n_6183));
 AOI21xp5_ASAP7_75t_L g214529 (.A1(n_4277),
    .A2(n_4287),
    .B(n_1660),
    .Y(n_6182));
 OAI21xp5_ASAP7_75t_SL g214530 (.A1(n_3846),
    .A2(n_4309),
    .B(n_1627),
    .Y(n_6180));
 OAI21xp5_ASAP7_75t_L g214531 (.A1(n_3845),
    .A2(n_4332),
    .B(n_1554),
    .Y(n_6177));
 NAND2xp5_ASAP7_75t_SL g214532 (.A(n_5527),
    .B(n_2397),
    .Y(n_6176));
 NAND2xp5_ASAP7_75t_SL g214533 (.A(n_1566),
    .B(n_5526),
    .Y(n_6174));
 NAND2xp5_ASAP7_75t_L g214534 (.A(n_1793),
    .B(n_1653),
    .Y(n_6173));
 AND2x2_ASAP7_75t_L g214535 (.A(n_2398),
    .B(n_5521),
    .Y(n_6172));
 AOI21xp5_ASAP7_75t_R g214536 (.A1(n_4307),
    .A2(n_4286),
    .B(n_1640),
    .Y(n_6171));
 OAI21xp5_ASAP7_75t_L g214537 (.A1(n_4322),
    .A2(n_4316),
    .B(n_1449),
    .Y(n_6170));
 INVxp67_ASAP7_75t_R g214538 (.A(n_5794),
    .Y(n_5878));
 INVxp67_ASAP7_75t_R g214539 (.A(n_5737),
    .Y(n_5877));
 AOI211xp5_ASAP7_75t_L g214540 (.A1(n_1449),
    .A2(n_2505),
    .B(n_4957),
    .C(n_3789),
    .Y(n_5876));
 OAI22xp33_ASAP7_75t_R g214541 (.A1(n_2041),
    .A2(n_4229),
    .B1(n_2594),
    .B2(n_2395),
    .Y(n_5875));
 A2O1A1Ixp33_ASAP7_75t_R g214542 (.A1(n_2488),
    .A2(n_2110),
    .B(n_1363),
    .C(n_4873),
    .Y(n_5874));
 OAI21xp33_ASAP7_75t_L g214543 (.A1(n_2428),
    .A2(n_4026),
    .B(n_5303),
    .Y(n_5873));
 OAI22xp33_ASAP7_75t_R g214544 (.A1(n_2053),
    .A2(n_4238),
    .B1(n_2428),
    .B2(n_4284),
    .Y(n_5872));
 OAI22xp33_ASAP7_75t_R g214545 (.A1(n_4225),
    .A2(n_2441),
    .B1(n_1413),
    .B2(n_2440),
    .Y(n_5871));
 OAI22xp33_ASAP7_75t_R g214546 (.A1(n_4227),
    .A2(n_2449),
    .B1(n_2448),
    .B2(n_1348),
    .Y(n_5870));
 OAI221xp5_ASAP7_75t_L g214547 (.A1(n_2396),
    .A2(n_3438),
    .B1(n_2053),
    .B2(n_1704),
    .C(n_5031),
    .Y(n_5869));
 OAI22xp33_ASAP7_75t_R g214548 (.A1(n_2457),
    .A2(n_4226),
    .B1(n_2065),
    .B2(n_2456),
    .Y(n_5868));
 O2A1O1Ixp33_ASAP7_75t_R g214549 (.A1(n_2158),
    .A2(n_3421),
    .B(n_1343),
    .C(n_3753),
    .Y(n_5867));
 O2A1O1Ixp33_ASAP7_75t_R g214550 (.A1(n_2131),
    .A2(n_2891),
    .B(sa03[3]),
    .C(n_3751),
    .Y(n_5866));
 AOI22xp33_ASAP7_75t_R g214551 (.A1(sa03[3]),
    .A2(n_3849),
    .B1(n_1558),
    .B2(n_4230),
    .Y(n_5865));
 A2O1A1Ixp33_ASAP7_75t_R g214552 (.A1(n_1577),
    .A2(n_3189),
    .B(n_2484),
    .C(n_2752),
    .Y(n_5864));
 OAI221xp5_ASAP7_75t_R g214553 (.A1(n_2789),
    .A2(n_8177),
    .B1(n_2943),
    .B2(n_1367),
    .C(n_3836),
    .Y(n_5863));
 AOI221xp5_ASAP7_75t_SL g214554 (.A1(n_2922),
    .A2(n_1501),
    .B1(n_2816),
    .B2(sa21[3]),
    .C(n_3838),
    .Y(n_5862));
 AO221x1_ASAP7_75t_SL g214555 (.A1(n_3241),
    .A2(n_1984),
    .B1(n_3531),
    .B2(n_1933),
    .C(n_3837),
    .Y(n_5861));
 AOI222xp33_ASAP7_75t_L g214556 (.A1(n_3603),
    .A2(n_1518),
    .B1(n_1431),
    .B2(n_2175),
    .C1(n_3506),
    .C2(n_1404),
    .Y(n_5860));
 OAI221xp5_ASAP7_75t_L g214557 (.A1(n_3067),
    .A2(n_1512),
    .B1(n_1609),
    .B2(n_1583),
    .C(n_4263),
    .Y(n_5859));
 OAI222xp33_ASAP7_75t_R g214558 (.A1(n_2925),
    .A2(n_1346),
    .B1(n_3030),
    .B2(sa33[3]),
    .C1(n_2061),
    .C2(n_2127),
    .Y(n_5858));
 AOI222xp33_ASAP7_75t_R g214559 (.A1(n_2930),
    .A2(n_1459),
    .B1(n_3062),
    .B2(n_8210),
    .C1(n_2067),
    .C2(n_2129),
    .Y(n_5857));
 XNOR2xp5_ASAP7_75t_L g214561 (.A(n_4461),
    .B(n_1984),
    .Y(n_5856));
 AOI221xp5_ASAP7_75t_SL g214562 (.A1(n_3540),
    .A2(n_1555),
    .B1(n_1432),
    .B2(n_2131),
    .C(n_5182),
    .Y(n_5855));
 AOI222xp33_ASAP7_75t_L g214563 (.A1(n_2055),
    .A2(n_2589),
    .B1(n_2919),
    .B2(n_2410),
    .C1(n_2590),
    .C2(n_1653),
    .Y(n_5854));
 AOI21xp5_ASAP7_75t_L g214564 (.A1(n_4175),
    .A2(n_1577),
    .B(n_4789),
    .Y(n_5853));
 OAI22xp5_ASAP7_75t_L g214565 (.A1(sa03[3]),
    .A2(n_4594),
    .B1(n_1967),
    .B2(n_4595),
    .Y(n_5852));
 XNOR2xp5_ASAP7_75t_R g214566 (.A(n_3968),
    .B(sa33[3]),
    .Y(n_5851));
 OAI221xp5_ASAP7_75t_SL g214567 (.A1(n_4077),
    .A2(n_2083),
    .B1(n_1644),
    .B2(n_3586),
    .C(n_2772),
    .Y(n_5850));
 OAI22xp5_ASAP7_75t_SL g214568 (.A1(sa01[3]),
    .A2(n_3975),
    .B1(n_1859),
    .B2(n_3974),
    .Y(n_5849));
 AOI222xp33_ASAP7_75t_SL g214569 (.A1(n_3581),
    .A2(n_2429),
    .B1(n_1655),
    .B2(n_2187),
    .C1(n_4144),
    .C2(n_1576),
    .Y(n_5848));
 OAI221xp5_ASAP7_75t_L g214570 (.A1(n_4187),
    .A2(n_1381),
    .B1(n_1639),
    .B2(n_3719),
    .C(n_2769),
    .Y(n_5847));
 OAI222xp33_ASAP7_75t_L g214571 (.A1(n_4658),
    .A2(n_1418),
    .B1(n_1754),
    .B2(n_8691),
    .C1(n_1651),
    .C2(n_1609),
    .Y(n_5846));
 XOR2xp5_ASAP7_75t_L g214572 (.A(n_3733),
    .B(sa22[3]),
    .Y(n_5845));
 OAI22xp5_ASAP7_75t_SL g214573 (.A1(sa11[3]),
    .A2(n_3978),
    .B1(n_1986),
    .B2(n_3977),
    .Y(n_5844));
 AOI22xp33_ASAP7_75t_L g214574 (.A1(n_1467),
    .A2(n_3967),
    .B1(sa00[3]),
    .B2(n_3966),
    .Y(n_5843));
 OAI22xp33_ASAP7_75t_SL g214575 (.A1(n_1519),
    .A2(n_3948),
    .B1(n_1518),
    .B2(n_3947),
    .Y(n_5842));
 OAI22xp5_ASAP7_75t_L g214576 (.A1(n_1512),
    .A2(n_3980),
    .B1(n_1971),
    .B2(n_3981),
    .Y(n_5841));
 OAI221xp5_ASAP7_75t_SL g214577 (.A1(n_4538),
    .A2(n_2081),
    .B1(n_1442),
    .B2(n_3222),
    .C(n_2767),
    .Y(n_5840));
 OAI222xp33_ASAP7_75t_SL g214578 (.A1(n_3066),
    .A2(n_3511),
    .B1(n_3706),
    .B2(n_8702),
    .C1(n_1583),
    .C2(n_2575),
    .Y(n_5839));
 OAI222xp33_ASAP7_75t_SL g214579 (.A1(n_1543),
    .A2(n_3435),
    .B1(n_4533),
    .B2(n_1629),
    .C1(n_1376),
    .C2(n_2011),
    .Y(n_5838));
 AOI222xp33_ASAP7_75t_SL g214580 (.A1(n_1451),
    .A2(n_4482),
    .B1(n_2062),
    .B2(n_3490),
    .C1(n_2401),
    .C2(n_2014),
    .Y(n_5837));
 XOR2xp5_ASAP7_75t_L g214581 (.A(n_3732),
    .B(n_1343),
    .Y(n_5836));
 OAI211xp5_ASAP7_75t_SL g214582 (.A1(n_1580),
    .A2(n_3878),
    .B(n_4143),
    .C(n_4663),
    .Y(n_5835));
 AOI221xp5_ASAP7_75t_SL g214583 (.A1(n_3535),
    .A2(n_1433),
    .B1(n_1622),
    .B2(n_1484),
    .C(n_5147),
    .Y(n_5834));
 OAI221xp5_ASAP7_75t_L g214584 (.A1(n_3599),
    .A2(n_2395),
    .B1(n_1665),
    .B2(n_2100),
    .C(n_5202),
    .Y(n_5833));
 AOI221xp5_ASAP7_75t_L g214585 (.A1(n_4459),
    .A2(n_2429),
    .B1(n_1657),
    .B2(n_2015),
    .C(n_4256),
    .Y(n_5832));
 OAI21xp33_ASAP7_75t_L g214586 (.A1(n_1654),
    .A2(n_4487),
    .B(n_4811),
    .Y(n_5831));
 AOI222xp33_ASAP7_75t_R g214587 (.A1(n_1444),
    .A2(n_3488),
    .B1(n_1405),
    .B2(sa02[7]),
    .C1(n_4458),
    .C2(n_2400),
    .Y(n_5830));
 AOI222xp33_ASAP7_75t_SL g214588 (.A1(n_2040),
    .A2(n_3514),
    .B1(n_2387),
    .B2(n_1525),
    .C1(n_4512),
    .C2(n_2398),
    .Y(n_5829));
 OA222x2_ASAP7_75t_R g214589 (.A1(n_1582),
    .A2(n_3528),
    .B1(n_1651),
    .B2(n_2019),
    .C1(n_8702),
    .C2(n_4500),
    .Y(n_5828));
 AOI221xp5_ASAP7_75t_L g214590 (.A1(n_3497),
    .A2(n_1431),
    .B1(n_2421),
    .B2(sa13[7]),
    .C(n_5150),
    .Y(n_5827));
 OAI221xp5_ASAP7_75t_R g214591 (.A1(n_3839),
    .A2(n_2463),
    .B1(n_3066),
    .B2(sa12[7]),
    .C(n_2771),
    .Y(n_5826));
 AOI222xp33_ASAP7_75t_R g214592 (.A1(n_4311),
    .A2(n_2055),
    .B1(n_3058),
    .B2(n_1461),
    .C1(n_1653),
    .C2(n_2241),
    .Y(n_5825));
 AOI221xp5_ASAP7_75t_R g214593 (.A1(n_3055),
    .A2(sa31[6]),
    .B1(n_4319),
    .B2(n_1547),
    .C(n_2770),
    .Y(n_5824));
 AOI21xp33_ASAP7_75t_R g214594 (.A1(n_1561),
    .A2(n_4280),
    .B(n_4713),
    .Y(n_5823));
 AOI222xp33_ASAP7_75t_L g214595 (.A1(n_2735),
    .A2(n_1461),
    .B1(n_1652),
    .B2(n_2192),
    .C1(n_2055),
    .C2(n_2964),
    .Y(n_5822));
 AOI22xp5_ASAP7_75t_SL g214596 (.A1(n_2056),
    .A2(n_4364),
    .B1(n_1407),
    .B2(n_4363),
    .Y(n_5821));
 AOI221xp5_ASAP7_75t_L g214597 (.A1(n_2910),
    .A2(sa01[3]),
    .B1(n_3675),
    .B2(n_1465),
    .C(n_1638),
    .Y(n_5820));
 AOI322xp5_ASAP7_75t_SL g214598 (.A1(n_2788),
    .A2(n_2402),
    .A3(n_2279),
    .B1(n_1410),
    .B2(n_4483),
    .C1(n_1581),
    .C2(n_2014),
    .Y(n_5819));
 AOI221xp5_ASAP7_75t_SL g214599 (.A1(n_4057),
    .A2(n_4287),
    .B1(n_3057),
    .B2(sa11[6]),
    .C(n_2766),
    .Y(n_5818));
 AOI221xp5_ASAP7_75t_L g214600 (.A1(n_1570),
    .A2(n_8200),
    .B1(n_2507),
    .B2(n_1461),
    .C(n_5349),
    .Y(n_5817));
 AOI22xp33_ASAP7_75t_L g214601 (.A1(n_2047),
    .A2(n_3866),
    .B1(n_2066),
    .B2(n_3867),
    .Y(n_5816));
 AO22x1_ASAP7_75t_SL g214602 (.A1(n_3443),
    .A2(n_1784),
    .B1(n_3478),
    .B2(n_4399),
    .Y(n_5815));
 AOI22xp33_ASAP7_75t_R g214603 (.A1(n_1560),
    .A2(n_3888),
    .B1(n_1567),
    .B2(n_3889),
    .Y(n_5814));
 OAI221xp5_ASAP7_75t_L g214604 (.A1(n_3012),
    .A2(n_3313),
    .B1(n_2488),
    .B2(n_1972),
    .C(n_4670),
    .Y(n_5813));
 OAI22xp33_ASAP7_75t_L g214605 (.A1(n_3909),
    .A2(n_1542),
    .B1(n_3908),
    .B2(n_1446),
    .Y(n_5812));
 OAI222xp33_ASAP7_75t_L g214606 (.A1(n_3587),
    .A2(n_1363),
    .B1(n_2973),
    .B2(n_2395),
    .C1(n_2041),
    .C2(n_2307),
    .Y(n_5811));
 AOI221xp5_ASAP7_75t_SL g214607 (.A1(n_1559),
    .A2(n_2302),
    .B1(n_2970),
    .B2(n_2050),
    .C(n_4234),
    .Y(n_5810));
 AOI221xp5_ASAP7_75t_L g214608 (.A1(n_2447),
    .A2(n_1859),
    .B1(n_2831),
    .B2(n_3031),
    .C(n_4527),
    .Y(n_5809));
 OAI221xp5_ASAP7_75t_SL g214609 (.A1(n_2855),
    .A2(n_3006),
    .B1(n_2494),
    .B2(n_1343),
    .C(n_4547),
    .Y(n_5808));
 OAI222xp33_ASAP7_75t_R g214610 (.A1(n_2073),
    .A2(n_3154),
    .B1(n_1628),
    .B2(n_3064),
    .C1(n_1543),
    .C2(n_2312),
    .Y(n_5807));
 AOI221xp5_ASAP7_75t_L g214611 (.A1(n_2588),
    .A2(n_1439),
    .B1(n_2942),
    .B2(n_3087),
    .C(n_3752),
    .Y(n_5806));
 OAI221xp5_ASAP7_75t_L g214612 (.A1(n_4014),
    .A2(n_2495),
    .B1(n_2968),
    .B2(n_3498),
    .C(n_1980),
    .Y(n_5805));
 AOI322xp5_ASAP7_75t_SL g214613 (.A1(n_2777),
    .A2(n_1625),
    .A3(n_1620),
    .B1(sa30[6]),
    .B2(n_1774),
    .C1(n_1391),
    .C2(n_1484),
    .Y(n_5804));
 OAI222xp33_ASAP7_75t_L g214614 (.A1(n_3055),
    .A2(n_1642),
    .B1(n_2955),
    .B2(n_1635),
    .C1(n_2083),
    .C2(n_2242),
    .Y(n_5803));
 OAI221xp5_ASAP7_75t_R g214615 (.A1(n_4004),
    .A2(n_2489),
    .B1(n_3081),
    .B2(n_2919),
    .C(sa00[0]),
    .Y(n_5802));
 OAI211xp5_ASAP7_75t_R g214616 (.A1(n_1590),
    .A2(n_3872),
    .B(n_4549),
    .C(n_4152),
    .Y(n_5801));
 OAI221xp5_ASAP7_75t_L g214617 (.A1(n_4521),
    .A2(n_2395),
    .B1(n_2346),
    .B2(n_1935),
    .C(n_4276),
    .Y(n_5800));
 OAI221xp5_ASAP7_75t_SL g214618 (.A1(n_1417),
    .A2(n_2675),
    .B1(n_1654),
    .B2(n_2906),
    .C(n_4247),
    .Y(n_5799));
 AOI221xp5_ASAP7_75t_SL g214619 (.A1(n_3527),
    .A2(n_1561),
    .B1(n_4519),
    .B2(n_1566),
    .C(n_3233),
    .Y(n_5798));
 OAI211xp5_ASAP7_75t_L g214620 (.A1(n_2088),
    .A2(n_1764),
    .B(n_4166),
    .C(n_4542),
    .Y(n_5797));
 OAI222xp33_ASAP7_75t_R g214621 (.A1(n_1354),
    .A2(n_3491),
    .B1(n_4511),
    .B2(n_2396),
    .C1(n_2337),
    .C2(n_1394),
    .Y(n_5796));
 AOI222xp33_ASAP7_75t_R g214622 (.A1(n_1438),
    .A2(n_1702),
    .B1(n_3373),
    .B2(n_2065),
    .C1(n_1557),
    .C2(n_2896),
    .Y(n_5795));
 OAI22xp33_ASAP7_75t_L g214623 (.A1(n_2083),
    .A2(n_4360),
    .B1(n_1642),
    .B2(n_3724),
    .Y(n_5794));
 AOI221xp5_ASAP7_75t_R g214624 (.A1(n_3489),
    .A2(n_1439),
    .B1(n_2339),
    .B2(n_1496),
    .C(n_5145),
    .Y(n_5793));
 OAI221xp5_ASAP7_75t_R g214625 (.A1(n_1548),
    .A2(n_2640),
    .B1(n_1644),
    .B2(n_2889),
    .C(n_4243),
    .Y(n_5792));
 AOI222xp33_ASAP7_75t_L g214626 (.A1(n_1352),
    .A2(n_2650),
    .B1(n_2420),
    .B2(n_3330),
    .C1(n_2392),
    .C2(n_2914),
    .Y(n_5791));
 OAI22xp5_ASAP7_75t_L g214627 (.A1(n_1344),
    .A2(n_3880),
    .B1(n_1662),
    .B2(n_3715),
    .Y(n_5790));
 OAI221xp5_ASAP7_75t_R g214628 (.A1(n_4539),
    .A2(n_1975),
    .B1(sa21[3]),
    .B2(n_2253),
    .C(n_2763),
    .Y(n_5789));
 AOI222xp33_ASAP7_75t_R g214629 (.A1(n_2401),
    .A2(n_3357),
    .B1(n_2416),
    .B2(n_2899),
    .C1(n_1419),
    .C2(n_1694),
    .Y(n_5788));
 AOI221xp5_ASAP7_75t_L g214630 (.A1(n_3031),
    .A2(n_2851),
    .B1(n_3598),
    .B2(n_1463),
    .C(n_3677),
    .Y(n_5787));
 AOI211xp5_ASAP7_75t_SL g214631 (.A1(n_1770),
    .A2(n_1345),
    .B(n_4261),
    .C(n_1877),
    .Y(n_5786));
 OAI22xp5_ASAP7_75t_L g214632 (.A1(n_1381),
    .A2(n_3897),
    .B1(n_1640),
    .B2(n_3714),
    .Y(n_5785));
 OAI21xp33_ASAP7_75t_SL g214633 (.A1(n_2080),
    .A2(n_3877),
    .B(n_5365),
    .Y(n_5784));
 AOI222xp33_ASAP7_75t_L g214634 (.A1(n_2400),
    .A2(n_3419),
    .B1(n_1444),
    .B2(n_2617),
    .C1(n_1405),
    .C2(n_3320),
    .Y(n_5783));
 OAI211xp5_ASAP7_75t_L g214635 (.A1(n_2070),
    .A2(n_3876),
    .B(n_4642),
    .C(n_3735),
    .Y(n_5782));
 OAI22xp33_ASAP7_75t_R g214636 (.A1(n_3461),
    .A2(n_2974),
    .B1(n_4396),
    .B2(n_1337),
    .Y(n_5781));
 OAI221xp5_ASAP7_75t_R g214637 (.A1(n_1658),
    .A2(n_1736),
    .B1(n_2901),
    .B2(n_1660),
    .C(n_2738),
    .Y(n_5780));
 AOI222xp33_ASAP7_75t_SL g214638 (.A1(n_2058),
    .A2(n_3475),
    .B1(n_2342),
    .B2(n_1464),
    .C1(n_4543),
    .C2(n_2390),
    .Y(n_5779));
 OAI211xp5_ASAP7_75t_L g214639 (.A1(n_2083),
    .A2(n_3896),
    .B(n_4654),
    .C(n_4151),
    .Y(n_5778));
 OAI211xp5_ASAP7_75t_L g214640 (.A1(n_1344),
    .A2(n_4432),
    .B(n_4705),
    .C(n_4165),
    .Y(n_5777));
 OAI22xp33_ASAP7_75t_L g214641 (.A1(n_3523),
    .A2(n_4497),
    .B1(sa03[1]),
    .B2(n_4439),
    .Y(n_5776));
 OAI22xp33_ASAP7_75t_L g214642 (.A1(n_3611),
    .A2(n_4407),
    .B1(n_3381),
    .B2(n_3547),
    .Y(n_5775));
 AO32x1_ASAP7_75t_SL g214643 (.A1(n_4141),
    .A2(n_2094),
    .A3(n_1455),
    .B1(n_3077),
    .B2(sa12[1]),
    .Y(n_5774));
 AOI21xp5_ASAP7_75t_L g214644 (.A1(n_3892),
    .A2(n_2090),
    .B(n_5364),
    .Y(n_5773));
 OAI211xp5_ASAP7_75t_L g214645 (.A1(n_1850),
    .A2(n_1758),
    .B(n_4222),
    .C(n_3551),
    .Y(n_5772));
 OAI221xp5_ASAP7_75t_L g214646 (.A1(n_2932),
    .A2(n_3366),
    .B1(n_3536),
    .B2(n_1460),
    .C(n_3690),
    .Y(n_5771));
 OAI211xp5_ASAP7_75t_R g214647 (.A1(n_2063),
    .A2(n_4683),
    .B(n_4685),
    .C(n_4118),
    .Y(n_5770));
 OAI221xp5_ASAP7_75t_L g214648 (.A1(n_3895),
    .A2(n_1634),
    .B1(n_2531),
    .B2(n_1933),
    .C(n_3157),
    .Y(n_5769));
 OAI221xp5_ASAP7_75t_L g214649 (.A1(n_3032),
    .A2(n_3417),
    .B1(n_3565),
    .B2(n_1933),
    .C(n_3572),
    .Y(n_5768));
 AOI221xp5_ASAP7_75t_SL g214650 (.A1(n_3007),
    .A2(n_3287),
    .B1(n_3542),
    .B2(n_1498),
    .C(n_3649),
    .Y(n_5767));
 AOI211xp5_ASAP7_75t_SL g214651 (.A1(n_3894),
    .A2(n_1424),
    .B(n_4525),
    .C(n_4140),
    .Y(n_5766));
 AOI221xp5_ASAP7_75t_R g214652 (.A1(n_3017),
    .A2(n_3281),
    .B1(n_3553),
    .B2(n_1395),
    .C(n_3626),
    .Y(n_5765));
 OAI211xp5_ASAP7_75t_L g214653 (.A1(n_2073),
    .A2(n_3906),
    .B(n_4699),
    .C(n_4154),
    .Y(n_5764));
 OAI221xp5_ASAP7_75t_R g214654 (.A1(n_3293),
    .A2(n_3008),
    .B1(n_3567),
    .B2(n_1404),
    .C(n_3621),
    .Y(n_5763));
 OAI211xp5_ASAP7_75t_L g214655 (.A1(n_1337),
    .A2(n_3898),
    .B(n_4137),
    .C(n_4689),
    .Y(n_5762));
 OAI221xp5_ASAP7_75t_SL g214656 (.A1(n_3999),
    .A2(n_2066),
    .B1(n_1558),
    .B2(n_1689),
    .C(n_3683),
    .Y(n_5761));
 AOI211xp5_ASAP7_75t_L g214657 (.A1(n_4397),
    .A2(n_2089),
    .B(n_4530),
    .C(n_4106),
    .Y(n_5760));
 OAI211xp5_ASAP7_75t_L g214658 (.A1(n_1656),
    .A2(n_3978),
    .B(n_3629),
    .C(n_3131),
    .Y(n_5759));
 OAI211xp5_ASAP7_75t_L g214659 (.A1(n_1634),
    .A2(n_4462),
    .B(n_3619),
    .C(n_3133),
    .Y(n_5758));
 OAI211xp5_ASAP7_75t_L g214660 (.A1(n_1624),
    .A2(n_3976),
    .B(n_3620),
    .C(n_3075),
    .Y(n_5757));
 OAI221xp5_ASAP7_75t_L g214661 (.A1(n_3333),
    .A2(n_3146),
    .B1(n_3563),
    .B2(n_1459),
    .C(n_3681),
    .Y(n_5756));
 AOI211xp5_ASAP7_75t_L g214662 (.A1(n_3969),
    .A2(n_2404),
    .B(n_3123),
    .C(n_3627),
    .Y(n_5755));
 OAI221xp5_ASAP7_75t_R g214663 (.A1(n_3477),
    .A2(n_2539),
    .B1(n_3168),
    .B2(n_2415),
    .C(n_4531),
    .Y(n_5754));
 AOI32xp33_ASAP7_75t_SL g214664 (.A1(n_1737),
    .A2(n_8703),
    .A3(n_3155),
    .B1(n_1783),
    .B2(n_1987),
    .Y(n_5753));
 AOI322xp5_ASAP7_75t_L g214665 (.A1(n_3247),
    .A2(n_2435),
    .A3(n_1619),
    .B1(sa02[7]),
    .B2(n_2075),
    .C1(n_4532),
    .C2(n_1458),
    .Y(n_5752));
 OAI22xp33_ASAP7_75t_R g214666 (.A1(n_3465),
    .A2(n_4481),
    .B1(n_1478),
    .B2(n_4424),
    .Y(n_5751));
 OAI221xp5_ASAP7_75t_L g214667 (.A1(n_4599),
    .A2(n_1844),
    .B1(n_2396),
    .B2(n_2548),
    .C(n_4215),
    .Y(n_5750));
 OAI211xp5_ASAP7_75t_R g214668 (.A1(n_1658),
    .A2(n_3865),
    .B(n_4705),
    .C(n_3410),
    .Y(n_5749));
 OAI22xp33_ASAP7_75t_SL g214669 (.A1(n_3606),
    .A2(n_4473),
    .B1(n_1524),
    .B2(n_4475),
    .Y(n_5748));
 OAI221xp5_ASAP7_75t_L g214670 (.A1(n_4207),
    .A2(n_1624),
    .B1(n_1434),
    .B2(n_2149),
    .C(n_1870),
    .Y(n_5747));
 AOI221xp5_ASAP7_75t_L g214671 (.A1(n_4025),
    .A2(n_1664),
    .B1(n_1550),
    .B2(n_2210),
    .C(n_4610),
    .Y(n_5746));
 OAI21xp33_ASAP7_75t_SL g214672 (.A1(n_2463),
    .A2(n_4493),
    .B(n_5353),
    .Y(n_5745));
 AOI221xp5_ASAP7_75t_SL g214673 (.A1(n_4119),
    .A2(n_2847),
    .B1(n_2976),
    .B2(n_1595),
    .C(n_4643),
    .Y(n_5744));
 OAI22xp5_ASAP7_75t_R g214674 (.A1(n_2935),
    .A2(n_2953),
    .B1(n_1678),
    .B2(n_4020),
    .Y(n_5743));
 OAI211xp5_ASAP7_75t_L g214675 (.A1(n_2860),
    .A2(n_4099),
    .B(n_3736),
    .C(sa30[2]),
    .Y(n_5742));
 OAI22xp5_ASAP7_75t_R g214676 (.A1(n_4466),
    .A2(n_4448),
    .B1(n_1676),
    .B2(n_4495),
    .Y(n_5741));
 AOI221xp5_ASAP7_75t_L g214677 (.A1(n_2933),
    .A2(n_2192),
    .B1(n_4109),
    .B2(n_2837),
    .C(n_4645),
    .Y(n_5740));
 OAI22xp5_ASAP7_75t_R g214678 (.A1(n_2952),
    .A2(n_4439),
    .B1(n_2588),
    .B2(n_4437),
    .Y(n_5739));
 AOI221xp5_ASAP7_75t_L g214679 (.A1(n_4035),
    .A2(n_1446),
    .B1(n_1545),
    .B2(n_2134),
    .C(sa21[0]),
    .Y(n_5738));
 OAI321xp33_ASAP7_75t_SL g214680 (.A1(n_2780),
    .A2(n_1408),
    .A3(n_1614),
    .B1(n_1460),
    .B2(n_4449),
    .C(n_3652),
    .Y(n_5737));
 AOI221xp5_ASAP7_75t_SL g214681 (.A1(n_2951),
    .A2(n_2065),
    .B1(n_3142),
    .B2(n_2444),
    .C(n_2125),
    .Y(n_5736));
 OAI321xp33_ASAP7_75t_R g214682 (.A1(n_3244),
    .A2(n_1651),
    .A3(n_2321),
    .B1(n_1456),
    .B2(n_4684),
    .C(n_3643),
    .Y(n_5735));
 OAI321xp33_ASAP7_75t_L g214683 (.A1(n_2804),
    .A2(n_1658),
    .A3(n_2288),
    .B1(n_1850),
    .B2(n_4433),
    .C(n_3653),
    .Y(n_5734));
 AOI321xp33_ASAP7_75t_SL g214684 (.A1(n_2807),
    .A2(n_1633),
    .A3(n_2291),
    .B1(n_4509),
    .B2(sa31[6]),
    .C(n_3658),
    .Y(n_5733));
 OAI221xp5_ASAP7_75t_L g214685 (.A1(n_4355),
    .A2(n_1418),
    .B1(n_8691),
    .B2(n_3707),
    .C(n_1965),
    .Y(n_5732));
 AOI211xp5_ASAP7_75t_L g214686 (.A1(n_3886),
    .A2(n_1423),
    .B(n_4220),
    .C(n_4192),
    .Y(n_5731));
 AOI221xp5_ASAP7_75t_SL g214687 (.A1(n_3665),
    .A2(n_1398),
    .B1(n_3881),
    .B2(n_1424),
    .C(sa22[0]),
    .Y(n_5730));
 OAI211xp5_ASAP7_75t_R g214688 (.A1(n_2445),
    .A2(n_4208),
    .B(n_1439),
    .C(n_1533),
    .Y(n_5729));
 AOI221xp5_ASAP7_75t_R g214689 (.A1(n_3672),
    .A2(n_1638),
    .B1(n_3862),
    .B2(n_2087),
    .C(sa01[0]),
    .Y(n_5728));
 AOI322xp5_ASAP7_75t_R g214690 (.A1(n_2910),
    .A2(n_1734),
    .A3(n_1589),
    .B1(sa01[3]),
    .B2(n_3598),
    .C1(n_1638),
    .C2(n_1384),
    .Y(n_5727));
 OAI321xp33_ASAP7_75t_R g214691 (.A1(n_1580),
    .A2(n_2818),
    .A3(n_3345),
    .B1(n_2278),
    .B2(n_2415),
    .C(n_3022),
    .Y(n_5726));
 OAI221xp5_ASAP7_75t_L g214692 (.A1(n_3888),
    .A2(n_2091),
    .B1(n_1565),
    .B2(n_3727),
    .C(n_8203),
    .Y(n_5725));
 AO22x1_ASAP7_75t_L g214693 (.A1(n_1641),
    .A2(n_4640),
    .B1(n_2042),
    .B2(n_4445),
    .Y(n_5724));
 OAI221xp5_ASAP7_75t_L g214694 (.A1(n_4576),
    .A2(n_1392),
    .B1(n_1644),
    .B2(n_2292),
    .C(n_2980),
    .Y(n_5723));
 AOI321xp33_ASAP7_75t_L g214695 (.A1(n_1745),
    .A2(n_3284),
    .A3(n_2092),
    .B1(n_2394),
    .B2(n_1618),
    .C(n_2975),
    .Y(n_5722));
 AOI22xp33_ASAP7_75t_R g214696 (.A1(n_1397),
    .A2(n_4006),
    .B1(n_2532),
    .B2(n_2040),
    .Y(n_5721));
 AOI221xp5_ASAP7_75t_L g214697 (.A1(n_3043),
    .A2(n_1405),
    .B1(n_3037),
    .B2(n_2464),
    .C(n_2179),
    .Y(n_5720));
 AOI322xp5_ASAP7_75t_R g214698 (.A1(n_3415),
    .A2(n_2064),
    .A3(n_1735),
    .B1(n_1512),
    .B2(n_3641),
    .C1(n_8703),
    .C2(n_1953),
    .Y(n_5719));
 AOI321xp33_ASAP7_75t_L g214699 (.A1(n_3257),
    .A2(n_3341),
    .A3(n_1424),
    .B1(n_2397),
    .B2(n_2295),
    .C(n_2985),
    .Y(n_5718));
 AOI221xp5_ASAP7_75t_R g214700 (.A1(n_2956),
    .A2(n_2387),
    .B1(n_3132),
    .B2(n_1682),
    .C(n_2625),
    .Y(n_5717));
 OAI322xp33_ASAP7_75t_SL g214701 (.A1(n_3347),
    .A2(n_2083),
    .A3(n_2904),
    .B1(n_8181),
    .B2(n_3565),
    .C1(n_1644),
    .C2(sa31[4]),
    .Y(n_5716));
 AOI32xp33_ASAP7_75t_L g214702 (.A1(n_4661),
    .A2(n_2092),
    .A3(n_2110),
    .B1(n_4521),
    .B2(n_2394),
    .Y(n_5715));
 AOI22xp33_ASAP7_75t_R g214703 (.A1(n_3447),
    .A2(n_2985),
    .B1(n_1683),
    .B2(n_4008),
    .Y(n_5714));
 AOI21xp5_ASAP7_75t_SL g214704 (.A1(n_4539),
    .A2(n_1401),
    .B(n_3780),
    .Y(n_5713));
 AOI32xp33_ASAP7_75t_R g214705 (.A1(n_4608),
    .A2(n_1366),
    .A3(n_1595),
    .B1(n_4508),
    .B2(n_2046),
    .Y(n_5712));
 AOI211xp5_ASAP7_75t_SL g214706 (.A1(n_3007),
    .A2(n_2205),
    .B(n_4160),
    .C(n_1981),
    .Y(n_5711));
 OAI221xp5_ASAP7_75t_R g214707 (.A1(n_4483),
    .A2(n_1578),
    .B1(n_2415),
    .B2(n_3490),
    .C(n_4041),
    .Y(n_5710));
 OAI322xp33_ASAP7_75t_L g214708 (.A1(n_3424),
    .A2(n_2081),
    .A3(n_3369),
    .B1(n_3552),
    .B2(n_1985),
    .C1(n_2396),
    .C2(sa22[4]),
    .Y(n_5709));
 AOI32xp33_ASAP7_75t_R g214709 (.A1(n_2883),
    .A2(n_3367),
    .A3(n_2079),
    .B1(n_1445),
    .B2(n_1949),
    .Y(n_5708));
 OAI22xp5_ASAP7_75t_L g214710 (.A1(n_3988),
    .A2(n_1461),
    .B1(n_2508),
    .B2(n_2056),
    .Y(n_5707));
 AOI221xp5_ASAP7_75t_L g214711 (.A1(n_2054),
    .A2(n_2501),
    .B1(n_1398),
    .B2(n_3666),
    .C(n_8217),
    .Y(n_5706));
 AOI22xp33_ASAP7_75t_R g214712 (.A1(n_1456),
    .A2(n_4000),
    .B1(n_2510),
    .B2(n_2077),
    .Y(n_5705));
 OAI32xp33_ASAP7_75t_L g214713 (.A1(n_2885),
    .A2(n_3356),
    .A3(n_2073),
    .B1(n_1503),
    .B2(n_1628),
    .Y(n_5704));
 OAI311xp33_ASAP7_75t_R g214714 (.A1(n_3280),
    .A2(n_3423),
    .A3(n_2081),
    .B1(n_4032),
    .C1(n_4680),
    .Y(n_5703));
 AOI221xp5_ASAP7_75t_L g214715 (.A1(n_4120),
    .A2(n_2831),
    .B1(n_3031),
    .B2(n_2171),
    .C(n_1785),
    .Y(n_5702));
 OAI32xp33_ASAP7_75t_L g214716 (.A1(n_4453),
    .A2(n_3375),
    .A3(n_1571),
    .B1(n_4424),
    .B2(n_4506),
    .Y(n_5701));
 OAI221xp5_ASAP7_75t_L g214717 (.A1(n_2041),
    .A2(n_2594),
    .B1(n_3460),
    .B2(n_2430),
    .C(n_3826),
    .Y(n_5700));
 OAI221xp5_ASAP7_75t_R g214718 (.A1(n_1543),
    .A2(n_2523),
    .B1(n_1628),
    .B2(n_3717),
    .C(sa21[0]),
    .Y(n_5699));
 AO21x1_ASAP7_75t_L g214719 (.A1(n_2400),
    .A2(n_4621),
    .B(n_3783),
    .Y(n_5698));
 AOI221xp5_ASAP7_75t_L g214720 (.A1(n_3128),
    .A2(n_2494),
    .B1(n_3096),
    .B2(n_1569),
    .C(n_3585),
    .Y(n_5697));
 OAI311xp33_ASAP7_75t_R g214721 (.A1(n_3448),
    .A2(n_1590),
    .A3(n_2852),
    .B1(n_4180),
    .C1(n_4556),
    .Y(n_5696));
 AO32x1_ASAP7_75t_SL g214722 (.A1(n_4617),
    .A2(n_2095),
    .A3(n_1576),
    .B1(n_4460),
    .B2(n_2429),
    .Y(n_5695));
 AOI221xp5_ASAP7_75t_R g214723 (.A1(n_3221),
    .A2(n_2392),
    .B1(n_1431),
    .B2(n_2554),
    .C(n_8188),
    .Y(n_5694));
 AOI22xp33_ASAP7_75t_R g214724 (.A1(n_2223),
    .A2(n_3915),
    .B1(n_1447),
    .B2(n_3872),
    .Y(n_5693));
 OAI22xp33_ASAP7_75t_L g214725 (.A1(n_2430),
    .A2(n_4669),
    .B1(n_1551),
    .B2(n_4025),
    .Y(n_5692));
 OAI321xp33_ASAP7_75t_L g214726 (.A1(n_2797),
    .A2(n_2866),
    .A3(n_2088),
    .B1(n_2326),
    .B2(n_1553),
    .C(n_3086),
    .Y(n_5691));
 AO22x1_ASAP7_75t_SL g214727 (.A1(n_3025),
    .A2(n_4419),
    .B1(n_2561),
    .B2(n_4421),
    .Y(n_5690));
 AOI221xp5_ASAP7_75t_R g214728 (.A1(n_3130),
    .A2(n_2471),
    .B1(n_3025),
    .B2(n_1657),
    .C(n_3582),
    .Y(n_5689));
 AOI321xp33_ASAP7_75t_SL g214729 (.A1(n_3254),
    .A2(n_1412),
    .A3(n_3406),
    .B1(n_2050),
    .B2(n_2318),
    .C(n_2967),
    .Y(n_5688));
 OAI211xp5_ASAP7_75t_SL g214730 (.A1(n_1392),
    .A2(n_4509),
    .B(n_4535),
    .C(n_4202),
    .Y(n_5687));
 AOI221xp5_ASAP7_75t_R g214731 (.A1(n_3177),
    .A2(n_1352),
    .B1(n_2420),
    .B2(n_3506),
    .C(n_2565),
    .Y(n_5686));
 OAI322xp33_ASAP7_75t_R g214732 (.A1(n_2015),
    .A2(n_1850),
    .A3(n_2187),
    .B1(n_1986),
    .B2(n_2881),
    .C1(n_2096),
    .C2(n_3860),
    .Y(n_5685));
 AOI311xp33_ASAP7_75t_SL g214733 (.A1(n_3287),
    .A2(n_3425),
    .A3(n_1412),
    .B(n_4681),
    .C(n_4185),
    .Y(n_5684));
 OAI32xp33_ASAP7_75t_L g214734 (.A1(n_4582),
    .A2(n_1580),
    .A3(n_2102),
    .B1(n_1357),
    .B2(n_4482),
    .Y(n_5683));
 AOI211xp5_ASAP7_75t_SL g214735 (.A1(n_1763),
    .A2(n_1439),
    .B(n_2125),
    .C(n_3186),
    .Y(n_5682));
 AO32x1_ASAP7_75t_SL g214736 (.A1(n_4410),
    .A2(n_3392),
    .A3(n_2062),
    .B1(n_4425),
    .B2(n_4545),
    .Y(n_5681));
 OAI221xp5_ASAP7_75t_L g214737 (.A1(n_3851),
    .A2(sa30[6]),
    .B1(n_2043),
    .B2(n_2512),
    .C(n_1924),
    .Y(n_5680));
 AOI311xp33_ASAP7_75t_L g214738 (.A1(n_3450),
    .A2(n_3329),
    .A3(n_2092),
    .B(n_4203),
    .C(n_4666),
    .Y(n_5679));
 OAI211xp5_ASAP7_75t_L g214739 (.A1(n_1629),
    .A2(n_4566),
    .B(n_3196),
    .C(n_2649),
    .Y(n_5678));
 AOI211xp5_ASAP7_75t_SL g214740 (.A1(n_4605),
    .A2(n_8703),
    .B(n_3208),
    .C(n_1591),
    .Y(n_5677));
 AOI211xp5_ASAP7_75t_L g214741 (.A1(n_4591),
    .A2(n_2392),
    .B(n_3205),
    .C(n_2221),
    .Y(n_5676));
 AOI22xp33_ASAP7_75t_R g214742 (.A1(n_2174),
    .A2(n_3926),
    .B1(n_1431),
    .B2(n_3877),
    .Y(n_5675));
 OAI21xp33_ASAP7_75t_L g214743 (.A1(n_4436),
    .A2(n_4475),
    .B(n_4882),
    .Y(n_5674));
 AOI32xp33_ASAP7_75t_R g214744 (.A1(n_4505),
    .A2(n_3343),
    .A3(n_2089),
    .B1(n_4438),
    .B2(n_4588),
    .Y(n_5673));
 AOI22xp33_ASAP7_75t_L g214745 (.A1(n_1645),
    .A2(n_4476),
    .B1(n_1372),
    .B2(n_3033),
    .Y(n_5672));
 AOI321xp33_ASAP7_75t_SL g214746 (.A1(n_3262),
    .A2(n_2064),
    .A3(n_1746),
    .B1(n_8703),
    .B2(n_2320),
    .C(n_3065),
    .Y(n_5671));
 OAI22xp5_ASAP7_75t_SL g214747 (.A1(n_1747),
    .A2(n_4124),
    .B1(n_2063),
    .B2(n_2979),
    .Y(n_5670));
 AOI211xp5_ASAP7_75t_L g214748 (.A1(n_4553),
    .A2(n_2398),
    .B(n_3190),
    .C(n_2625),
    .Y(n_5669));
 OAI22xp5_ASAP7_75t_R g214749 (.A1(n_3095),
    .A2(n_4475),
    .B1(n_2530),
    .B2(n_4473),
    .Y(n_5668));
 OAI221xp5_ASAP7_75t_L g214750 (.A1(n_3975),
    .A2(n_1666),
    .B1(n_1590),
    .B2(sa01[7]),
    .C(n_3135),
    .Y(n_5667));
 OA211x2_ASAP7_75t_SL g214751 (.A1(n_1639),
    .A2(n_4563),
    .B(n_3193),
    .C(n_2273),
    .Y(n_5666));
 OAI211xp5_ASAP7_75t_R g214752 (.A1(n_2078),
    .A2(n_1774),
    .B(n_4690),
    .C(n_4172),
    .Y(n_5665));
 AOI22xp5_ASAP7_75t_R g214753 (.A1(n_3952),
    .A2(n_2172),
    .B1(n_3896),
    .B2(n_2040),
    .Y(n_5664));
 AOI22xp33_ASAP7_75t_R g214754 (.A1(n_1398),
    .A2(n_4373),
    .B1(n_3659),
    .B2(n_1424),
    .Y(n_5663));
 AOI22xp33_ASAP7_75t_L g214755 (.A1(n_1652),
    .A2(n_4507),
    .B1(n_1572),
    .B2(n_3723),
    .Y(n_5662));
 AOI321xp33_ASAP7_75t_SL g214756 (.A1(n_3246),
    .A2(n_1717),
    .A3(n_1570),
    .B1(n_1653),
    .B2(n_1613),
    .C(n_3080),
    .Y(n_5661));
 OAI22xp33_ASAP7_75t_R g214757 (.A1(n_1637),
    .A2(n_4492),
    .B1(n_1588),
    .B2(n_3699),
    .Y(n_5660));
 AOI22xp33_ASAP7_75t_L g214758 (.A1(n_1566),
    .A2(n_4435),
    .B1(n_2090),
    .B2(n_3705),
    .Y(n_5659));
 AOI321xp33_ASAP7_75t_SL g214759 (.A1(n_2807),
    .A2(n_2857),
    .A3(n_1645),
    .B1(n_3515),
    .B2(n_2084),
    .C(n_2626),
    .Y(n_5658));
 AOI22xp33_ASAP7_75t_SL g214760 (.A1(n_2394),
    .A2(n_4413),
    .B1(n_1374),
    .B2(n_3169),
    .Y(n_5657));
 OAI22xp33_ASAP7_75t_L g214761 (.A1(n_1639),
    .A2(n_4446),
    .B1(n_3140),
    .B2(n_1381),
    .Y(n_5656));
 OAI22xp33_ASAP7_75t_R g214762 (.A1(n_1660),
    .A2(n_4451),
    .B1(n_3126),
    .B2(n_1344),
    .Y(n_5655));
 OAI22xp5_ASAP7_75t_SL g214763 (.A1(n_2411),
    .A2(n_4571),
    .B1(n_2056),
    .B2(n_3964),
    .Y(n_5654));
 OAI211xp5_ASAP7_75t_L g214764 (.A1(n_2419),
    .A2(n_4571),
    .B(n_3194),
    .C(n_2258),
    .Y(n_5653));
 AOI21xp5_ASAP7_75t_R g214765 (.A1(n_4581),
    .A2(n_2429),
    .B(n_3768),
    .Y(n_5652));
 AOI311xp33_ASAP7_75t_R g214766 (.A1(n_3292),
    .A2(n_1752),
    .A3(n_1586),
    .B(n_4116),
    .C(n_4688),
    .Y(n_5651));
 AOI221xp5_ASAP7_75t_L g214767 (.A1(n_4051),
    .A2(n_2069),
    .B1(n_1659),
    .B2(n_1616),
    .C(n_2947),
    .Y(n_5650));
 AOI211xp5_ASAP7_75t_R g214768 (.A1(n_4631),
    .A2(n_2051),
    .B(n_3209),
    .C(n_2266),
    .Y(n_5649));
 AO21x1_ASAP7_75t_L g214769 (.A1(n_1587),
    .A2(n_4044),
    .B(n_3782),
    .Y(n_5648));
 OAI221xp5_ASAP7_75t_R g214770 (.A1(n_4552),
    .A2(n_2078),
    .B1(n_1639),
    .B2(n_2333),
    .C(n_3085),
    .Y(n_5647));
 AOI311xp33_ASAP7_75t_R g214771 (.A1(n_3334),
    .A2(n_2886),
    .A3(n_1423),
    .B(n_4163),
    .C(n_4673),
    .Y(n_5646));
 OAI221xp5_ASAP7_75t_L g214772 (.A1(n_1583),
    .A2(n_1953),
    .B1(n_2895),
    .B2(n_1455),
    .C(n_1608),
    .Y(n_5645));
 AOI221xp5_ASAP7_75t_R g214773 (.A1(n_2913),
    .A2(n_1404),
    .B1(n_1431),
    .B2(n_1504),
    .C(n_2201),
    .Y(n_5644));
 AOI221xp5_ASAP7_75t_R g214774 (.A1(n_3418),
    .A2(n_1459),
    .B1(n_2067),
    .B2(n_1954),
    .C(n_2225),
    .Y(n_5643));
 OAI321xp33_ASAP7_75t_R g214775 (.A1(n_2074),
    .A2(n_3282),
    .A3(n_3525),
    .B1(n_2322),
    .B2(n_2399),
    .C(n_3059),
    .Y(n_5642));
 OAI22xp33_ASAP7_75t_R g214776 (.A1(n_2393),
    .A2(n_4466),
    .B1(n_3151),
    .B2(n_2080),
    .Y(n_5641));
 AOI221xp5_ASAP7_75t_R g214777 (.A1(n_2901),
    .A2(n_1850),
    .B1(n_2044),
    .B2(n_1387),
    .C(n_2190),
    .Y(n_5640));
 AOI221xp5_ASAP7_75t_L g214778 (.A1(n_4054),
    .A2(n_2512),
    .B1(n_3036),
    .B2(sa30[6]),
    .C(n_3613),
    .Y(n_5639));
 OAI22xp33_ASAP7_75t_R g214779 (.A1(n_2830),
    .A2(n_3946),
    .B1(n_2584),
    .B2(n_3545),
    .Y(n_5638));
 AOI22xp33_ASAP7_75t_R g214780 (.A1(n_1440),
    .A2(n_4373),
    .B1(n_1424),
    .B2(n_4374),
    .Y(n_5637));
 OAI221xp5_ASAP7_75t_L g214781 (.A1(n_3069),
    .A2(n_1473),
    .B1(n_3178),
    .B2(n_2393),
    .C(n_4702),
    .Y(n_5636));
 AOI22xp33_ASAP7_75t_R g214782 (.A1(n_1587),
    .A2(n_4315),
    .B1(n_1638),
    .B2(n_4290),
    .Y(n_5635));
 AOI22xp33_ASAP7_75t_L g214783 (.A1(n_1643),
    .A2(n_4554),
    .B1(n_1682),
    .B2(n_2387),
    .Y(n_5634));
 OAI22xp5_ASAP7_75t_R g214784 (.A1(n_8702),
    .A2(n_4696),
    .B1(n_2063),
    .B2(n_4465),
    .Y(n_5633));
 AOI322xp5_ASAP7_75t_R g214785 (.A1(n_2100),
    .A2(n_1935),
    .A3(n_1921),
    .B1(n_1972),
    .B2(n_3429),
    .C1(n_3273),
    .C2(n_3184),
    .Y(n_5632));
 OAI22xp33_ASAP7_75t_L g214786 (.A1(n_1546),
    .A2(n_4509),
    .B1(n_2559),
    .B2(n_1632),
    .Y(n_5631));
 AOI221xp5_ASAP7_75t_L g214787 (.A1(n_1424),
    .A2(n_1610),
    .B1(n_2982),
    .B2(n_2427),
    .C(n_3831),
    .Y(n_5630));
 OAI22xp33_ASAP7_75t_R g214788 (.A1(n_4422),
    .A2(n_4675),
    .B1(n_2489),
    .B2(n_4481),
    .Y(n_5629));
 OAI322xp33_ASAP7_75t_R g214789 (.A1(n_2437),
    .A2(n_2506),
    .A3(n_8180),
    .B1(n_1379),
    .B2(n_2099),
    .C1(n_4322),
    .C2(n_2041),
    .Y(n_5628));
 OAI22xp5_ASAP7_75t_L g214790 (.A1(n_1628),
    .A2(n_4384),
    .B1(n_1678),
    .B2(n_2424),
    .Y(n_5627));
 OAI22xp5_ASAP7_75t_R g214791 (.A1(n_2041),
    .A2(n_4414),
    .B1(n_2487),
    .B2(n_2430),
    .Y(n_5626));
 OAI22xp33_ASAP7_75t_L g214792 (.A1(n_1666),
    .A2(n_4490),
    .B1(n_2057),
    .B2(n_2813),
    .Y(n_5625));
 OAI221xp5_ASAP7_75t_R g214793 (.A1(n_2973),
    .A2(n_2430),
    .B1(n_1363),
    .B2(n_2212),
    .C(n_3829),
    .Y(n_5624));
 OAI221xp5_ASAP7_75t_R g214794 (.A1(n_3345),
    .A2(n_4098),
    .B1(n_1580),
    .B2(n_3029),
    .C(n_1869),
    .Y(n_5623));
 OAI322xp33_ASAP7_75t_R g214795 (.A1(n_4292),
    .A2(n_3263),
    .A3(n_1582),
    .B1(n_2063),
    .B2(sa12[4]),
    .C1(n_2509),
    .C2(n_1456),
    .Y(n_5622));
 OAI22xp5_ASAP7_75t_L g214796 (.A1(n_1578),
    .A2(n_4404),
    .B1(n_1679),
    .B2(n_1647),
    .Y(n_5621));
 OAI322xp33_ASAP7_75t_L g214797 (.A1(n_4288),
    .A2(n_3269),
    .A3(n_2045),
    .B1(n_1344),
    .B2(n_1387),
    .C1(n_2519),
    .C2(n_1850),
    .Y(n_5620));
 AOI221xp5_ASAP7_75t_R g214798 (.A1(n_2064),
    .A2(n_2019),
    .B1(n_3981),
    .B2(n_2413),
    .C(n_3134),
    .Y(n_5619));
 OA211x2_ASAP7_75t_L g214799 (.A1(n_2073),
    .A2(n_4491),
    .B(n_4537),
    .C(n_4033),
    .Y(n_5618));
 AOI221xp5_ASAP7_75t_R g214800 (.A1(n_3645),
    .A2(n_1627),
    .B1(n_3519),
    .B2(n_1542),
    .C(n_3662),
    .Y(n_5617));
 AOI322xp5_ASAP7_75t_R g214801 (.A1(n_4300),
    .A2(n_3276),
    .A3(n_1352),
    .B1(n_1505),
    .B2(n_1586),
    .C1(n_2504),
    .C2(n_1934),
    .Y(n_5616));
 OAI22xp33_ASAP7_75t_R g214802 (.A1(n_2078),
    .A2(n_4443),
    .B1(n_1671),
    .B2(n_1623),
    .Y(n_5615));
 AOI22xp33_ASAP7_75t_R g214803 (.A1(n_4286),
    .A2(n_1625),
    .B1(n_1391),
    .B2(n_2551),
    .Y(n_5614));
 AOI22xp5_ASAP7_75t_L g214804 (.A1(n_4287),
    .A2(n_1655),
    .B1(n_2069),
    .B2(n_2592),
    .Y(n_5613));
 OAI221xp5_ASAP7_75t_R g214805 (.A1(n_1408),
    .A2(n_3966),
    .B1(n_1573),
    .B2(n_1483),
    .C(n_3078),
    .Y(n_5612));
 OAI32xp33_ASAP7_75t_L g214806 (.A1(n_4450),
    .A2(n_1738),
    .A3(n_1575),
    .B1(n_4635),
    .B2(n_4420),
    .Y(n_5611));
 OAI22xp33_ASAP7_75t_R g214807 (.A1(n_1408),
    .A2(n_4487),
    .B1(n_2490),
    .B2(n_1342),
    .Y(n_5610));
 AOI322xp5_ASAP7_75t_R g214808 (.A1(n_2865),
    .A2(n_2571),
    .A3(n_2062),
    .B1(n_1410),
    .B2(n_3079),
    .C1(n_1451),
    .C2(n_1905),
    .Y(n_5609));
 OAI322xp33_ASAP7_75t_L g214809 (.A1(n_2594),
    .A2(n_2487),
    .A3(n_8180),
    .B1(n_2972),
    .B2(n_1551),
    .C1(n_2395),
    .C2(n_2111),
    .Y(n_5608));
 OAI32xp33_ASAP7_75t_R g214810 (.A1(n_3245),
    .A2(n_1408),
    .A3(n_2838),
    .B1(n_1478),
    .B2(n_3078),
    .Y(n_5607));
 OAI221xp5_ASAP7_75t_SL g214811 (.A1(n_3948),
    .A2(n_2423),
    .B1(n_1584),
    .B2(sa13[7]),
    .C(n_3069),
    .Y(n_5606));
 OAI32xp33_ASAP7_75t_L g214812 (.A1(n_1543),
    .A2(n_2786),
    .A3(n_3356),
    .B1(n_4383),
    .B2(n_2073),
    .Y(n_5605));
 OAI32xp33_ASAP7_75t_L g214813 (.A1(n_2783),
    .A2(n_2052),
    .A3(n_2449),
    .B1(n_1568),
    .B2(n_4632),
    .Y(n_5604));
 OAI21xp5_ASAP7_75t_L g214814 (.A1(n_1442),
    .A2(n_4624),
    .B(n_3773),
    .Y(n_5603));
 AOI22xp33_ASAP7_75t_L g214815 (.A1(n_1432),
    .A2(n_3996),
    .B1(n_2588),
    .B2(n_1555),
    .Y(n_5602));
 AOI322xp5_ASAP7_75t_SL g214816 (.A1(n_2464),
    .A2(n_2557),
    .A3(n_1458),
    .B1(n_2067),
    .B2(n_3044),
    .C1(n_2400),
    .C2(n_1605),
    .Y(n_5601));
 OAI322xp33_ASAP7_75t_R g214817 (.A1(n_2560),
    .A2(n_1681),
    .A3(n_1933),
    .B1(n_1548),
    .B2(n_2956),
    .C1(n_1644),
    .C2(n_2104),
    .Y(n_5600));
 OAI22xp5_ASAP7_75t_L g214818 (.A1(n_1635),
    .A2(n_4513),
    .B1(n_1682),
    .B2(n_2083),
    .Y(n_5599));
 OAI21xp33_ASAP7_75t_L g214819 (.A1(n_2908),
    .A2(n_4129),
    .B(n_5027),
    .Y(n_5598));
 AOI322xp5_ASAP7_75t_L g214820 (.A1(n_2549),
    .A2(n_2458),
    .A3(n_1934),
    .B1(n_2178),
    .B2(n_1436),
    .C1(n_3046),
    .C2(n_1352),
    .Y(n_5597));
 AOI22xp33_ASAP7_75t_R g214821 (.A1(n_1667),
    .A2(n_4117),
    .B1(n_2584),
    .B2(n_2390),
    .Y(n_5596));
 AOI22xp33_ASAP7_75t_L g214822 (.A1(n_2427),
    .A2(n_4510),
    .B1(n_2492),
    .B2(n_2082),
    .Y(n_5595));
 AOI22xp33_ASAP7_75t_R g214823 (.A1(n_2413),
    .A2(n_4499),
    .B1(n_2463),
    .B2(n_2064),
    .Y(n_5594));
 OAI32xp33_ASAP7_75t_R g214824 (.A1(n_1727),
    .A2(n_1429),
    .A3(n_2451),
    .B1(n_2423),
    .B2(n_4590),
    .Y(n_5593));
 OAI22xp33_ASAP7_75t_R g214825 (.A1(n_2424),
    .A2(n_4566),
    .B1(n_2786),
    .B2(n_3045),
    .Y(n_5592));
 OAI22xp5_ASAP7_75t_L g214826 (.A1(n_2423),
    .A2(n_4496),
    .B1(n_1675),
    .B2(n_2080),
    .Y(n_5591));
 OAI22xp33_ASAP7_75t_R g214827 (.A1(n_1651),
    .A2(n_4657),
    .B1(n_2575),
    .B2(n_8691),
    .Y(n_5590));
 AOI22xp33_ASAP7_75t_R g214828 (.A1(n_3961),
    .A2(n_2392),
    .B1(n_1585),
    .B2(n_3574),
    .Y(n_5589));
 AOI22xp33_ASAP7_75t_R g214829 (.A1(n_2401),
    .A2(n_4482),
    .B1(n_1679),
    .B2(n_1577),
    .Y(n_5588));
 OAI22xp33_ASAP7_75t_L g214830 (.A1(n_2422),
    .A2(n_4196),
    .B1(n_2553),
    .B2(n_1429),
    .Y(n_5587));
 OAI22xp5_ASAP7_75t_SL g214831 (.A1(n_1634),
    .A2(n_4078),
    .B1(n_2568),
    .B2(n_1642),
    .Y(n_5586));
 AOI211xp5_ASAP7_75t_L g214832 (.A1(n_2781),
    .A2(n_1441),
    .B(n_4140),
    .C(n_8217),
    .Y(n_5585));
 AOI22xp33_ASAP7_75t_R g214833 (.A1(n_2089),
    .A2(n_3845),
    .B1(n_2046),
    .B2(n_4332),
    .Y(n_5584));
 AOI22xp33_ASAP7_75t_R g214834 (.A1(n_1349),
    .A2(n_4470),
    .B1(n_2530),
    .B2(n_1566),
    .Y(n_5583));
 AOI22xp33_ASAP7_75t_SL g214835 (.A1(n_3073),
    .A2(n_4101),
    .B1(n_3118),
    .B2(n_3077),
    .Y(n_5582));
 OA21x2_ASAP7_75t_L g214836 (.A1(n_3313),
    .A2(n_4168),
    .B(n_4865),
    .Y(n_5581));
 AOI22xp33_ASAP7_75t_L g214837 (.A1(n_1655),
    .A2(n_4145),
    .B1(n_2562),
    .B2(n_1659),
    .Y(n_5580));
 AOI22xp33_ASAP7_75t_L g214838 (.A1(n_2429),
    .A2(n_4551),
    .B1(n_2069),
    .B2(n_2814),
    .Y(n_5579));
 OAI211xp5_ASAP7_75t_R g214839 (.A1(n_1560),
    .A2(n_2783),
    .B(n_4149),
    .C(n_1980),
    .Y(n_5578));
 AOI22xp5_ASAP7_75t_R g214840 (.A1(n_2084),
    .A2(n_1778),
    .B1(n_2398),
    .B2(n_4320),
    .Y(n_5577));
 AOI221xp5_ASAP7_75t_L g214841 (.A1(n_3610),
    .A2(n_2503),
    .B1(n_4353),
    .B2(n_1585),
    .C(n_1966),
    .Y(n_5576));
 OAI22xp5_ASAP7_75t_L g214842 (.A1(n_1656),
    .A2(n_4460),
    .B1(n_2471),
    .B2(n_1575),
    .Y(n_5575));
 AO221x1_ASAP7_75t_L g214843 (.A1(n_4087),
    .A2(n_3260),
    .B1(n_3169),
    .B2(n_8180),
    .C(n_4203),
    .Y(n_5574));
 AOI221xp5_ASAP7_75t_R g214844 (.A1(n_2927),
    .A2(n_1569),
    .B1(n_3076),
    .B2(n_2090),
    .C(n_2609),
    .Y(n_5573));
 OAI211xp5_ASAP7_75t_L g214845 (.A1(n_1571),
    .A2(n_3990),
    .B(n_4178),
    .C(sa00[0]),
    .Y(n_5572));
 OAI22xp33_ASAP7_75t_R g214846 (.A1(n_2434),
    .A2(n_4637),
    .B1(n_2521),
    .B2(n_2399),
    .Y(n_5571));
 AOI22xp33_ASAP7_75t_R g214847 (.A1(n_1581),
    .A2(n_4297),
    .B1(n_1453),
    .B2(n_4293),
    .Y(n_5570));
 AOI22xp33_ASAP7_75t_R g214848 (.A1(n_1399),
    .A2(n_4598),
    .B1(n_1844),
    .B2(n_3438),
    .Y(n_5569));
 OAI221xp5_ASAP7_75t_R g214849 (.A1(n_4085),
    .A2(n_1729),
    .B1(n_3704),
    .B2(n_1498),
    .C(n_4184),
    .Y(n_5568));
 AOI22xp33_ASAP7_75t_L g214850 (.A1(n_1446),
    .A2(n_4136),
    .B1(n_2524),
    .B2(n_1350),
    .Y(n_5567));
 AOI22xp33_ASAP7_75t_L g214851 (.A1(n_1566),
    .A2(n_4638),
    .B1(n_1499),
    .B2(n_1749),
    .Y(n_5566));
 AOI221xp5_ASAP7_75t_L g214852 (.A1(n_4079),
    .A2(n_2807),
    .B1(n_3725),
    .B2(n_1933),
    .C(n_4201),
    .Y(n_5565));
 AOI22xp33_ASAP7_75t_R g214853 (.A1(n_4396),
    .A2(n_2394),
    .B1(n_3372),
    .B2(n_8180),
    .Y(n_5564));
 AOI221xp5_ASAP7_75t_L g214854 (.A1(n_3150),
    .A2(n_1403),
    .B1(n_4091),
    .B2(n_3258),
    .C(n_4116),
    .Y(n_5563));
 OAI221xp5_ASAP7_75t_R g214855 (.A1(n_4066),
    .A2(n_2787),
    .B1(n_3172),
    .B2(n_1346),
    .C(n_4041),
    .Y(n_5562));
 OA21x2_ASAP7_75t_L g214856 (.A1(n_2465),
    .A2(n_4484),
    .B(n_4934),
    .Y(n_5561));
 OAI211xp5_ASAP7_75t_SL g214857 (.A1(n_1442),
    .A2(n_3936),
    .B(n_4251),
    .C(n_4183),
    .Y(n_5560));
 AOI22xp33_ASAP7_75t_L g214858 (.A1(n_1445),
    .A2(n_4562),
    .B1(n_1353),
    .B2(n_1719),
    .Y(n_5559));
 AOI22xp33_ASAP7_75t_R g214859 (.A1(n_1627),
    .A2(n_4150),
    .B1(n_1501),
    .B2(n_2915),
    .Y(n_5558));
 AOI221xp5_ASAP7_75t_L g214860 (.A1(n_4080),
    .A2(n_2805),
    .B1(n_3125),
    .B2(n_1850),
    .C(n_4164),
    .Y(n_5557));
 OAI221xp5_ASAP7_75t_L g214861 (.A1(n_4074),
    .A2(n_1714),
    .B1(n_3699),
    .B2(n_1463),
    .C(n_4180),
    .Y(n_5556));
 AOI211xp5_ASAP7_75t_L g214862 (.A1(n_1772),
    .A2(n_2390),
    .B(n_3185),
    .C(n_2244),
    .Y(n_5555));
 OAI22xp33_ASAP7_75t_L g214863 (.A1(n_4195),
    .A2(n_2081),
    .B1(n_1354),
    .B2(n_3253),
    .Y(n_5554));
 OAI32xp33_ASAP7_75t_L g214864 (.A1(n_3293),
    .A2(n_1429),
    .A3(n_2504),
    .B1(n_2080),
    .B2(n_4440),
    .Y(n_5553));
 AOI221xp5_ASAP7_75t_SL g214865 (.A1(n_4089),
    .A2(n_2777),
    .B1(n_3139),
    .B2(n_1353),
    .C(n_4171),
    .Y(n_5552));
 OAI221xp5_ASAP7_75t_SL g214866 (.A1(n_2780),
    .A2(n_4070),
    .B1(n_3722),
    .B2(n_1461),
    .C(n_4134),
    .Y(n_5551));
 AOI22xp33_ASAP7_75t_R g214867 (.A1(n_4186),
    .A2(n_1423),
    .B1(n_3248),
    .B2(n_1444),
    .Y(n_5550));
 AO22x1_ASAP7_75t_SL g214868 (.A1(n_1372),
    .A2(n_4059),
    .B1(n_2040),
    .B2(n_2806),
    .Y(n_5549));
 AOI22xp33_ASAP7_75t_R g214869 (.A1(n_1370),
    .A2(n_4045),
    .B1(n_2077),
    .B2(n_3244),
    .Y(n_5548));
 AOI221xp5_ASAP7_75t_R g214870 (.A1(n_2906),
    .A2(n_1460),
    .B1(n_4653),
    .B2(n_1653),
    .C(n_2183),
    .Y(n_5547));
 AOI22xp33_ASAP7_75t_L g214871 (.A1(n_4050),
    .A2(n_2072),
    .B1(n_2786),
    .B2(n_1542),
    .Y(n_5546));
 AOI22xp33_ASAP7_75t_R g214872 (.A1(n_1577),
    .A2(n_4173),
    .B1(n_2787),
    .B2(n_1419),
    .Y(n_5545));
 AOI22xp33_ASAP7_75t_R g214873 (.A1(n_1552),
    .A2(n_4611),
    .B1(n_2437),
    .B2(n_1664),
    .Y(n_5544));
 AOI221xp5_ASAP7_75t_R g214874 (.A1(n_3682),
    .A2(n_1689),
    .B1(n_3918),
    .B2(n_2130),
    .C(n_1510),
    .Y(n_5543));
 OAI22xp33_ASAP7_75t_R g214875 (.A1(n_4001),
    .A2(n_1418),
    .B1(n_3274),
    .B2(n_1582),
    .Y(n_5542));
 AOI22xp33_ASAP7_75t_R g214876 (.A1(n_1586),
    .A2(n_4024),
    .B1(n_1431),
    .B2(n_1726),
    .Y(n_5541));
 AOI32xp33_ASAP7_75t_R g214877 (.A1(n_2781),
    .A2(n_2397),
    .A3(n_2440),
    .B1(n_4623),
    .B2(n_2427),
    .Y(n_5540));
 AO32x1_ASAP7_75t_SL g214878 (.A1(n_1712),
    .A2(n_2389),
    .A3(n_2442),
    .B1(n_1772),
    .B2(n_2431),
    .Y(n_5539));
 OAI321xp33_ASAP7_75t_L g214879 (.A1(n_3244),
    .A2(n_3290),
    .A3(n_2063),
    .B1(n_1454),
    .B2(n_3137),
    .C(n_4118),
    .Y(n_5538));
 OAI22xp33_ASAP7_75t_R g214880 (.A1(n_1580),
    .A2(n_3979),
    .B1(n_2793),
    .B2(n_2061),
    .Y(n_5537));
 AOI221xp5_ASAP7_75t_L g214881 (.A1(n_3937),
    .A2(n_1424),
    .B1(n_3659),
    .B2(n_1844),
    .C(n_4031),
    .Y(n_5536));
 INVxp67_ASAP7_75t_L g214882 (.A(n_5242),
    .Y(n_5533));
 INVxp67_ASAP7_75t_R g214883 (.A(n_5531),
    .Y(n_5532));
 INVxp33_ASAP7_75t_R g214884 (.A(n_5528),
    .Y(n_5529));
 INVxp33_ASAP7_75t_R g214886 (.A(n_5519),
    .Y(n_5520));
 INVxp67_ASAP7_75t_R g214887 (.A(n_5517),
    .Y(n_5518));
 INVxp67_ASAP7_75t_R g214888 (.A(n_5498),
    .Y(n_5499));
 INVxp67_ASAP7_75t_L g214889 (.A(n_5491),
    .Y(n_5492));
 INVxp67_ASAP7_75t_L g214890 (.A(n_5489),
    .Y(n_5490));
 INVxp67_ASAP7_75t_R g214891 (.A(n_5485),
    .Y(n_5486));
 INVxp67_ASAP7_75t_R g214892 (.A(n_5482),
    .Y(n_5483));
 INVxp33_ASAP7_75t_R g214893 (.A(n_5479),
    .Y(n_5480));
 INVxp67_ASAP7_75t_R g214894 (.A(n_5477),
    .Y(n_5478));
 INVx1_ASAP7_75t_L g214895 (.A(n_5473),
    .Y(n_5474));
 INVxp33_ASAP7_75t_R g214896 (.A(n_5468),
    .Y(n_5469));
 INVxp67_ASAP7_75t_R g214897 (.A(n_5466),
    .Y(n_5467));
 INVxp67_ASAP7_75t_R g214898 (.A(n_5464),
    .Y(n_5465));
 INVxp33_ASAP7_75t_R g214899 (.A(n_5459),
    .Y(n_5460));
 INVxp33_ASAP7_75t_R g214900 (.A(n_5449),
    .Y(n_5450));
 INVxp33_ASAP7_75t_R g214901 (.A(n_5447),
    .Y(n_5448));
 INVxp67_ASAP7_75t_R g214902 (.A(n_5435),
    .Y(n_5436));
 INVxp67_ASAP7_75t_L g214903 (.A(n_5433),
    .Y(n_5434));
 INVxp67_ASAP7_75t_R g214904 (.A(n_5430),
    .Y(n_5431));
 INVxp33_ASAP7_75t_R g214905 (.A(n_5425),
    .Y(n_5426));
 INVxp33_ASAP7_75t_R g214906 (.A(n_5422),
    .Y(n_5423));
 INVxp67_ASAP7_75t_L g214907 (.A(n_5419),
    .Y(n_5420));
 INVxp67_ASAP7_75t_L g214908 (.A(n_5418),
    .Y(n_5417));
 INVxp67_ASAP7_75t_R g214909 (.A(n_5412),
    .Y(n_5413));
 INVxp67_ASAP7_75t_R g214910 (.A(n_5409),
    .Y(n_5410));
 INVxp67_ASAP7_75t_SL g214911 (.A(n_5407),
    .Y(n_5408));
 INVxp67_ASAP7_75t_L g214913 (.A(n_5403),
    .Y(n_5404));
 INVxp67_ASAP7_75t_R g214915 (.A(n_1791),
    .Y(n_5402));
 INVx1_ASAP7_75t_R g214916 (.A(n_5400),
    .Y(n_5401));
 INVx1_ASAP7_75t_L g214917 (.A(n_5398),
    .Y(n_5399));
 INVxp67_ASAP7_75t_R g214918 (.A(n_5396),
    .Y(n_5395));
 INVxp67_ASAP7_75t_R g214919 (.A(n_5393),
    .Y(n_5392));
 INVxp67_ASAP7_75t_R g214920 (.A(n_5390),
    .Y(n_5391));
 INVxp67_ASAP7_75t_R g214922 (.A(n_1790),
    .Y(n_5389));
 INVx1_ASAP7_75t_SL g214923 (.A(n_5386),
    .Y(n_5387));
 INVxp67_ASAP7_75t_R g214924 (.A(n_5381),
    .Y(n_5382));
 INVxp33_ASAP7_75t_R g214925 (.A(n_5379),
    .Y(n_5380));
 INVxp67_ASAP7_75t_R g214926 (.A(n_5377),
    .Y(n_5376));
 INVxp33_ASAP7_75t_R g214927 (.A(n_5374),
    .Y(n_5375));
 OAI21xp33_ASAP7_75t_R g214928 (.A1(n_3158),
    .A2(n_2073),
    .B(n_2475),
    .Y(n_5373));
 NOR2xp33_ASAP7_75t_SL g214929 (.A(n_3595),
    .B(n_4555),
    .Y(n_5372));
 OAI221xp5_ASAP7_75t_R g214931 (.A1(n_3111),
    .A2(sa02[1]),
    .B1(n_2068),
    .B2(n_2293),
    .C(n_3681),
    .Y(n_5371));
 NOR2xp33_ASAP7_75t_R g214932 (.A(n_1634),
    .B(n_3861),
    .Y(n_5370));
 OR2x2_ASAP7_75t_L g214933 (.A(n_1647),
    .B(n_3869),
    .Y(n_5369));
 NOR2xp33_ASAP7_75t_R g214934 (.A(n_2724),
    .B(n_4585),
    .Y(n_5368));
 NAND2xp33_ASAP7_75t_L g214935 (.A(n_4157),
    .B(n_4574),
    .Y(n_5367));
 AOI21xp33_ASAP7_75t_R g214936 (.A1(n_3093),
    .A2(n_1667),
    .B(n_3543),
    .Y(n_5366));
 NOR2xp33_ASAP7_75t_L g214937 (.A(n_4540),
    .B(n_4199),
    .Y(n_5365));
 NAND2xp33_ASAP7_75t_L g214938 (.A(n_4529),
    .B(n_4149),
    .Y(n_5364));
 NOR2xp33_ASAP7_75t_R g214939 (.A(n_2714),
    .B(n_4697),
    .Y(n_5363));
 NAND2xp5_ASAP7_75t_L g214940 (.A(n_2730),
    .B(n_4639),
    .Y(n_5362));
 NAND2xp33_ASAP7_75t_R g214941 (.A(n_2729),
    .B(n_4679),
    .Y(n_5361));
 NAND2xp33_ASAP7_75t_R g214942 (.A(n_4672),
    .B(n_3702),
    .Y(n_5360));
 OR2x2_ASAP7_75t_R g214943 (.A(n_2339),
    .B(n_4398),
    .Y(n_5359));
 AND2x2_ASAP7_75t_R g214944 (.A(n_3399),
    .B(n_4556),
    .Y(n_5358));
 NOR2xp33_ASAP7_75t_R g214945 (.A(sa23[3]),
    .B(n_4056),
    .Y(n_5357));
 NOR2xp33_ASAP7_75t_L g214946 (.A(n_3503),
    .B(n_4309),
    .Y(n_5356));
 NOR2xp33_ASAP7_75t_R g214947 (.A(n_1364),
    .B(n_4367),
    .Y(n_5355));
 NOR2xp33_ASAP7_75t_R g214948 (.A(n_4614),
    .B(n_3924),
    .Y(n_5354));
 NAND2xp5_ASAP7_75t_L g214949 (.A(n_4488),
    .B(n_1783),
    .Y(n_5353));
 NAND2xp33_ASAP7_75t_R g214950 (.A(n_4704),
    .B(n_4134),
    .Y(n_5352));
 NOR2xp33_ASAP7_75t_SL g214951 (.A(n_8177),
    .B(n_3850),
    .Y(n_5351));
 OAI21xp33_ASAP7_75t_R g214952 (.A1(n_2078),
    .A2(n_3179),
    .B(n_2477),
    .Y(n_5350));
 NOR2xp33_ASAP7_75t_L g214953 (.A(n_2411),
    .B(n_3875),
    .Y(n_5349));
 NAND2xp33_ASAP7_75t_R g214954 (.A(n_2421),
    .B(n_3877),
    .Y(n_5348));
 NAND2xp33_ASAP7_75t_R g214955 (.A(n_4029),
    .B(n_1972),
    .Y(n_5347));
 NAND2xp33_ASAP7_75t_R g214956 (.A(n_1432),
    .B(n_1764),
    .Y(n_5346));
 NOR2xp33_ASAP7_75t_L g214957 (.A(n_3431),
    .B(n_4688),
    .Y(n_5345));
 NAND2xp33_ASAP7_75t_R g214958 (.A(n_1349),
    .B(n_3893),
    .Y(n_5344));
 OAI21xp33_ASAP7_75t_R g214959 (.A1(n_2068),
    .A2(n_3167),
    .B(n_2596),
    .Y(n_5343));
 AND2x2_ASAP7_75t_R g214960 (.A(n_1664),
    .B(n_3898),
    .Y(n_5342));
 OAI21xp33_ASAP7_75t_L g214961 (.A1(n_3356),
    .A2(n_3434),
    .B(n_2072),
    .Y(n_5341));
 AOI211xp5_ASAP7_75t_L g214962 (.A1(n_2055),
    .A2(n_1593),
    .B(n_4687),
    .C(sa00[0]),
    .Y(n_5340));
 OAI21xp33_ASAP7_75t_R g214963 (.A1(n_3216),
    .A2(n_2080),
    .B(n_2450),
    .Y(n_5339));
 OAI21xp33_ASAP7_75t_L g214964 (.A1(n_2070),
    .A2(n_3211),
    .B(n_2473),
    .Y(n_5338));
 AOI211xp5_ASAP7_75t_R g214965 (.A1(n_2077),
    .A2(n_2133),
    .B(n_4691),
    .C(sa12[0]),
    .Y(n_5337));
 NAND2xp33_ASAP7_75t_R g214966 (.A(sa22[3]),
    .B(n_1761),
    .Y(n_5336));
 OAI21xp33_ASAP7_75t_R g214967 (.A1(n_1590),
    .A2(n_3001),
    .B(n_2442),
    .Y(n_5335));
 AO21x1_ASAP7_75t_SL g214968 (.A1(n_2829),
    .A2(n_3702),
    .B(n_2363),
    .Y(n_5334));
 OAI21xp33_ASAP7_75t_R g214969 (.A1(n_2083),
    .A2(n_3210),
    .B(n_2485),
    .Y(n_5333));
 OR2x2_ASAP7_75t_L g214970 (.A(n_4382),
    .B(n_4093),
    .Y(n_5332));
 OAI211xp5_ASAP7_75t_L g214971 (.A1(n_2153),
    .A2(n_2057),
    .B(n_4520),
    .C(n_1877),
    .Y(n_5331));
 NOR2xp33_ASAP7_75t_R g214972 (.A(n_1860),
    .B(n_4198),
    .Y(n_5330));
 NOR2xp33_ASAP7_75t_R g214973 (.A(n_8210),
    .B(n_4197),
    .Y(n_5329));
 OAI21xp5_ASAP7_75t_SL g214974 (.A1(n_1501),
    .A2(n_3518),
    .B(n_3657),
    .Y(n_5328));
 AOI21xp33_ASAP7_75t_R g214975 (.A1(n_2095),
    .A2(n_2519),
    .B(n_4485),
    .Y(n_5327));
 NOR2xp33_ASAP7_75t_R g214976 (.A(n_2068),
    .B(n_3887),
    .Y(n_5326));
 NAND2xp33_ASAP7_75t_R g214977 (.A(n_2413),
    .B(n_4348),
    .Y(n_5325));
 NAND2xp33_ASAP7_75t_R g214978 (.A(n_2462),
    .B(n_4415),
    .Y(n_5324));
 AOI21xp33_ASAP7_75t_R g214979 (.A1(n_2537),
    .A2(n_2205),
    .B(n_4441),
    .Y(n_5323));
 AOI221xp5_ASAP7_75t_L g214980 (.A1(n_3637),
    .A2(n_2128),
    .B1(n_1444),
    .B2(n_2123),
    .C(sa02[0]),
    .Y(n_5322));
 AO21x1_ASAP7_75t_R g214981 (.A1(n_2178),
    .A2(n_2503),
    .B(n_4495),
    .Y(n_5321));
 AND2x2_ASAP7_75t_R g214982 (.A(n_2931),
    .B(n_3935),
    .Y(n_5320));
 OAI211xp5_ASAP7_75t_L g214983 (.A1(n_2107),
    .A2(n_1450),
    .B(n_4560),
    .C(n_8182),
    .Y(n_5319));
 NAND2xp33_ASAP7_75t_R g214984 (.A(n_1687),
    .B(n_4405),
    .Y(n_5318));
 AOI21xp33_ASAP7_75t_SL g214985 (.A1(n_2496),
    .A2(n_1605),
    .B(n_4484),
    .Y(n_5317));
 NOR2xp33_ASAP7_75t_R g214986 (.A(n_2041),
    .B(n_3898),
    .Y(n_5316));
 AOI21xp5_ASAP7_75t_L g214987 (.A1(n_2917),
    .A2(n_2095),
    .B(n_4641),
    .Y(n_5315));
 AND2x2_ASAP7_75t_R g214988 (.A(n_1550),
    .B(n_3898),
    .Y(n_5314));
 AOI211xp5_ASAP7_75t_L g214989 (.A1(n_1547),
    .A2(n_2146),
    .B(n_4564),
    .C(n_1866),
    .Y(n_5313));
 OA211x2_ASAP7_75t_L g214990 (.A1(n_2279),
    .A2(n_2415),
    .B(n_3477),
    .C(n_3112),
    .Y(n_5312));
 OAI21xp33_ASAP7_75t_R g214991 (.A1(n_1602),
    .A2(n_2533),
    .B(n_4498),
    .Y(n_5311));
 AOI21xp33_ASAP7_75t_R g214992 (.A1(n_2509),
    .A2(n_1603),
    .B(n_4493),
    .Y(n_5310));
 OAI21xp33_ASAP7_75t_L g214993 (.A1(n_1759),
    .A2(n_2393),
    .B(n_3578),
    .Y(n_5309));
 AND2x2_ASAP7_75t_L g214994 (.A(n_2500),
    .B(n_4380),
    .Y(n_5308));
 AOI21xp33_ASAP7_75t_R g214995 (.A1(n_1689),
    .A2(n_1595),
    .B(n_4497),
    .Y(n_5307));
 NAND3xp33_ASAP7_75t_R g214996 (.A(n_2796),
    .B(n_1439),
    .C(n_1532),
    .Y(n_5306));
 NAND2xp33_ASAP7_75t_R g214997 (.A(n_1682),
    .B(n_4372),
    .Y(n_5305));
 AOI21xp33_ASAP7_75t_R g214998 (.A1(n_8690),
    .A2(n_3640),
    .B(n_3661),
    .Y(n_5304));
 AOI211xp5_ASAP7_75t_R g214999 (.A1(n_2054),
    .A2(n_1601),
    .B(n_4627),
    .C(sa22[0]),
    .Y(n_5303));
 NOR2xp33_ASAP7_75t_R g215000 (.A(n_2447),
    .B(n_4337),
    .Y(n_5302));
 OAI21xp33_ASAP7_75t_R g215001 (.A1(n_3654),
    .A2(n_2052),
    .B(n_3674),
    .Y(n_5301));
 AOI211xp5_ASAP7_75t_R g215002 (.A1(n_1627),
    .A2(n_2253),
    .B(n_2832),
    .C(n_1968),
    .Y(n_5300));
 OAI21xp33_ASAP7_75t_R g215003 (.A1(n_3655),
    .A2(n_1442),
    .B(n_3618),
    .Y(n_5299));
 NAND2xp5_ASAP7_75t_L g215004 (.A(n_2427),
    .B(n_4358),
    .Y(n_5298));
 O2A1O1Ixp33_ASAP7_75t_R g215005 (.A1(n_1839),
    .A2(n_2540),
    .B(n_2415),
    .C(n_2924),
    .Y(n_5297));
 NAND2xp33_ASAP7_75t_R g215006 (.A(n_1343),
    .B(n_3854),
    .Y(n_5296));
 OAI211xp5_ASAP7_75t_R g215007 (.A1(n_2235),
    .A2(n_2399),
    .B(n_3283),
    .C(sa02[0]),
    .Y(n_5295));
 A2O1A1Ixp33_ASAP7_75t_R g215008 (.A1(n_1935),
    .A2(n_2212),
    .B(n_2394),
    .C(sa10[1]),
    .Y(n_5294));
 A2O1A1Ixp33_ASAP7_75t_R g215009 (.A1(n_1500),
    .A2(n_2524),
    .B(n_1627),
    .C(n_2923),
    .Y(n_5293));
 O2A1O1Ixp33_ASAP7_75t_R g215010 (.A1(n_1457),
    .A2(n_2521),
    .B(n_2399),
    .C(n_2930),
    .Y(n_5292));
 A2O1A1Ixp33_ASAP7_75t_L g215011 (.A1(n_1395),
    .A2(n_2501),
    .B(n_1398),
    .C(n_2936),
    .Y(n_5291));
 OAI211xp5_ASAP7_75t_SL g215012 (.A1(n_2186),
    .A2(n_2047),
    .B(n_4650),
    .C(n_1509),
    .Y(n_5290));
 OAI21xp33_ASAP7_75t_R g215013 (.A1(n_3164),
    .A2(n_3642),
    .B(n_4348),
    .Y(n_5289));
 A2O1A1Ixp33_ASAP7_75t_R g215014 (.A1(n_1455),
    .A2(n_2196),
    .B(n_1351),
    .C(sa12[1]),
    .Y(n_5288));
 NAND2xp5_ASAP7_75t_R g215015 (.A(n_1622),
    .B(n_4362),
    .Y(n_5287));
 NOR2xp33_ASAP7_75t_R g215016 (.A(n_1678),
    .B(n_4217),
    .Y(n_5286));
 A2O1A1Ixp33_ASAP7_75t_R g215017 (.A1(sa11[6]),
    .A2(n_2562),
    .B(n_1659),
    .C(n_2918),
    .Y(n_5285));
 O2A1O1Ixp33_ASAP7_75t_R g215018 (.A1(n_1499),
    .A2(n_2529),
    .B(n_1565),
    .C(n_2927),
    .Y(n_5284));
 OAI211xp5_ASAP7_75t_L g215019 (.A1(n_2249),
    .A2(n_2052),
    .B(n_3254),
    .C(n_1980),
    .Y(n_5283));
 OA21x2_ASAP7_75t_R g215020 (.A1(n_3320),
    .A2(n_3488),
    .B(n_2075),
    .Y(n_5282));
 A2O1A1Ixp33_ASAP7_75t_R g215021 (.A1(sa30[6]),
    .A2(n_2555),
    .B(n_1445),
    .C(n_2943),
    .Y(n_5281));
 OAI21xp33_ASAP7_75t_SL g215022 (.A1(n_1546),
    .A2(n_3515),
    .B(n_3575),
    .Y(n_5280));
 A2O1A1Ixp33_ASAP7_75t_L g215023 (.A1(sa31[6]),
    .A2(n_2567),
    .B(n_1643),
    .C(n_3530),
    .Y(n_5279));
 AOI21xp33_ASAP7_75t_R g215024 (.A1(n_3485),
    .A2(n_3321),
    .B(n_1337),
    .Y(n_5278));
 OAI211xp5_ASAP7_75t_R g215025 (.A1(n_1610),
    .A2(n_2396),
    .B(n_3257),
    .C(sa22[0]),
    .Y(n_5277));
 A2O1A1Ixp33_ASAP7_75t_R g215026 (.A1(n_1935),
    .A2(n_2506),
    .B(n_2394),
    .C(n_3593),
    .Y(n_5276));
 OAI211xp5_ASAP7_75t_SL g215027 (.A1(n_2503),
    .A2(n_2393),
    .B(n_1769),
    .C(n_3609),
    .Y(n_5275));
 A2O1A1Ixp33_ASAP7_75t_R g215028 (.A1(n_1463),
    .A2(n_2584),
    .B(n_2389),
    .C(n_2920),
    .Y(n_5274));
 OA21x2_ASAP7_75t_R g215029 (.A1(n_3386),
    .A2(n_3527),
    .B(n_2090),
    .Y(n_5273));
 NAND2xp33_ASAP7_75t_R g215030 (.A(n_1704),
    .B(n_4284),
    .Y(n_5272));
 NAND2xp33_ASAP7_75t_R g215031 (.A(n_2089),
    .B(n_4385),
    .Y(n_5271));
 O2A1O1Ixp33_ASAP7_75t_R g215032 (.A1(n_1456),
    .A2(n_2575),
    .B(n_8691),
    .C(n_1753),
    .Y(n_5270));
 AO21x1_ASAP7_75t_L g215033 (.A1(n_3370),
    .A2(n_3491),
    .B(n_2081),
    .Y(n_5269));
 NOR2xp33_ASAP7_75t_R g215034 (.A(n_2489),
    .B(n_4344),
    .Y(n_5268));
 NAND2xp5_ASAP7_75t_R g215035 (.A(n_1465),
    .B(n_4043),
    .Y(n_5267));
 NAND3xp33_ASAP7_75t_R g215036 (.A(n_1728),
    .B(n_3406),
    .C(n_1498),
    .Y(n_5266));
 NOR2xp33_ASAP7_75t_SL g215037 (.A(n_2620),
    .B(n_4279),
    .Y(n_5265));
 NOR2xp33_ASAP7_75t_R g215038 (.A(n_2634),
    .B(n_4278),
    .Y(n_5264));
 A2O1A1Ixp33_ASAP7_75t_L g215039 (.A1(n_1934),
    .A2(n_2554),
    .B(n_1436),
    .C(n_3505),
    .Y(n_5263));
 OAI21xp33_ASAP7_75t_R g215040 (.A1(n_3368),
    .A2(n_3535),
    .B(n_1391),
    .Y(n_5262));
 NAND2xp33_ASAP7_75t_R g215041 (.A(n_2410),
    .B(n_4365),
    .Y(n_5261));
 NAND2xp33_ASAP7_75t_R g215042 (.A(n_1775),
    .B(n_2490),
    .Y(n_5535));
 NAND2xp33_ASAP7_75t_R g215043 (.A(n_4317),
    .B(n_2436),
    .Y(n_5260));
 OR3x1_ASAP7_75t_L g215044 (.A(n_4282),
    .B(n_3602),
    .C(n_2617),
    .Y(n_5259));
 OAI211xp5_ASAP7_75t_R g215045 (.A1(n_2496),
    .A2(n_2399),
    .B(n_4007),
    .C(n_3630),
    .Y(n_5258));
 AOI21xp33_ASAP7_75t_R g215046 (.A1(n_3036),
    .A2(sa30[3]),
    .B(n_3445),
    .Y(n_5257));
 AO21x1_ASAP7_75t_R g215047 (.A1(n_2394),
    .A2(n_3664),
    .B(n_1527),
    .Y(n_5256));
 OAI221xp5_ASAP7_75t_R g215048 (.A1(n_1551),
    .A2(n_2308),
    .B1(n_2395),
    .B2(n_1871),
    .C(n_4689),
    .Y(n_5255));
 OA21x2_ASAP7_75t_R g215049 (.A1(n_3373),
    .A2(n_3489),
    .B(n_2089),
    .Y(n_5254));
 OA21x2_ASAP7_75t_R g215050 (.A1(n_3347),
    .A2(n_3514),
    .B(n_2084),
    .Y(n_5253));
 NOR2xp33_ASAP7_75t_L g215051 (.A(n_3261),
    .B(n_4316),
    .Y(n_5252));
 O2A1O1Ixp33_ASAP7_75t_R g215052 (.A1(n_1460),
    .A2(n_2585),
    .B(n_2419),
    .C(n_3465),
    .Y(n_5251));
 NAND2xp33_ASAP7_75t_R g215053 (.A(n_1432),
    .B(n_4503),
    .Y(n_5250));
 OAI21xp5_ASAP7_75t_R g215054 (.A1(n_1742),
    .A2(n_3487),
    .B(n_1572),
    .Y(n_5249));
 OAI21xp33_ASAP7_75t_R g215055 (.A1(n_1654),
    .A2(n_3710),
    .B(n_8196),
    .Y(n_5248));
 NOR2xp33_ASAP7_75t_L g215056 (.A(n_1674),
    .B(n_4303),
    .Y(n_5534));
 OA211x2_ASAP7_75t_R g215057 (.A1(n_2014),
    .A2(n_2415),
    .B(n_3112),
    .C(n_2931),
    .Y(n_5247));
 AOI21xp5_ASAP7_75t_R g215058 (.A1(n_3530),
    .A2(n_2386),
    .B(n_3650),
    .Y(n_5246));
 O2A1O1Ixp33_ASAP7_75t_R g215059 (.A1(n_2731),
    .A2(n_2538),
    .B(n_1498),
    .C(n_1981),
    .Y(n_5245));
 NOR2xp33_ASAP7_75t_R g215060 (.A(n_1358),
    .B(n_4492),
    .Y(n_5244));
 A2O1A1Ixp33_ASAP7_75t_R g215061 (.A1(n_2715),
    .A2(n_1691),
    .B(n_1464),
    .C(sa01[2]),
    .Y(n_5243));
 O2A1O1Ixp33_ASAP7_75t_L g215062 (.A1(n_8177),
    .A2(n_2271),
    .B(n_3197),
    .C(n_4552),
    .Y(n_5242));
 NOR2xp33_ASAP7_75t_R g215063 (.A(n_1541),
    .B(n_4491),
    .Y(n_5241));
 OA21x2_ASAP7_75t_R g215064 (.A1(n_1669),
    .A2(n_2921),
    .B(n_3545),
    .Y(n_5240));
 NAND2xp33_ASAP7_75t_R g215065 (.A(n_1683),
    .B(n_4498),
    .Y(n_5239));
 AOI21xp33_ASAP7_75t_R g215066 (.A1(n_1754),
    .A2(n_2413),
    .B(n_4177),
    .Y(n_5238));
 AO21x1_ASAP7_75t_R g215067 (.A1(n_3165),
    .A2(n_3653),
    .B(n_3864),
    .Y(n_5237));
 NOR2xp33_ASAP7_75t_SL g215068 (.A(n_4269),
    .B(n_4366),
    .Y(n_5236));
 A2O1A1Ixp33_ASAP7_75t_R g215069 (.A1(n_2726),
    .A2(n_2534),
    .B(n_1844),
    .C(sa22[2]),
    .Y(n_5235));
 OA21x2_ASAP7_75t_L g215070 (.A1(n_2329),
    .A2(n_2045),
    .B(n_4642),
    .Y(n_5234));
 AOI221xp5_ASAP7_75t_L g215071 (.A1(n_3215),
    .A2(n_2001),
    .B1(n_1352),
    .B2(n_2137),
    .C(n_1966),
    .Y(n_5233));
 OA21x2_ASAP7_75t_SL g215072 (.A1(n_2296),
    .A2(n_1546),
    .B(n_4654),
    .Y(n_5232));
 OAI21xp33_ASAP7_75t_R g215073 (.A1(n_3494),
    .A2(n_2948),
    .B(sa11[0]),
    .Y(n_5231));
 NOR2xp33_ASAP7_75t_SL g215074 (.A(n_3442),
    .B(n_4399),
    .Y(n_5230));
 OAI211xp5_ASAP7_75t_L g215075 (.A1(sa12[4]),
    .A2(n_1512),
    .B(n_4647),
    .C(n_1455),
    .Y(n_5229));
 NOR2xp33_ASAP7_75t_R g215076 (.A(n_2558),
    .B(n_4007),
    .Y(n_5228));
 OAI21xp33_ASAP7_75t_R g215077 (.A1(n_2934),
    .A2(n_3085),
    .B(sa30[0]),
    .Y(n_5227));
 OAI221xp5_ASAP7_75t_L g215078 (.A1(n_2448),
    .A2(n_1507),
    .B1(n_1343),
    .B2(n_1491),
    .C(n_4351),
    .Y(n_5226));
 OAI211xp5_ASAP7_75t_SL g215079 (.A1(n_1506),
    .A2(n_1519),
    .B(n_1787),
    .C(n_1934),
    .Y(n_5225));
 OAI211xp5_ASAP7_75t_SL g215080 (.A1(n_1954),
    .A2(n_1860),
    .B(n_1786),
    .C(n_1458),
    .Y(n_5224));
 OA211x2_ASAP7_75t_SL g215081 (.A1(n_1387),
    .A2(sa11[3]),
    .B(n_4659),
    .C(n_1377),
    .Y(n_5223));
 NOR2xp33_ASAP7_75t_R g215082 (.A(n_2421),
    .B(n_4354),
    .Y(n_5222));
 NAND2xp33_ASAP7_75t_R g215083 (.A(n_3276),
    .B(n_4300),
    .Y(n_5221));
 AOI211xp5_ASAP7_75t_L g215084 (.A1(n_1467),
    .A2(n_8200),
    .B(n_4655),
    .C(n_1845),
    .Y(n_5220));
 NOR2xp33_ASAP7_75t_L g215085 (.A(n_3412),
    .B(n_4306),
    .Y(n_5219));
 NOR2xp33_ASAP7_75t_R g215086 (.A(n_2387),
    .B(n_4360),
    .Y(n_5218));
 NOR2xp33_ASAP7_75t_R g215087 (.A(n_1667),
    .B(n_3863),
    .Y(n_5217));
 OAI31xp33_ASAP7_75t_R g215088 (.A1(n_2876),
    .A2(n_1867),
    .A3(n_1888),
    .B(n_2694),
    .Y(n_5216));
 NAND2xp33_ASAP7_75t_R g215089 (.A(n_3283),
    .B(n_4295),
    .Y(n_5215));
 NOR2xp33_ASAP7_75t_R g215090 (.A(n_1669),
    .B(n_3991),
    .Y(n_5214));
 NOR2xp33_ASAP7_75t_R g215091 (.A(n_1655),
    .B(n_3880),
    .Y(n_5213));
 NAND2xp5_ASAP7_75t_L g215092 (.A(n_2851),
    .B(n_4575),
    .Y(n_5212));
 NOR2xp33_ASAP7_75t_L g215093 (.A(n_1625),
    .B(n_3897),
    .Y(n_5211));
 O2A1O1Ixp33_ASAP7_75t_L g215094 (.A1(n_2015),
    .A2(n_2591),
    .B(n_2429),
    .C(sa11[0]),
    .Y(n_5210));
 NAND2xp33_ASAP7_75t_R g215095 (.A(n_1745),
    .B(n_4323),
    .Y(n_5209));
 OAI211xp5_ASAP7_75t_L g215096 (.A1(n_2299),
    .A2(n_2059),
    .B(n_4541),
    .C(n_3621),
    .Y(n_5208));
 NOR2xp33_ASAP7_75t_R g215097 (.A(n_2829),
    .B(n_3971),
    .Y(n_5207));
 OAI211xp5_ASAP7_75t_SL g215098 (.A1(sa30[3]),
    .A2(n_1375),
    .B(n_4662),
    .C(n_1367),
    .Y(n_5206));
 OAI211xp5_ASAP7_75t_L g215099 (.A1(n_1851),
    .A2(sa33[3]),
    .B(n_4682),
    .C(n_1346),
    .Y(n_5205));
 NOR2xp33_ASAP7_75t_L g215100 (.A(n_3407),
    .B(n_1773),
    .Y(n_5204));
 NAND2xp5_ASAP7_75t_R g215101 (.A(n_1439),
    .B(n_4083),
    .Y(n_5203));
 NAND2xp33_ASAP7_75t_R g215102 (.A(n_2092),
    .B(n_4660),
    .Y(n_5202));
 NAND2xp33_ASAP7_75t_R g215103 (.A(n_4346),
    .B(n_2420),
    .Y(n_5201));
 NAND2xp33_ASAP7_75t_R g215104 (.A(n_3341),
    .B(n_4284),
    .Y(n_5200));
 NAND2xp33_ASAP7_75t_R g215105 (.A(n_4205),
    .B(n_2044),
    .Y(n_5199));
 NAND2xp33_ASAP7_75t_R g215106 (.A(n_4364),
    .B(n_2357),
    .Y(n_5198));
 NAND2xp33_ASAP7_75t_R g215107 (.A(n_4045),
    .B(n_2077),
    .Y(n_5197));
 NOR2xp33_ASAP7_75t_R g215108 (.A(n_1379),
    .B(n_4593),
    .Y(n_5196));
 NAND2xp33_ASAP7_75t_R g215109 (.A(n_1582),
    .B(n_4355),
    .Y(n_5195));
 NAND2xp33_ASAP7_75t_R g215110 (.A(n_2444),
    .B(n_4018),
    .Y(n_5194));
 NAND2xp5_ASAP7_75t_L g215111 (.A(n_1433),
    .B(n_4112),
    .Y(n_5193));
 NOR2xp33_ASAP7_75t_R g215112 (.A(n_2434),
    .B(n_4342),
    .Y(n_5192));
 NAND2xp33_ASAP7_75t_R g215113 (.A(n_4516),
    .B(n_1453),
    .Y(n_5191));
 AND2x2_ASAP7_75t_R g215114 (.A(n_1444),
    .B(n_4186),
    .Y(n_5190));
 NAND2xp33_ASAP7_75t_R g215115 (.A(n_1446),
    .B(n_4350),
    .Y(n_5189));
 NAND2xp5_ASAP7_75t_R g215116 (.A(n_1398),
    .B(n_4511),
    .Y(n_5188));
 NAND2xp33_ASAP7_75t_R g215117 (.A(n_2355),
    .B(n_4354),
    .Y(n_5187));
 NOR2xp33_ASAP7_75t_R g215118 (.A(n_2778),
    .B(n_4285),
    .Y(n_5186));
 NAND2xp5_ASAP7_75t_L g215119 (.A(n_3329),
    .B(n_4156),
    .Y(n_5185));
 NAND2xp33_ASAP7_75t_R g215120 (.A(n_2352),
    .B(n_4360),
    .Y(n_5184));
 NOR2xp33_ASAP7_75t_R g215121 (.A(n_2158),
    .B(n_3963),
    .Y(n_5183));
 NOR2xp33_ASAP7_75t_L g215122 (.A(n_2088),
    .B(n_3996),
    .Y(n_5182));
 NAND2xp5_ASAP7_75t_L g215123 (.A(n_2061),
    .B(n_3885),
    .Y(n_5181));
 NOR2xp33_ASAP7_75t_SL g215124 (.A(n_1442),
    .B(n_4026),
    .Y(n_5180));
 NOR2xp33_ASAP7_75t_R g215125 (.A(n_1381),
    .B(n_4286),
    .Y(n_5179));
 NAND2xp5_ASAP7_75t_L g215126 (.A(n_2366),
    .B(n_3866),
    .Y(n_5178));
 NAND2xp33_ASAP7_75t_R g215127 (.A(n_1445),
    .B(n_4306),
    .Y(n_5177));
 NOR2xp33_ASAP7_75t_R g215128 (.A(n_2852),
    .B(n_3946),
    .Y(n_5176));
 NAND2xp33_ASAP7_75t_R g215129 (.A(n_2800),
    .B(n_3844),
    .Y(n_5175));
 NOR2xp33_ASAP7_75t_R g215130 (.A(n_2344),
    .B(n_3927),
    .Y(n_5174));
 NOR2xp33_ASAP7_75t_R g215131 (.A(n_4301),
    .B(n_8702),
    .Y(n_5173));
 NAND2xp5_ASAP7_75t_R g215132 (.A(n_2354),
    .B(n_3885),
    .Y(n_5172));
 NAND2xp5_ASAP7_75t_L g215133 (.A(n_1554),
    .B(n_3985),
    .Y(n_5171));
 NAND2xp33_ASAP7_75t_R g215134 (.A(n_2367),
    .B(n_3880),
    .Y(n_5170));
 NOR2xp33_ASAP7_75t_R g215135 (.A(n_2457),
    .B(n_3917),
    .Y(n_5169));
 NAND2xp5_ASAP7_75t_L g215136 (.A(n_2128),
    .B(n_1766),
    .Y(n_5168));
 OAI21xp33_ASAP7_75t_R g215137 (.A1(n_3241),
    .A2(n_2104),
    .B(n_1372),
    .Y(n_5167));
 NOR2xp33_ASAP7_75t_R g215138 (.A(n_2474),
    .B(n_3860),
    .Y(n_5166));
 NOR2xp33_ASAP7_75t_L g215139 (.A(n_2806),
    .B(n_1778),
    .Y(n_5165));
 NAND2xp33_ASAP7_75t_R g215140 (.A(n_2079),
    .B(n_4130),
    .Y(n_5164));
 NAND2xp5_ASAP7_75t_R g215141 (.A(n_1440),
    .B(n_3882),
    .Y(n_5163));
 NAND2xp5_ASAP7_75t_R g215142 (.A(n_2477),
    .B(n_3956),
    .Y(n_5162));
 NOR2xp33_ASAP7_75t_R g215143 (.A(n_2341),
    .B(n_3902),
    .Y(n_5161));
 NAND2xp33_ASAP7_75t_R g215144 (.A(n_3888),
    .B(n_1621),
    .Y(n_5160));
 OR2x2_ASAP7_75t_L g215145 (.A(n_2484),
    .B(n_3905),
    .Y(n_5159));
 NAND2xp33_ASAP7_75t_R g215146 (.A(n_3915),
    .B(n_2442),
    .Y(n_5158));
 NOR2xp33_ASAP7_75t_R g215147 (.A(n_1660),
    .B(n_4277),
    .Y(n_5157));
 NOR2xp33_ASAP7_75t_R g215148 (.A(n_2468),
    .B(n_3874),
    .Y(n_5156));
 NOR2xp33_ASAP7_75t_R g215149 (.A(n_2449),
    .B(n_3963),
    .Y(n_5155));
 NOR2xp33_ASAP7_75t_R g215150 (.A(n_1565),
    .B(n_4280),
    .Y(n_5154));
 NOR2xp33_ASAP7_75t_R g215151 (.A(n_2399),
    .B(n_4048),
    .Y(n_5153));
 NAND2xp5_ASAP7_75t_R g215152 (.A(n_2343),
    .B(n_3911),
    .Y(n_5152));
 NOR2xp33_ASAP7_75t_SL g215153 (.A(n_2868),
    .B(n_4290),
    .Y(n_5151));
 NOR2xp33_ASAP7_75t_L g215154 (.A(n_1429),
    .B(n_4496),
    .Y(n_5150));
 NAND2xp33_ASAP7_75t_R g215155 (.A(n_8690),
    .B(n_4039),
    .Y(n_5149));
 NOR2xp33_ASAP7_75t_R g215156 (.A(n_1382),
    .B(n_4375),
    .Y(n_5148));
 NOR2xp33_ASAP7_75t_L g215157 (.A(n_1640),
    .B(n_4494),
    .Y(n_5147));
 NAND2xp33_ASAP7_75t_R g215158 (.A(n_3926),
    .B(n_2450),
    .Y(n_5146));
 NOR2xp33_ASAP7_75t_R g215159 (.A(n_1558),
    .B(n_4508),
    .Y(n_5145));
 NAND2xp33_ASAP7_75t_R g215160 (.A(n_1641),
    .B(n_4206),
    .Y(n_5144));
 NAND2xp33_ASAP7_75t_R g215161 (.A(n_3944),
    .B(n_1659),
    .Y(n_5143));
 NAND2xp33_ASAP7_75t_R g215162 (.A(n_2416),
    .B(n_1767),
    .Y(n_5142));
 NAND2xp5_ASAP7_75t_R g215163 (.A(n_1411),
    .B(n_4325),
    .Y(n_5141));
 NOR2xp33_ASAP7_75t_R g215164 (.A(n_2335),
    .B(n_4423),
    .Y(n_5140));
 NOR2xp33_ASAP7_75t_R g215165 (.A(n_2353),
    .B(n_3936),
    .Y(n_5139));
 NOR2xp33_ASAP7_75t_R g215166 (.A(n_3303),
    .B(n_4334),
    .Y(n_5138));
 NAND2xp5_ASAP7_75t_R g215167 (.A(n_2371),
    .B(n_3890),
    .Y(n_5137));
 NOR2xp33_ASAP7_75t_R g215168 (.A(n_1337),
    .B(n_4411),
    .Y(n_5136));
 NAND2xp5_ASAP7_75t_R g215169 (.A(n_1399),
    .B(n_1776),
    .Y(n_5135));
 NAND2xp33_ASAP7_75t_R g215170 (.A(n_3253),
    .B(n_4324),
    .Y(n_5134));
 NAND2xp5_ASAP7_75t_L g215171 (.A(n_1449),
    .B(n_4345),
    .Y(n_5531));
 NOR2xp33_ASAP7_75t_SL g215172 (.A(n_1642),
    .B(n_3861),
    .Y(n_5530));
 NAND2xp5_ASAP7_75t_R g215173 (.A(n_4333),
    .B(n_4305),
    .Y(n_5528));
 NAND2xp5_ASAP7_75t_R g215174 (.A(n_4324),
    .B(n_4284),
    .Y(n_5527));
 NAND2xp5_ASAP7_75t_SL g215175 (.A(n_4326),
    .B(n_4280),
    .Y(n_5526));
 NAND2xp5_ASAP7_75t_R g215176 (.A(n_2416),
    .B(n_3868),
    .Y(n_5525));
 NAND2xp5_ASAP7_75t_L g215177 (.A(n_2400),
    .B(n_1780),
    .Y(n_5524));
 NOR2xp33_ASAP7_75t_SL g215178 (.A(n_1662),
    .B(n_3864),
    .Y(n_5523));
 NAND2xp5_ASAP7_75t_SL g215179 (.A(n_1775),
    .B(n_4328),
    .Y(n_1793));
 NAND2xp5_ASAP7_75t_R g215180 (.A(n_2392),
    .B(n_4346),
    .Y(n_5522));
 NAND2xp5_ASAP7_75t_R g215181 (.A(n_1777),
    .B(n_4318),
    .Y(n_5521));
 NAND2xp33_ASAP7_75t_R g215182 (.A(n_4369),
    .B(n_2389),
    .Y(n_5519));
 NAND2xp5_ASAP7_75t_L g215183 (.A(n_3970),
    .B(n_4300),
    .Y(n_5517));
 NOR2xp67_ASAP7_75t_L g215184 (.A(n_4330),
    .B(n_4313),
    .Y(n_5516));
 NOR2xp33_ASAP7_75t_SL g215185 (.A(n_1558),
    .B(n_4367),
    .Y(n_5133));
 NAND2xp5_ASAP7_75t_L g215186 (.A(n_4295),
    .B(n_3972),
    .Y(n_5515));
 NAND2xp5_ASAP7_75t_L g215187 (.A(n_2079),
    .B(n_4649),
    .Y(n_5514));
 NOR2xp33_ASAP7_75t_L g215188 (.A(n_4315),
    .B(n_3946),
    .Y(n_5513));
 NOR2xp33_ASAP7_75t_R g215189 (.A(n_3845),
    .B(n_4332),
    .Y(n_5132));
 NAND2xp5_ASAP7_75t_R g215190 (.A(n_1433),
    .B(n_4307),
    .Y(n_5512));
 NAND2xp33_ASAP7_75t_R g215191 (.A(n_4307),
    .B(n_4286),
    .Y(n_5131));
 NAND2xp5_ASAP7_75t_R g215192 (.A(n_2054),
    .B(n_4284),
    .Y(n_5511));
 NAND2xp5_ASAP7_75t_R g215193 (.A(n_1447),
    .B(n_4289),
    .Y(n_5510));
 NAND2xp5_ASAP7_75t_L g215194 (.A(n_2072),
    .B(n_4618),
    .Y(n_5509));
 NAND2xp33_ASAP7_75t_R g215195 (.A(n_4294),
    .B(n_2062),
    .Y(n_5508));
 NAND2xp5_ASAP7_75t_L g215196 (.A(n_4298),
    .B(n_4294),
    .Y(n_5507));
 NOR2xp33_ASAP7_75t_R g215197 (.A(n_1443),
    .B(n_4375),
    .Y(n_5130));
 NAND2xp5_ASAP7_75t_R g215198 (.A(n_1422),
    .B(n_4394),
    .Y(n_5506));
 NAND2xp5_ASAP7_75t_R g215199 (.A(n_1399),
    .B(n_1761),
    .Y(n_5505));
 NAND2xp5_ASAP7_75t_R g215200 (.A(n_1641),
    .B(n_3851),
    .Y(n_5504));
 NOR2xp33_ASAP7_75t_R g215201 (.A(n_3846),
    .B(n_4309),
    .Y(n_5129));
 NAND2xp5_ASAP7_75t_L g215202 (.A(n_2389),
    .B(n_3856),
    .Y(n_5503));
 NAND2xp33_ASAP7_75t_R g215203 (.A(n_3854),
    .B(n_2051),
    .Y(n_5502));
 NAND2xp5_ASAP7_75t_L g215204 (.A(n_3849),
    .B(n_2046),
    .Y(n_5501));
 NAND2xp5_ASAP7_75t_R g215205 (.A(n_1627),
    .B(n_4350),
    .Y(n_5500));
 NAND2xp5_ASAP7_75t_R g215206 (.A(n_1627),
    .B(n_3858),
    .Y(n_5498));
 NAND2xp5_ASAP7_75t_L g215207 (.A(n_3871),
    .B(sa23[3]),
    .Y(n_5497));
 NOR2xp33_ASAP7_75t_R g215208 (.A(n_1354),
    .B(n_3852),
    .Y(n_5128));
 NAND2xp5_ASAP7_75t_R g215209 (.A(n_1449),
    .B(n_4412),
    .Y(n_5496));
 NAND2xp33_ASAP7_75t_R g215210 (.A(n_1448),
    .B(n_3856),
    .Y(n_5127));
 NOR2xp33_ASAP7_75t_L g215211 (.A(n_3959),
    .B(n_4297),
    .Y(n_5495));
 NAND2xp5_ASAP7_75t_L g215212 (.A(n_1436),
    .B(n_1782),
    .Y(n_5494));
 NAND2xp5_ASAP7_75t_R g215213 (.A(n_2042),
    .B(n_3851),
    .Y(n_5493));
 NOR2xp67_ASAP7_75t_L g215214 (.A(n_1560),
    .B(n_3853),
    .Y(n_5491));
 NAND2xp5_ASAP7_75t_L g215215 (.A(n_2050),
    .B(n_4434),
    .Y(n_5489));
 NOR2xp67_ASAP7_75t_L g215216 (.A(n_1541),
    .B(n_3857),
    .Y(n_5488));
 NAND2xp5_ASAP7_75t_L g215217 (.A(n_1438),
    .B(n_3849),
    .Y(n_5487));
 NOR2xp33_ASAP7_75t_L g215218 (.A(n_1662),
    .B(n_4450),
    .Y(n_5485));
 NAND2xp33_ASAP7_75t_R g215219 (.A(n_1627),
    .B(n_4376),
    .Y(n_5484));
 OAI21xp5_ASAP7_75t_L g215220 (.A1(n_3245),
    .A2(n_2586),
    .B(n_1653),
    .Y(n_5482));
 NAND2xp33_ASAP7_75t_R g215221 (.A(n_8690),
    .B(n_4464),
    .Y(n_5481));
 NAND2xp33_ASAP7_75t_R g215222 (.A(n_4287),
    .B(n_4277),
    .Y(n_5126));
 NOR2xp33_ASAP7_75t_R g215223 (.A(n_4296),
    .B(n_4282),
    .Y(n_5125));
 NOR2xp33_ASAP7_75t_SL g215224 (.A(n_3320),
    .B(n_4282),
    .Y(n_5479));
 NOR2xp33_ASAP7_75t_L g215225 (.A(n_3337),
    .B(n_4278),
    .Y(n_5477));
 NOR2xp33_ASAP7_75t_R g215226 (.A(n_2415),
    .B(n_4404),
    .Y(n_5124));
 NAND2xp5_ASAP7_75t_L g215227 (.A(n_1734),
    .B(n_4289),
    .Y(n_5476));
 NAND2xp5_ASAP7_75t_L g215228 (.A(n_1643),
    .B(n_4456),
    .Y(n_5475));
 NOR2x1_ASAP7_75t_L g215229 (.A(n_4299),
    .B(n_4303),
    .Y(n_5473));
 NAND2xp33_ASAP7_75t_R g215230 (.A(n_4301),
    .B(n_4291),
    .Y(n_5123));
 NAND2xp33_ASAP7_75t_R g215231 (.A(n_1741),
    .B(n_4294),
    .Y(n_5472));
 NOR2xp33_ASAP7_75t_L g215232 (.A(n_3356),
    .B(n_4309),
    .Y(n_5471));
 NOR2xp33_ASAP7_75t_R g215233 (.A(n_1640),
    .B(n_4443),
    .Y(n_5470));
 NAND2xp33_ASAP7_75t_R g215234 (.A(n_4314),
    .B(n_4289),
    .Y(n_5122));
 NAND2xp5_ASAP7_75t_R g215235 (.A(n_1552),
    .B(n_4668),
    .Y(n_5468));
 NAND2xp5_ASAP7_75t_L g215236 (.A(n_3367),
    .B(n_4307),
    .Y(n_5466));
 NOR2xp33_ASAP7_75t_L g215237 (.A(n_3330),
    .B(n_4303),
    .Y(n_5464));
 NAND2xp5_ASAP7_75t_SL g215238 (.A(n_3844),
    .B(n_4126),
    .Y(n_5463));
 NAND2xp5_ASAP7_75t_SL g215239 (.A(n_1735),
    .B(n_4301),
    .Y(n_5462));
 NAND2xp5_ASAP7_75t_R g215240 (.A(n_4323),
    .B(n_3321),
    .Y(n_5461));
 NAND2xp5_ASAP7_75t_R g215241 (.A(n_1638),
    .B(n_4489),
    .Y(n_5459));
 NOR2xp33_ASAP7_75t_L g215242 (.A(n_3386),
    .B(n_4279),
    .Y(n_5458));
 NOR2xp67_ASAP7_75t_L g215243 (.A(n_2430),
    .B(n_4668),
    .Y(n_5457));
 NOR2xp33_ASAP7_75t_L g215244 (.A(n_3373),
    .B(n_4332),
    .Y(n_5456));
 NAND2xp5_ASAP7_75t_R g215245 (.A(n_3346),
    .B(n_4319),
    .Y(n_5455));
 NOR2xp33_ASAP7_75t_R g215246 (.A(n_3349),
    .B(n_4313),
    .Y(n_5454));
 NOR2xp33_ASAP7_75t_SL g215247 (.A(n_3355),
    .B(n_4304),
    .Y(n_5453));
 NAND2xp33_ASAP7_75t_R g215248 (.A(n_4317),
    .B(n_4323),
    .Y(n_5121));
 NOR2xp33_ASAP7_75t_R g215249 (.A(n_1556),
    .B(n_4504),
    .Y(n_5452));
 NAND2xp5_ASAP7_75t_R g215250 (.A(n_1641),
    .B(n_4362),
    .Y(n_5120));
 NAND2xp5_ASAP7_75t_L g215251 (.A(n_1419),
    .B(n_4524),
    .Y(n_5451));
 NOR2xp33_ASAP7_75t_R g215252 (.A(n_1647),
    .B(n_4524),
    .Y(n_5449));
 NAND2xp33_ASAP7_75t_R g215253 (.A(n_1775),
    .B(n_1743),
    .Y(n_5447));
 NOR2x1_ASAP7_75t_L g215254 (.A(n_2396),
    .B(n_4359),
    .Y(n_5446));
 AOI21xp5_ASAP7_75t_SL g215255 (.A1(n_3275),
    .A2(n_1953),
    .B(n_2482),
    .Y(n_5445));
 NAND2xp33_ASAP7_75t_R g215256 (.A(n_1699),
    .B(n_4307),
    .Y(n_5119));
 NAND2xp5_ASAP7_75t_R g215257 (.A(n_2042),
    .B(n_4567),
    .Y(n_5444));
 NAND2xp33_ASAP7_75t_R g215258 (.A(n_1622),
    .B(n_4568),
    .Y(n_5118));
 NAND2xp5_ASAP7_75t_L g215259 (.A(n_1545),
    .B(n_4569),
    .Y(n_5443));
 NOR2xp33_ASAP7_75t_SL g215260 (.A(n_2424),
    .B(n_4569),
    .Y(n_5442));
 NAND2xp5_ASAP7_75t_L g215261 (.A(n_1655),
    .B(n_4580),
    .Y(n_5441));
 NAND2xp5_ASAP7_75t_L g215262 (.A(n_2044),
    .B(n_4579),
    .Y(n_5440));
 NAND2xp33_ASAP7_75t_R g215263 (.A(n_2387),
    .B(n_4573),
    .Y(n_5117));
 NAND2xp5_ASAP7_75t_L g215264 (.A(n_2040),
    .B(n_4572),
    .Y(n_5439));
 NAND2xp5_ASAP7_75t_L g215265 (.A(n_8690),
    .B(n_4348),
    .Y(n_5438));
 AOI21xp5_ASAP7_75t_R g215266 (.A1(n_2792),
    .A2(n_8189),
    .B(n_2484),
    .Y(n_5437));
 NAND2xp5_ASAP7_75t_L g215267 (.A(n_1432),
    .B(n_4584),
    .Y(n_5116));
 NAND2xp5_ASAP7_75t_R g215268 (.A(n_4583),
    .B(n_1439),
    .Y(n_5435));
 NOR2xp33_ASAP7_75t_SL g215269 (.A(n_1565),
    .B(n_4352),
    .Y(n_5433));
 NAND2xp5_ASAP7_75t_R g215270 (.A(n_2643),
    .B(n_4305),
    .Y(n_5432));
 OAI21xp5_ASAP7_75t_L g215271 (.A1(n_1503),
    .A2(n_2817),
    .B(n_2475),
    .Y(n_5430));
 AOI21xp33_ASAP7_75t_R g215272 (.A1(n_3251),
    .A2(n_1505),
    .B(n_2451),
    .Y(n_5115));
 NOR2x1_ASAP7_75t_R g215273 (.A(n_2478),
    .B(n_4382),
    .Y(n_5429));
 NOR2xp33_ASAP7_75t_L g215274 (.A(n_2423),
    .B(n_4602),
    .Y(n_5428));
 NAND2xp5_ASAP7_75t_R g215275 (.A(n_1431),
    .B(n_4602),
    .Y(n_5427));
 OAI21xp5_ASAP7_75t_L g215276 (.A1(sa23[4]),
    .A2(n_3266),
    .B(n_2469),
    .Y(n_5425));
 NOR2xp33_ASAP7_75t_L g215277 (.A(n_2434),
    .B(n_4622),
    .Y(n_5114));
 NAND2xp5_ASAP7_75t_L g215278 (.A(n_1444),
    .B(n_4622),
    .Y(n_5424));
 OAI21xp33_ASAP7_75t_R g215279 (.A1(sa22[4]),
    .A2(n_2782),
    .B(n_2440),
    .Y(n_5113));
 OAI21xp5_ASAP7_75t_L g215280 (.A1(n_1425),
    .A2(n_1732),
    .B(n_2456),
    .Y(n_5422));
 NAND2xp5_ASAP7_75t_SL g215281 (.A(n_1559),
    .B(n_4629),
    .Y(n_5421));
 NAND2xp5_ASAP7_75t_L g215282 (.A(n_1349),
    .B(n_4630),
    .Y(n_5419));
 OAI21xp5_ASAP7_75t_R g215283 (.A1(n_1387),
    .A2(n_2814),
    .B(n_2473),
    .Y(n_5418));
 NOR2xp33_ASAP7_75t_R g215284 (.A(n_2056),
    .B(n_1340),
    .Y(n_5416));
 NOR2xp33_ASAP7_75t_L g215285 (.A(n_1408),
    .B(n_4620),
    .Y(n_5415));
 NOR2xp33_ASAP7_75t_R g215286 (.A(n_2486),
    .B(n_4371),
    .Y(n_5414));
 AOI21xp33_ASAP7_75t_R g215287 (.A1(n_2784),
    .A2(n_8912),
    .B(n_2449),
    .Y(n_5112));
 NAND2xp5_ASAP7_75t_R g215288 (.A(n_4628),
    .B(n_2414),
    .Y(n_5412));
 AND2x2_ASAP7_75t_R g215289 (.A(n_2452),
    .B(n_4380),
    .Y(n_5411));
 NOR2xp33_ASAP7_75t_R g215290 (.A(n_1582),
    .B(n_4628),
    .Y(n_5409));
 NAND2xp5_ASAP7_75t_L g215291 (.A(n_1653),
    .B(n_4365),
    .Y(n_5407));
 AOI21xp33_ASAP7_75t_L g215292 (.A1(n_2803),
    .A2(n_8212),
    .B(n_2438),
    .Y(n_5406));
 NAND2xp5_ASAP7_75t_SL g215293 (.A(sa11[3]),
    .B(n_3987),
    .Y(n_5405));
 NOR2xp67_ASAP7_75t_L g215294 (.A(n_2660),
    .B(n_4313),
    .Y(n_1792));
 NAND2xp5_ASAP7_75t_SL g215295 (.A(n_1512),
    .B(n_4001),
    .Y(n_5403));
 NOR2xp67_ASAP7_75t_L g215296 (.A(n_1706),
    .B(n_4321),
    .Y(n_1791));
 NAND2xp5_ASAP7_75t_SL g215297 (.A(n_2645),
    .B(n_4323),
    .Y(n_5400));
 OA21x2_ASAP7_75t_SL g215298 (.A1(n_2438),
    .A2(n_3418),
    .B(n_1860),
    .Y(n_5398));
 NOR2x1_ASAP7_75t_SL g215299 (.A(n_1518),
    .B(n_4024),
    .Y(n_5397));
 AND2x2_ASAP7_75t_SL g215300 (.A(sa33[3]),
    .B(n_3979),
    .Y(n_5396));
 NOR2xp67_ASAP7_75t_L g215301 (.A(n_2636),
    .B(n_4309),
    .Y(n_5394));
 NAND2xp5_ASAP7_75t_L g215302 (.A(n_4324),
    .B(n_3257),
    .Y(n_5393));
 NAND2xp5_ASAP7_75t_R g215303 (.A(n_2675),
    .B(n_1775),
    .Y(n_5390));
 NOR2x1_ASAP7_75t_SL g215304 (.A(n_1707),
    .B(n_4302),
    .Y(n_1790));
 NOR2xp67_ASAP7_75t_L g215305 (.A(n_8181),
    .B(n_4006),
    .Y(n_5388));
 NOR2x1_ASAP7_75t_SL g215306 (.A(n_1467),
    .B(n_3989),
    .Y(n_5386));
 NAND2xp5_ASAP7_75t_L g215307 (.A(sa20[3]),
    .B(n_1771),
    .Y(n_5385));
 AND2x2_ASAP7_75t_L g215308 (.A(n_3284),
    .B(n_4317),
    .Y(n_5384));
 NAND2xp5_ASAP7_75t_L g215309 (.A(n_2833),
    .B(n_3847),
    .Y(n_5383));
 NOR2x1_ASAP7_75t_R g215310 (.A(n_3327),
    .B(n_4330),
    .Y(n_5381));
 NOR2x1_ASAP7_75t_L g215311 (.A(n_2856),
    .B(n_1778),
    .Y(n_5379));
 NAND2xp5_ASAP7_75t_L g215312 (.A(n_3246),
    .B(n_4328),
    .Y(n_5378));
 NOR2x1_ASAP7_75t_SL g215313 (.A(n_3255),
    .B(n_4325),
    .Y(n_5377));
 AND2x2_ASAP7_75t_L g215314 (.A(n_3324),
    .B(n_4333),
    .Y(n_5374));
 INVx1_ASAP7_75t_L g215315 (.A(n_4914),
    .Y(n_5110));
 INVxp67_ASAP7_75t_R g215316 (.A(n_4853),
    .Y(n_5109));
 INVxp67_ASAP7_75t_L g215317 (.A(n_5101),
    .Y(n_5102));
 INVxp67_ASAP7_75t_R g215319 (.A(n_5093),
    .Y(n_5094));
 INVxp67_ASAP7_75t_R g215320 (.A(n_5091),
    .Y(n_5092));
 INVxp67_ASAP7_75t_R g215321 (.A(n_5089),
    .Y(n_5090));
 INVxp67_ASAP7_75t_R g215322 (.A(n_5080),
    .Y(n_5081));
 INVxp33_ASAP7_75t_R g215323 (.A(n_5078),
    .Y(n_5079));
 INVxp67_ASAP7_75t_R g215324 (.A(n_5073),
    .Y(n_5074));
 INVxp67_ASAP7_75t_R g215325 (.A(n_5070),
    .Y(n_5071));
 INVxp67_ASAP7_75t_R g215326 (.A(n_5066),
    .Y(n_5067));
 INVxp33_ASAP7_75t_R g215327 (.A(n_5061),
    .Y(n_5062));
 INVxp33_ASAP7_75t_R g215329 (.A(n_5059),
    .Y(n_5060));
 INVxp33_ASAP7_75t_R g215330 (.A(n_5057),
    .Y(n_5058));
 INVxp67_ASAP7_75t_R g215331 (.A(n_5055),
    .Y(n_5056));
 INVxp33_ASAP7_75t_R g215332 (.A(n_5053),
    .Y(n_5054));
 INVxp67_ASAP7_75t_R g215333 (.A(n_5051),
    .Y(n_5052));
 INVxp67_ASAP7_75t_R g215334 (.A(n_5049),
    .Y(n_5050));
 INVxp67_ASAP7_75t_L g215335 (.A(n_5048),
    .Y(n_5047));
 OA21x2_ASAP7_75t_L g215336 (.A1(n_1647),
    .A2(n_3088),
    .B(n_3548),
    .Y(n_5046));
 OA21x2_ASAP7_75t_SL g215337 (.A1(n_2424),
    .A2(n_3143),
    .B(n_3559),
    .Y(n_5045));
 AOI22xp33_ASAP7_75t_L g215338 (.A1(n_1446),
    .A2(n_3003),
    .B1(n_2826),
    .B2(n_1545),
    .Y(n_5044));
 AOI21xp5_ASAP7_75t_R g215339 (.A1(n_3115),
    .A2(n_1625),
    .B(n_3074),
    .Y(n_5043));
 OAI21xp33_ASAP7_75t_R g215340 (.A1(n_3297),
    .A2(n_3602),
    .B(n_2369),
    .Y(n_5042));
 OAI21xp33_ASAP7_75t_L g215341 (.A1(n_2428),
    .A2(n_3099),
    .B(n_3557),
    .Y(n_5041));
 NAND3xp33_ASAP7_75t_R g215342 (.A(n_4415),
    .B(n_3308),
    .C(n_2414),
    .Y(n_5040));
 OAI22xp33_ASAP7_75t_L g215343 (.A1(n_2998),
    .A2(n_1382),
    .B1(n_3361),
    .B2(n_1354),
    .Y(n_5039));
 NAND3xp33_ASAP7_75t_L g215344 (.A(n_3310),
    .B(n_2420),
    .C(n_4408),
    .Y(n_5038));
 OAI21xp33_ASAP7_75t_L g215345 (.A1(n_2083),
    .A2(n_3605),
    .B(n_2615),
    .Y(n_5037));
 AO21x1_ASAP7_75t_R g215346 (.A1(n_1609),
    .A2(n_3415),
    .B(n_1971),
    .Y(n_5036));
 AO22x1_ASAP7_75t_L g215347 (.A1(n_1569),
    .A2(n_3076),
    .B1(n_1559),
    .B2(n_2855),
    .Y(n_5035));
 AO21x1_ASAP7_75t_R g215348 (.A1(n_1439),
    .A2(n_3483),
    .B(n_3951),
    .Y(n_5034));
 AOI22xp33_ASAP7_75t_R g215349 (.A1(n_2431),
    .A2(n_3042),
    .B1(n_1448),
    .B2(n_2830),
    .Y(n_5111));
 AOI22xp5_ASAP7_75t_R g215350 (.A1(n_3056),
    .A2(n_1625),
    .B1(n_2860),
    .B2(n_2042),
    .Y(n_5033));
 NOR3xp33_ASAP7_75t_L g215351 (.A(n_4402),
    .B(n_3279),
    .C(n_2428),
    .Y(n_5032));
 AOI22xp33_ASAP7_75t_R g215352 (.A1(n_2427),
    .A2(n_3369),
    .B1(n_3361),
    .B2(n_1424),
    .Y(n_5031));
 AOI211xp5_ASAP7_75t_R g215353 (.A1(n_2803),
    .A2(n_8212),
    .B(n_3301),
    .C(n_2434),
    .Y(n_5030));
 AO22x1_ASAP7_75t_R g215354 (.A1(n_3541),
    .A2(n_1664),
    .B1(n_3313),
    .B2(n_1549),
    .Y(n_5029));
 OAI21xp33_ASAP7_75t_R g215355 (.A1(n_1450),
    .A2(n_2843),
    .B(sa11[0]),
    .Y(n_5028));
 AOI21xp33_ASAP7_75t_L g215356 (.A1(n_2993),
    .A2(n_2069),
    .B(sa11[0]),
    .Y(n_5027));
 O2A1O1Ixp33_ASAP7_75t_R g215357 (.A1(n_1938),
    .A2(n_2271),
    .B(n_2078),
    .C(n_2323),
    .Y(n_5026));
 OAI22xp33_ASAP7_75t_R g215358 (.A1(n_1632),
    .A2(n_3605),
    .B1(n_1546),
    .B2(n_2857),
    .Y(n_5025));
 AOI32xp33_ASAP7_75t_L g215359 (.A1(n_2790),
    .A2(n_1445),
    .A3(n_2477),
    .B1(n_3070),
    .B2(n_2777),
    .Y(n_5024));
 OAI32xp33_ASAP7_75t_L g215360 (.A1(n_2802),
    .A2(n_2399),
    .A3(n_2438),
    .B1(n_3248),
    .B2(n_2977),
    .Y(n_5023));
 AOI22xp33_ASAP7_75t_R g215361 (.A1(n_2420),
    .A2(n_3104),
    .B1(n_2299),
    .B2(n_1431),
    .Y(n_5022));
 OAI22xp33_ASAP7_75t_L g215362 (.A1(n_1647),
    .A2(n_2925),
    .B1(n_1380),
    .B2(n_3168),
    .Y(n_5021));
 AOI21xp5_ASAP7_75t_R g215363 (.A1(n_3047),
    .A2(n_2509),
    .B(n_4612),
    .Y(n_5020));
 OAI211xp5_ASAP7_75t_R g215364 (.A1(n_1425),
    .A2(n_1732),
    .B(n_3314),
    .C(n_2065),
    .Y(n_5019));
 A2O1A1Ixp33_ASAP7_75t_R g215365 (.A1(n_1463),
    .A2(n_2256),
    .B(n_2087),
    .C(n_2331),
    .Y(n_5018));
 NOR2xp33_ASAP7_75t_R g215366 (.A(n_4255),
    .B(n_3930),
    .Y(n_5017));
 A2O1A1Ixp33_ASAP7_75t_R g215367 (.A1(n_1497),
    .A2(n_2228),
    .B(n_2089),
    .C(n_2305),
    .Y(n_5016));
 A2O1A1Ixp33_ASAP7_75t_R g215368 (.A1(n_1336),
    .A2(n_2252),
    .B(n_2072),
    .C(n_2312),
    .Y(n_5015));
 A2O1A1Ixp33_ASAP7_75t_R g215369 (.A1(n_1395),
    .A2(n_1610),
    .B(n_2082),
    .C(n_2309),
    .Y(n_5014));
 O2A1O1Ixp33_ASAP7_75t_SL g215370 (.A1(n_1671),
    .A2(n_2552),
    .B(n_1433),
    .C(n_3352),
    .Y(n_5013));
 AO21x1_ASAP7_75t_R g215371 (.A1(n_3290),
    .A2(n_3712),
    .B(n_2359),
    .Y(n_5012));
 OAI22xp33_ASAP7_75t_R g215372 (.A1(n_1408),
    .A2(n_2987),
    .B1(n_2419),
    .B2(n_2966),
    .Y(n_5011));
 O2A1O1Ixp33_ASAP7_75t_R g215373 (.A1(n_1839),
    .A2(n_2275),
    .B(n_1578),
    .C(n_2304),
    .Y(n_5010));
 AOI21xp33_ASAP7_75t_R g215374 (.A1(n_2072),
    .A2(n_3003),
    .B(n_1700),
    .Y(n_5009));
 OAI22xp33_ASAP7_75t_R g215375 (.A1(n_2979),
    .A2(n_1651),
    .B1(n_8691),
    .B2(n_3000),
    .Y(n_5008));
 A2O1A1Ixp33_ASAP7_75t_R g215376 (.A1(sa11[6]),
    .A2(n_2227),
    .B(n_2069),
    .C(n_2330),
    .Y(n_5007));
 O2A1O1Ixp33_ASAP7_75t_R g215377 (.A1(n_1845),
    .A2(n_1612),
    .B(n_1571),
    .C(n_2315),
    .Y(n_5006));
 O2A1O1Ixp33_ASAP7_75t_R g215378 (.A1(n_8180),
    .A2(n_2212),
    .B(n_1363),
    .C(n_2308),
    .Y(n_5005));
 AOI21xp33_ASAP7_75t_R g215379 (.A1(n_2860),
    .A2(sa30[6]),
    .B(n_1445),
    .Y(n_5004));
 AOI22xp33_ASAP7_75t_R g215380 (.A1(n_2425),
    .A2(n_3356),
    .B1(n_2827),
    .B2(n_2072),
    .Y(n_5003));
 A2O1A1Ixp33_ASAP7_75t_R g215381 (.A1(sa31[6]),
    .A2(n_2243),
    .B(n_2084),
    .C(n_2297),
    .Y(n_5002));
 O2A1O1Ixp33_ASAP7_75t_R g215382 (.A1(n_1457),
    .A2(n_2234),
    .B(n_2074),
    .C(n_2293),
    .Y(n_5001));
 A2O1A1Ixp33_ASAP7_75t_R g215383 (.A1(n_2015),
    .A2(n_1986),
    .B(n_2842),
    .C(sa11[6]),
    .Y(n_5000));
 OAI21xp33_ASAP7_75t_R g215384 (.A1(n_1844),
    .A2(n_3361),
    .B(n_1442),
    .Y(n_4999));
 O2A1O1Ixp33_ASAP7_75t_L g215385 (.A1(n_1395),
    .A2(n_2141),
    .B(n_1354),
    .C(n_3280),
    .Y(n_4998));
 A2O1A1Ixp33_ASAP7_75t_R g215386 (.A1(n_1465),
    .A2(n_2564),
    .B(n_3180),
    .C(n_1670),
    .Y(n_4997));
 O2A1O1Ixp33_ASAP7_75t_L g215387 (.A1(sa11[6]),
    .A2(n_2187),
    .B(n_1450),
    .C(n_3379),
    .Y(n_4996));
 NAND2xp33_ASAP7_75t_R g215388 (.A(n_1680),
    .B(n_3821),
    .Y(n_4995));
 A2O1A1Ixp33_ASAP7_75t_R g215389 (.A1(sa30[6]),
    .A2(n_2551),
    .B(n_3187),
    .C(n_1673),
    .Y(n_4994));
 A2O1A1Ixp33_ASAP7_75t_R g215390 (.A1(n_1460),
    .A2(n_2241),
    .B(n_2055),
    .C(n_3365),
    .Y(n_4993));
 O2A1O1Ixp33_ASAP7_75t_R g215391 (.A1(n_1456),
    .A2(n_2196),
    .B(n_2063),
    .C(n_2281),
    .Y(n_4992));
 AOI22xp33_ASAP7_75t_R g215392 (.A1(n_1655),
    .A2(n_2993),
    .B1(n_1659),
    .B2(n_3014),
    .Y(n_4991));
 AOI22xp33_ASAP7_75t_L g215393 (.A1(n_2392),
    .A2(n_3051),
    .B1(n_2231),
    .B2(n_1586),
    .Y(n_4990));
 OAI21xp33_ASAP7_75t_R g215394 (.A1(n_1501),
    .A2(n_2827),
    .B(n_1628),
    .Y(n_4989));
 O2A1O1Ixp33_ASAP7_75t_R g215395 (.A1(n_1404),
    .A2(n_2230),
    .B(n_2080),
    .C(n_2299),
    .Y(n_4988));
 AOI21xp5_ASAP7_75t_R g215396 (.A1(n_1350),
    .A2(n_3154),
    .B(n_2631),
    .Y(n_4987));
 AOI21xp33_ASAP7_75t_R g215397 (.A1(n_2829),
    .A2(n_1934),
    .B(n_1436),
    .Y(n_4986));
 OAI21xp5_ASAP7_75t_R g215398 (.A1(n_1457),
    .A2(n_3297),
    .B(n_1389),
    .Y(n_4985));
 OAI21xp33_ASAP7_75t_R g215399 (.A1(n_1464),
    .A2(n_2831),
    .B(n_1637),
    .Y(n_4984));
 OAI21xp33_ASAP7_75t_R g215400 (.A1(n_1499),
    .A2(n_1715),
    .B(n_1565),
    .Y(n_4983));
 OAI21xp33_ASAP7_75t_R g215401 (.A1(n_1460),
    .A2(n_2837),
    .B(n_2419),
    .Y(n_4982));
 AOI21xp5_ASAP7_75t_L g215402 (.A1(n_2858),
    .A2(sa31[6]),
    .B(n_2398),
    .Y(n_4981));
 A2O1A1Ixp33_ASAP7_75t_SL g215403 (.A1(n_1336),
    .A2(n_2574),
    .B(n_3192),
    .C(n_1677),
    .Y(n_4980));
 OAI21xp33_ASAP7_75t_R g215404 (.A1(n_1588),
    .A2(n_3041),
    .B(n_2603),
    .Y(n_4979));
 O2A1O1Ixp33_ASAP7_75t_L g215405 (.A1(sa30[6]),
    .A2(n_2168),
    .B(n_2043),
    .C(n_4068),
    .Y(n_4978));
 AOI21xp33_ASAP7_75t_L g215406 (.A1(n_1424),
    .A2(n_2997),
    .B(n_1696),
    .Y(n_4977));
 O2A1O1Ixp33_ASAP7_75t_L g215407 (.A1(n_1599),
    .A2(sa30[6]),
    .B(n_1390),
    .C(n_4306),
    .Y(n_4976));
 O2A1O1Ixp33_ASAP7_75t_R g215408 (.A1(n_1336),
    .A2(n_2143),
    .B(n_1543),
    .C(n_4002),
    .Y(n_4975));
 NAND3xp33_ASAP7_75t_R g215409 (.A(n_1581),
    .B(n_1693),
    .C(n_4294),
    .Y(n_4974));
 AO21x1_ASAP7_75t_R g215410 (.A1(n_2575),
    .A2(n_8703),
    .B(n_3924),
    .Y(n_4973));
 AOI21xp33_ASAP7_75t_R g215411 (.A1(n_2416),
    .A2(n_3030),
    .B(n_2164),
    .Y(n_4972));
 AO21x1_ASAP7_75t_R g215412 (.A1(n_2556),
    .A2(n_1641),
    .B(n_3941),
    .Y(n_4971));
 NOR3xp33_ASAP7_75t_R g215413 (.A(n_4282),
    .B(n_2074),
    .C(n_2617),
    .Y(n_4970));
 AOI21xp5_ASAP7_75t_R g215414 (.A1(n_2378),
    .A2(n_2854),
    .B(n_1938),
    .Y(n_4969));
 OA21x2_ASAP7_75t_L g215415 (.A1(n_2554),
    .A2(n_2393),
    .B(n_3925),
    .Y(n_4968));
 O2A1O1Ixp33_ASAP7_75t_L g215416 (.A1(n_2154),
    .A2(n_1465),
    .B(n_2057),
    .C(n_4290),
    .Y(n_4967));
 OAI22xp5_ASAP7_75t_L g215417 (.A1(n_1626),
    .A2(n_2943),
    .B1(n_2043),
    .B2(n_3161),
    .Y(n_4966));
 OAI21xp5_ASAP7_75t_L g215418 (.A1(n_3366),
    .A2(n_3245),
    .B(n_1461),
    .Y(n_4965));
 O2A1O1Ixp33_ASAP7_75t_R g215419 (.A1(n_1461),
    .A2(n_1593),
    .B(n_2056),
    .C(n_4310),
    .Y(n_4964));
 O2A1O1Ixp33_ASAP7_75t_L g215420 (.A1(n_2146),
    .A2(sa31[6]),
    .B(n_1548),
    .C(n_4320),
    .Y(n_4963));
 O2A1O1Ixp33_ASAP7_75t_L g215421 (.A1(n_2134),
    .A2(n_1336),
    .B(n_1543),
    .C(n_4309),
    .Y(n_4962));
 OA21x2_ASAP7_75t_L g215422 (.A1(n_1548),
    .A2(n_3242),
    .B(n_4151),
    .Y(n_4961));
 O2A1O1Ixp33_ASAP7_75t_R g215423 (.A1(n_1935),
    .A2(n_2099),
    .B(n_2041),
    .C(n_3992),
    .Y(n_4960));
 AOI21xp33_ASAP7_75t_R g215424 (.A1(n_2089),
    .A2(n_3556),
    .B(n_2600),
    .Y(n_4959));
 A2O1A1Ixp33_ASAP7_75t_L g215425 (.A1(n_1535),
    .A2(n_2534),
    .B(n_2396),
    .C(n_4009),
    .Y(n_4958));
 OAI21xp33_ASAP7_75t_R g215426 (.A1(n_1551),
    .A2(n_2971),
    .B(n_3942),
    .Y(n_4957));
 OAI21xp33_ASAP7_75t_R g215427 (.A1(n_2342),
    .A2(n_2825),
    .B(n_1465),
    .Y(n_4956));
 AO21x1_ASAP7_75t_R g215428 (.A1(n_2346),
    .A2(n_3289),
    .B(n_8180),
    .Y(n_4955));
 AOI21xp33_ASAP7_75t_R g215429 (.A1(n_3278),
    .A2(n_2337),
    .B(n_1844),
    .Y(n_4954));
 OAI21xp5_ASAP7_75t_R g215430 (.A1(n_3256),
    .A2(n_3280),
    .B(n_1395),
    .Y(n_4953));
 O2A1O1Ixp33_ASAP7_75t_R g215431 (.A1(n_2137),
    .A2(n_1934),
    .B(n_2059),
    .C(n_4303),
    .Y(n_4952));
 AOI22xp33_ASAP7_75t_R g215432 (.A1(n_2044),
    .A2(n_2815),
    .B1(n_1659),
    .B2(n_3219),
    .Y(n_4951));
 OAI21xp33_ASAP7_75t_R g215433 (.A1(n_2187),
    .A2(n_2881),
    .B(n_1659),
    .Y(n_4950));
 O2A1O1Ixp33_ASAP7_75t_R g215434 (.A1(n_1497),
    .A2(n_2131),
    .B(n_2047),
    .C(n_3999),
    .Y(n_4949));
 AO21x1_ASAP7_75t_R g215435 (.A1(n_2360),
    .A2(n_2845),
    .B(n_1499),
    .Y(n_4948));
 AOI21xp33_ASAP7_75t_R g215436 (.A1(n_3310),
    .A2(n_2374),
    .B(n_1403),
    .Y(n_4947));
 AOI21xp33_ASAP7_75t_R g215437 (.A1(n_3302),
    .A2(n_2380),
    .B(n_1459),
    .Y(n_4946));
 AOI21xp33_ASAP7_75t_R g215438 (.A1(n_2840),
    .A2(n_2382),
    .B(n_1839),
    .Y(n_4945));
 OAI21xp33_ASAP7_75t_R g215439 (.A1(n_2339),
    .A2(n_3315),
    .B(n_1497),
    .Y(n_4944));
 AOI21xp33_ASAP7_75t_R g215440 (.A1(n_3254),
    .A2(n_3287),
    .B(n_1499),
    .Y(n_4943));
 OA21x2_ASAP7_75t_L g215441 (.A1(n_1390),
    .A2(n_2789),
    .B(n_4157),
    .Y(n_4942));
 A2O1A1Ixp33_ASAP7_75t_R g215442 (.A1(n_1403),
    .A2(n_2174),
    .B(n_1431),
    .C(n_4125),
    .Y(n_4941));
 O2A1O1Ixp33_ASAP7_75t_R g215443 (.A1(n_1458),
    .A2(n_2129),
    .B(n_2068),
    .C(n_4114),
    .Y(n_4940));
 O2A1O1Ixp33_ASAP7_75t_R g215444 (.A1(n_1483),
    .A2(n_2507),
    .B(n_1653),
    .C(n_4005),
    .Y(n_4939));
 AND3x1_ASAP7_75t_R g215445 (.A(n_3450),
    .B(n_3329),
    .C(n_2346),
    .Y(n_4938));
 A2O1A1Ixp33_ASAP7_75t_L g215446 (.A1(n_2122),
    .A2(n_1459),
    .B(n_1444),
    .C(n_4281),
    .Y(n_4937));
 AOI22xp33_ASAP7_75t_R g215447 (.A1(n_1446),
    .A2(n_2922),
    .B1(n_1545),
    .B2(n_3217),
    .Y(n_4936));
 OAI21xp5_ASAP7_75t_R g215448 (.A1(n_2175),
    .A2(n_2874),
    .B(n_2392),
    .Y(n_4935));
 NAND3xp33_ASAP7_75t_L g215449 (.A(n_4394),
    .B(n_1740),
    .C(n_1423),
    .Y(n_4934));
 OA21x2_ASAP7_75t_L g215450 (.A1(n_2524),
    .A2(n_1629),
    .B(n_3945),
    .Y(n_4933));
 A2O1A1Ixp33_ASAP7_75t_L g215451 (.A1(n_1490),
    .A2(n_2537),
    .B(n_2052),
    .C(n_4014),
    .Y(n_4932));
 OAI21xp33_ASAP7_75t_L g215452 (.A1(n_2490),
    .A2(n_1408),
    .B(n_4526),
    .Y(n_4931));
 OAI21xp33_ASAP7_75t_L g215453 (.A1(n_2563),
    .A2(n_2825),
    .B(n_1447),
    .Y(n_4930));
 AOI21xp33_ASAP7_75t_R g215454 (.A1(n_3314),
    .A2(n_2579),
    .B(n_1378),
    .Y(n_4929));
 A2O1A1Ixp33_ASAP7_75t_L g215455 (.A1(n_1464),
    .A2(n_2223),
    .B(n_1447),
    .C(n_4073),
    .Y(n_4928));
 O2A1O1Ixp33_ASAP7_75t_R g215456 (.A1(sa12[7]),
    .A2(n_2510),
    .B(n_8690),
    .C(n_4022),
    .Y(n_4927));
 AOI21xp5_ASAP7_75t_R g215457 (.A1(n_3100),
    .A2(n_1440),
    .B(n_3921),
    .Y(n_4926));
 AO21x1_ASAP7_75t_L g215458 (.A1(n_1444),
    .A2(n_2803),
    .B(n_4192),
    .Y(n_4925));
 OAI21xp33_ASAP7_75t_R g215459 (.A1(n_2560),
    .A2(n_3307),
    .B(n_1547),
    .Y(n_4924));
 A2O1A1Ixp33_ASAP7_75t_L g215460 (.A1(n_8180),
    .A2(n_2211),
    .B(n_1550),
    .C(n_4323),
    .Y(n_4923));
 A2O1A1Ixp33_ASAP7_75t_SL g215461 (.A1(n_2167),
    .A2(n_1683),
    .B(n_2081),
    .C(n_3004),
    .Y(n_4922));
 NAND3xp33_ASAP7_75t_R g215462 (.A(n_3422),
    .B(n_2337),
    .C(n_3281),
    .Y(n_4921));
 OAI21xp33_ASAP7_75t_R g215463 (.A1(n_2591),
    .A2(n_2842),
    .B(n_2044),
    .Y(n_4920));
 A2O1A1Ixp33_ASAP7_75t_R g215464 (.A1(n_2205),
    .A2(n_2494),
    .B(n_2091),
    .C(n_2994),
    .Y(n_4919));
 A2O1A1Ixp33_ASAP7_75t_R g215465 (.A1(n_2444),
    .A2(n_1595),
    .B(n_2088),
    .C(n_3018),
    .Y(n_4918));
 O2A1O1Ixp33_ASAP7_75t_L g215466 (.A1(n_1455),
    .A2(n_2246),
    .B(n_1582),
    .C(n_3958),
    .Y(n_4917));
 OAI21xp33_ASAP7_75t_R g215467 (.A1(n_2544),
    .A2(n_3309),
    .B(n_2077),
    .Y(n_4916));
 A2O1A1Ixp33_ASAP7_75t_R g215468 (.A1(n_1485),
    .A2(n_2512),
    .B(n_1639),
    .C(n_4012),
    .Y(n_4915));
 A2O1A1Ixp33_ASAP7_75t_SL g215469 (.A1(n_2192),
    .A2(n_2490),
    .B(n_1342),
    .C(n_1721),
    .Y(n_4914));
 OA21x2_ASAP7_75t_L g215470 (.A1(n_3094),
    .A2(n_2396),
    .B(n_4183),
    .Y(n_4913));
 O2A1O1Ixp33_ASAP7_75t_L g215471 (.A1(n_2015),
    .A2(n_2520),
    .B(n_1659),
    .C(n_4011),
    .Y(n_4912));
 AOI22xp5_ASAP7_75t_R g215472 (.A1(n_3523),
    .A2(n_2065),
    .B1(n_3152),
    .B2(n_1439),
    .Y(n_4911));
 AOI21xp33_ASAP7_75t_R g215473 (.A1(n_2100),
    .A2(n_3429),
    .B(n_2395),
    .Y(n_4910));
 OAI21xp33_ASAP7_75t_R g215474 (.A1(n_2552),
    .A2(n_2853),
    .B(n_1435),
    .Y(n_4909));
 OAI22xp33_ASAP7_75t_R g215475 (.A1(n_2743),
    .A2(n_1669),
    .B1(n_2388),
    .B2(n_2584),
    .Y(n_4908));
 O2A1O1Ixp33_ASAP7_75t_R g215476 (.A1(n_2472),
    .A2(n_2096),
    .B(n_2069),
    .C(n_2937),
    .Y(n_4907));
 AOI21xp33_ASAP7_75t_R g215477 (.A1(n_2845),
    .A2(n_2545),
    .B(n_1560),
    .Y(n_4906));
 AOI21xp33_ASAP7_75t_R g215478 (.A1(n_2835),
    .A2(n_2574),
    .B(n_1544),
    .Y(n_4905));
 AOI21xp33_ASAP7_75t_R g215479 (.A1(n_2779),
    .A2(n_2589),
    .B(n_1408),
    .Y(n_4904));
 AO21x1_ASAP7_75t_R g215480 (.A1(n_1638),
    .A2(n_3170),
    .B(n_1785),
    .Y(n_4903));
 OA21x2_ASAP7_75t_SL g215481 (.A1(n_1381),
    .A2(n_2789),
    .B(n_2957),
    .Y(n_4902));
 O2A1O1Ixp33_ASAP7_75t_R g215482 (.A1(n_2198),
    .A2(n_2463),
    .B(n_2064),
    .C(n_3026),
    .Y(n_4901));
 O2A1O1Ixp33_ASAP7_75t_L g215483 (.A1(n_1525),
    .A2(n_2532),
    .B(n_2398),
    .C(n_4015),
    .Y(n_4900));
 OAI32xp33_ASAP7_75t_R g215484 (.A1(n_1418),
    .A2(n_1591),
    .A3(n_3290),
    .B1(n_1735),
    .B2(n_3072),
    .Y(n_4899));
 OAI21xp33_ASAP7_75t_R g215485 (.A1(n_2570),
    .A2(n_2787),
    .B(n_2404),
    .Y(n_4898));
 OAI21xp33_ASAP7_75t_R g215486 (.A1(n_3412),
    .A2(n_2778),
    .B(n_1625),
    .Y(n_4897));
 OAI21xp33_ASAP7_75t_R g215487 (.A1(n_2591),
    .A2(n_2804),
    .B(n_1655),
    .Y(n_4896));
 OAI22xp33_ASAP7_75t_R g215488 (.A1(n_2747),
    .A2(n_1632),
    .B1(n_2567),
    .B2(n_1644),
    .Y(n_4895));
 AOI21xp5_ASAP7_75t_R g215489 (.A1(n_2816),
    .A2(n_2072),
    .B(n_3002),
    .Y(n_4894));
 AO21x1_ASAP7_75t_R g215490 (.A1(n_1676),
    .A2(n_2421),
    .B(n_4601),
    .Y(n_4893));
 OR3x1_ASAP7_75t_R g215491 (.A(n_3448),
    .B(n_2852),
    .C(n_2342),
    .Y(n_4892));
 A2O1A1Ixp33_ASAP7_75t_R g215492 (.A1(n_1605),
    .A2(n_2464),
    .B(n_2074),
    .C(n_2962),
    .Y(n_4891));
 AO21x1_ASAP7_75t_R g215493 (.A1(n_2956),
    .A2(n_1547),
    .B(n_3923),
    .Y(n_4890));
 AO21x1_ASAP7_75t_L g215494 (.A1(n_2463),
    .A2(n_2414),
    .B(n_4607),
    .Y(n_4889));
 AOI22xp33_ASAP7_75t_L g215495 (.A1(n_3162),
    .A2(n_1641),
    .B1(n_2079),
    .B2(n_3413),
    .Y(n_4888));
 AOI22xp33_ASAP7_75t_L g215496 (.A1(n_3275),
    .A2(n_3164),
    .B1(n_3243),
    .B2(n_3047),
    .Y(n_4887));
 AOI21xp33_ASAP7_75t_R g215497 (.A1(n_2042),
    .A2(n_3414),
    .B(n_3941),
    .Y(n_4886));
 OAI21xp33_ASAP7_75t_R g215498 (.A1(n_2594),
    .A2(n_3261),
    .B(n_1664),
    .Y(n_4885));
 NAND3xp33_ASAP7_75t_R g215499 (.A(n_4314),
    .B(n_2823),
    .C(n_1447),
    .Y(n_4884));
 OAI21xp33_ASAP7_75t_R g215500 (.A1(n_2550),
    .A2(n_3259),
    .B(n_2421),
    .Y(n_4883));
 NAND3xp33_ASAP7_75t_L g215501 (.A(n_4434),
    .B(n_3358),
    .C(n_1411),
    .Y(n_4882));
 OAI21xp33_ASAP7_75t_R g215502 (.A1(n_2548),
    .A2(n_3252),
    .B(n_2427),
    .Y(n_4881));
 OAI21xp33_ASAP7_75t_L g215503 (.A1(n_2399),
    .A2(n_3167),
    .B(n_4522),
    .Y(n_4880));
 AO21x1_ASAP7_75t_R g215504 (.A1(n_2413),
    .A2(n_3127),
    .B(n_1591),
    .Y(n_4879));
 OAI21xp33_ASAP7_75t_R g215505 (.A1(n_2546),
    .A2(n_1729),
    .B(n_1349),
    .Y(n_4878));
 AOI22xp33_ASAP7_75t_L g215506 (.A1(n_1633),
    .A2(n_3033),
    .B1(n_2296),
    .B2(n_2040),
    .Y(n_4877));
 OAI22xp33_ASAP7_75t_R g215507 (.A1(n_1408),
    .A2(n_1756),
    .B1(n_2837),
    .B2(n_2056),
    .Y(n_4876));
 OA21x2_ASAP7_75t_SL g215508 (.A1(n_3046),
    .A2(n_2423),
    .B(n_2220),
    .Y(n_4875));
 OAI22xp5_ASAP7_75t_R g215509 (.A1(n_1567),
    .A2(n_2969),
    .B1(n_1565),
    .B2(n_3050),
    .Y(n_4874));
 OAI21xp5_ASAP7_75t_SL g215510 (.A1(n_2437),
    .A2(n_3713),
    .B(n_2394),
    .Y(n_4873));
 AOI21xp33_ASAP7_75t_R g215511 (.A1(n_3253),
    .A2(n_3341),
    .B(n_2428),
    .Y(n_4872));
 AOI32xp33_ASAP7_75t_R g215512 (.A1(n_2521),
    .A2(n_2439),
    .A3(n_1458),
    .B1(n_1422),
    .B2(n_2128),
    .Y(n_4871));
 AOI211xp5_ASAP7_75t_R g215513 (.A1(n_3275),
    .A2(n_2064),
    .B(n_3208),
    .C(n_3026),
    .Y(n_4870));
 AOI21xp33_ASAP7_75t_L g215514 (.A1(n_2386),
    .A2(n_1681),
    .B(n_4065),
    .Y(n_4869));
 OAI22xp5_ASAP7_75t_R g215515 (.A1(n_1656),
    .A2(n_2918),
    .B1(n_3023),
    .B2(n_1344),
    .Y(n_4868));
 OAI32xp33_ASAP7_75t_R g215516 (.A1(n_2580),
    .A2(n_2445),
    .A3(n_1496),
    .B1(n_1594),
    .B2(n_1556),
    .Y(n_4867));
 AO21x1_ASAP7_75t_L g215517 (.A1(n_2465),
    .A2(n_2435),
    .B(n_4053),
    .Y(n_4866));
 OA21x2_ASAP7_75t_L g215518 (.A1(n_2111),
    .A2(n_3012),
    .B(n_4155),
    .Y(n_4865));
 AO22x1_ASAP7_75t_R g215519 (.A1(n_2930),
    .A2(n_1405),
    .B1(n_2075),
    .B2(n_3034),
    .Y(n_4864));
 AOI32xp33_ASAP7_75t_R g215520 (.A1(n_2475),
    .A2(n_2523),
    .A3(n_1500),
    .B1(n_1350),
    .B2(n_2142),
    .Y(n_4863));
 OAI21xp33_ASAP7_75t_L g215521 (.A1(n_1673),
    .A2(n_1623),
    .B(n_4204),
    .Y(n_4862));
 OA21x2_ASAP7_75t_L g215522 (.A1(n_1683),
    .A2(n_1382),
    .B(n_4194),
    .Y(n_4861));
 OA21x2_ASAP7_75t_L g215523 (.A1(n_2471),
    .A2(n_1656),
    .B(n_4200),
    .Y(n_4860));
 NOR4xp25_ASAP7_75t_R g215524 (.A(n_4278),
    .B(n_1450),
    .C(n_8182),
    .D(n_2634),
    .Y(n_4859));
 AOI21xp5_ASAP7_75t_R g215525 (.A1(n_3698),
    .A2(n_1496),
    .B(n_4106),
    .Y(n_4858));
 AOI22xp33_ASAP7_75t_R g215526 (.A1(n_2413),
    .A2(n_2999),
    .B1(n_2195),
    .B2(n_2064),
    .Y(n_4857));
 NAND3xp33_ASAP7_75t_R g215527 (.A(n_2777),
    .B(n_2859),
    .C(n_2350),
    .Y(n_4856));
 OAI21xp33_ASAP7_75t_L g215528 (.A1(n_1680),
    .A2(n_1646),
    .B(n_4105),
    .Y(n_4855));
 OR3x1_ASAP7_75t_L g215529 (.A(n_2787),
    .B(n_3345),
    .C(n_1839),
    .Y(n_4854));
 OAI22xp33_ASAP7_75t_R g215530 (.A1(n_1626),
    .A2(n_3035),
    .B1(n_2270),
    .B2(n_2078),
    .Y(n_4853));
 AOI21xp33_ASAP7_75t_R g215531 (.A1(n_2815),
    .A2(n_2473),
    .B(n_1344),
    .Y(n_4852));
 AOI21xp33_ASAP7_75t_R g215532 (.A1(n_1595),
    .A2(n_1732),
    .B(n_2088),
    .Y(n_4851));
 AOI22xp33_ASAP7_75t_R g215533 (.A1(n_2401),
    .A2(n_2946),
    .B1(n_2274),
    .B2(n_1577),
    .Y(n_4850));
 AOI21xp33_ASAP7_75t_R g215534 (.A1(n_2897),
    .A2(n_1496),
    .B(n_2276),
    .Y(n_4849));
 AOI21xp33_ASAP7_75t_R g215535 (.A1(n_2892),
    .A2(n_1464),
    .B(n_2151),
    .Y(n_4848));
 OAI21xp33_ASAP7_75t_L g215536 (.A1(n_2170),
    .A2(n_2808),
    .B(n_1587),
    .Y(n_4847));
 OAI21xp33_ASAP7_75t_R g215537 (.A1(n_2504),
    .A2(n_3293),
    .B(n_1586),
    .Y(n_4846));
 AOI21xp33_ASAP7_75t_L g215538 (.A1(n_3147),
    .A2(n_1457),
    .B(n_4163),
    .Y(n_4845));
 AOI21xp5_ASAP7_75t_R g215539 (.A1(n_3275),
    .A2(n_2481),
    .B(n_1418),
    .Y(n_4844));
 OAI21xp33_ASAP7_75t_R g215540 (.A1(n_3272),
    .A2(n_2111),
    .B(n_1374),
    .Y(n_4843));
 OAI21xp33_ASAP7_75t_R g215541 (.A1(n_2120),
    .A2(n_2816),
    .B(n_2072),
    .Y(n_4842));
 OAI21xp33_ASAP7_75t_R g215542 (.A1(n_2803),
    .A2(n_1604),
    .B(n_2075),
    .Y(n_4841));
 OAI21xp33_ASAP7_75t_R g215543 (.A1(n_2815),
    .A2(n_2096),
    .B(n_1576),
    .Y(n_4840));
 NAND3xp33_ASAP7_75t_L g215544 (.A(n_1730),
    .B(n_1621),
    .C(n_1715),
    .Y(n_4839));
 NOR3xp33_ASAP7_75t_R g215545 (.A(n_2881),
    .B(n_1344),
    .C(n_3337),
    .Y(n_4838));
 AOI21xp33_ASAP7_75t_R g215546 (.A1(n_2917),
    .A2(n_2471),
    .B(n_3859),
    .Y(n_4837));
 OR3x1_ASAP7_75t_L g215547 (.A(n_2786),
    .B(n_2826),
    .C(n_2347),
    .Y(n_4836));
 OA21x2_ASAP7_75t_R g215548 (.A1(n_1337),
    .A2(n_3273),
    .B(n_3204),
    .Y(n_4835));
 OAI21xp5_ASAP7_75t_L g215549 (.A1(n_1336),
    .A2(n_3200),
    .B(n_4033),
    .Y(n_4834));
 NAND3xp33_ASAP7_75t_R g215550 (.A(n_3258),
    .B(n_2828),
    .C(n_2355),
    .Y(n_4833));
 NAND3xp33_ASAP7_75t_R g215551 (.A(n_3297),
    .B(n_2364),
    .C(n_3247),
    .Y(n_4832));
 NAND3xp33_ASAP7_75t_R g215552 (.A(n_3243),
    .B(n_3291),
    .C(n_2370),
    .Y(n_4831));
 AOI21xp33_ASAP7_75t_R g215553 (.A1(n_2192),
    .A2(n_1711),
    .B(n_1342),
    .Y(n_4830));
 AOI21xp33_ASAP7_75t_R g215554 (.A1(n_3246),
    .A2(n_2837),
    .B(n_1417),
    .Y(n_4829));
 AOI21xp5_ASAP7_75t_R g215555 (.A1(n_2808),
    .A2(n_1587),
    .B(n_3185),
    .Y(n_4828));
 AOI21xp33_ASAP7_75t_R g215556 (.A1(n_2792),
    .A2(n_1577),
    .B(n_2736),
    .Y(n_4827));
 AOI21xp5_ASAP7_75t_L g215557 (.A1(n_2784),
    .A2(n_2090),
    .B(n_3209),
    .Y(n_4826));
 OAI21xp33_ASAP7_75t_R g215558 (.A1(n_1573),
    .A2(n_1711),
    .B(n_3194),
    .Y(n_4825));
 A2O1A1Ixp33_ASAP7_75t_R g215559 (.A1(n_2439),
    .A2(n_2521),
    .B(n_2399),
    .C(n_2765),
    .Y(n_4824));
 OAI21xp33_ASAP7_75t_R g215560 (.A1(n_2850),
    .A2(n_2818),
    .B(n_2062),
    .Y(n_4823));
 OAI21xp5_ASAP7_75t_R g215561 (.A1(n_2830),
    .A2(n_2822),
    .B(n_2058),
    .Y(n_4822));
 O2A1O1Ixp33_ASAP7_75t_R g215562 (.A1(n_2465),
    .A2(n_2558),
    .B(n_1860),
    .C(n_4257),
    .Y(n_4821));
 AOI22xp5_ASAP7_75t_L g215563 (.A1(n_2753),
    .A2(n_1627),
    .B1(n_2252),
    .B2(n_2072),
    .Y(n_4820));
 AOI22xp33_ASAP7_75t_R g215564 (.A1(n_2749),
    .A2(n_2079),
    .B1(n_3179),
    .B2(n_1445),
    .Y(n_4819));
 AOI221xp5_ASAP7_75t_L g215565 (.A1(n_2940),
    .A2(n_2505),
    .B1(n_1552),
    .B2(n_2212),
    .C(n_3235),
    .Y(n_4818));
 OAI221xp5_ASAP7_75t_SL g215566 (.A1(n_3024),
    .A2(n_2501),
    .B1(n_1354),
    .B2(n_1610),
    .C(n_3232),
    .Y(n_4817));
 OAI22xp33_ASAP7_75t_R g215567 (.A1(n_1460),
    .A2(n_3628),
    .B1(n_1467),
    .B2(n_2879),
    .Y(n_4816));
 OAI21xp33_ASAP7_75t_SL g215568 (.A1(n_1498),
    .A2(n_2926),
    .B(n_3841),
    .Y(n_4815));
 AOI22xp33_ASAP7_75t_R g215569 (.A1(n_1455),
    .A2(n_3634),
    .B1(n_1512),
    .B2(n_3415),
    .Y(n_4814));
 OAI221xp5_ASAP7_75t_SL g215570 (.A1(n_2936),
    .A2(n_1395),
    .B1(n_2053),
    .B2(n_2140),
    .C(n_2764),
    .Y(n_4813));
 AOI22xp33_ASAP7_75t_R g215571 (.A1(n_3671),
    .A2(n_2389),
    .B1(n_1448),
    .B2(n_2584),
    .Y(n_4812));
 AOI22xp33_ASAP7_75t_SL g215572 (.A1(n_1416),
    .A2(n_3487),
    .B1(n_1483),
    .B2(n_2410),
    .Y(n_4811));
 AOI221xp5_ASAP7_75t_R g215573 (.A1(n_3084),
    .A2(n_2431),
    .B1(n_1448),
    .B2(n_2255),
    .C(n_3234),
    .Y(n_4810));
 OAI221xp5_ASAP7_75t_L g215574 (.A1(n_1582),
    .A2(n_2195),
    .B1(n_2196),
    .B2(n_1512),
    .C(n_3805),
    .Y(n_4809));
 OAI221xp5_ASAP7_75t_L g215575 (.A1(n_2047),
    .A2(n_2228),
    .B1(n_2229),
    .B2(sa03[3]),
    .C(n_3840),
    .Y(n_4808));
 AOI22xp33_ASAP7_75t_L g215576 (.A1(n_2398),
    .A2(n_3724),
    .B1(n_2567),
    .B2(n_1547),
    .Y(n_4807));
 AOI22xp33_ASAP7_75t_R g215577 (.A1(n_2390),
    .A2(n_3696),
    .B1(n_2222),
    .B2(n_1668),
    .Y(n_4806));
 OAI22xp33_ASAP7_75t_L g215578 (.A1(n_1660),
    .A2(n_3716),
    .B1(n_2561),
    .B2(n_1450),
    .Y(n_4805));
 AOI221xp5_ASAP7_75t_R g215579 (.A1(n_2497),
    .A2(n_1458),
    .B1(n_1423),
    .B2(n_8212),
    .C(n_8208),
    .Y(n_4804));
 AO22x1_ASAP7_75t_L g215580 (.A1(n_1641),
    .A2(n_3714),
    .B1(n_2555),
    .B2(n_2042),
    .Y(n_4803));
 OAI221xp5_ASAP7_75t_L g215581 (.A1(n_2056),
    .A2(n_1611),
    .B1(n_1612),
    .B2(sa00[3]),
    .C(n_3812),
    .Y(n_4802));
 OAI221xp5_ASAP7_75t_R g215582 (.A1(n_1548),
    .A2(n_2243),
    .B1(n_2242),
    .B2(n_1984),
    .C(n_3796),
    .Y(n_4801));
 OAI22xp33_ASAP7_75t_R g215583 (.A1(n_3711),
    .A2(n_2419),
    .B1(n_1417),
    .B2(n_2585),
    .Y(n_4800));
 AOI22xp33_ASAP7_75t_R g215584 (.A1(n_2431),
    .A2(n_2958),
    .B1(n_2256),
    .B2(n_1589),
    .Y(n_4799));
 OAI22xp33_ASAP7_75t_R g215585 (.A1(n_1536),
    .A2(n_2986),
    .B1(n_1602),
    .B2(n_2396),
    .Y(n_4798));
 AOI22xp33_ASAP7_75t_R g215586 (.A1(n_2089),
    .A2(n_2945),
    .B1(n_2306),
    .B2(n_2048),
    .Y(n_4797));
 AOI22xp33_ASAP7_75t_SL g215587 (.A1(n_2398),
    .A2(n_3160),
    .B1(n_2039),
    .B2(n_3586),
    .Y(n_4796));
 AOI221xp5_ASAP7_75t_SL g215588 (.A1(n_1444),
    .A2(n_2234),
    .B1(n_2235),
    .B2(n_8210),
    .C(n_4221),
    .Y(n_4795));
 AOI22xp33_ASAP7_75t_R g215589 (.A1(n_1467),
    .A2(n_2995),
    .B1(n_2055),
    .B2(n_2240),
    .Y(n_4794));
 OAI22xp33_ASAP7_75t_R g215590 (.A1(sa01[3]),
    .A2(n_3082),
    .B1(n_2057),
    .B2(n_2223),
    .Y(n_4793));
 OAI21xp33_ASAP7_75t_L g215591 (.A1(n_3395),
    .A2(n_3116),
    .B(n_4274),
    .Y(n_4792));
 AOI22xp33_ASAP7_75t_R g215592 (.A1(n_1986),
    .A2(n_3028),
    .B1(n_2044),
    .B2(n_2187),
    .Y(n_4791));
 OAI222xp33_ASAP7_75t_L g215593 (.A1(n_1562),
    .A2(n_2249),
    .B1(n_1568),
    .B2(n_3049),
    .C1(n_2248),
    .C2(n_1343),
    .Y(n_4790));
 OAI22xp33_ASAP7_75t_L g215594 (.A1(n_3731),
    .A2(n_2415),
    .B1(n_2127),
    .B2(n_1647),
    .Y(n_4789));
 AOI22xp33_ASAP7_75t_L g215595 (.A1(n_1566),
    .A2(n_3144),
    .B1(n_1561),
    .B2(n_1757),
    .Y(n_4788));
 AOI221xp5_ASAP7_75t_L g215596 (.A1(n_2231),
    .A2(n_1518),
    .B1(n_2421),
    .B2(n_3052),
    .C(n_2768),
    .Y(n_4787));
 AOI22xp33_ASAP7_75t_R g215597 (.A1(n_1653),
    .A2(n_3223),
    .B1(n_2240),
    .B2(n_2410),
    .Y(n_4786));
 AOI211xp5_ASAP7_75t_L g215598 (.A1(n_2940),
    .A2(n_3329),
    .B(n_3121),
    .C(n_3678),
    .Y(n_4785));
 AOI22xp5_ASAP7_75t_SL g215599 (.A1(n_2394),
    .A2(n_3101),
    .B1(n_1549),
    .B2(n_3599),
    .Y(n_4784));
 AOI22xp33_ASAP7_75t_L g215600 (.A1(n_8178),
    .A2(n_3588),
    .B1(n_1552),
    .B2(n_2099),
    .Y(n_4783));
 OAI211xp5_ASAP7_75t_R g215601 (.A1(n_3280),
    .A2(n_3024),
    .B(n_3113),
    .C(n_3687),
    .Y(n_4782));
 AOI211xp5_ASAP7_75t_L g215602 (.A1(n_3109),
    .A2(n_3287),
    .B(n_3128),
    .C(n_3660),
    .Y(n_4781));
 OAI22xp33_ASAP7_75t_L g215603 (.A1(n_2393),
    .A2(n_3709),
    .B1(n_2174),
    .B2(n_2423),
    .Y(n_4780));
 OAI221xp5_ASAP7_75t_L g215604 (.A1(n_2061),
    .A2(n_2274),
    .B1(n_2275),
    .B2(sa33[3]),
    .C(n_3794),
    .Y(n_4779));
 OAI22xp33_ASAP7_75t_R g215605 (.A1(n_2052),
    .A2(n_1757),
    .B1(n_2157),
    .B2(n_1567),
    .Y(n_4778));
 AOI22xp33_ASAP7_75t_L g215606 (.A1(n_1424),
    .A2(n_3730),
    .B1(n_2310),
    .B2(n_1440),
    .Y(n_4777));
 AO22x1_ASAP7_75t_L g215607 (.A1(n_1423),
    .A2(n_3062),
    .B1(n_2293),
    .B2(n_2067),
    .Y(n_4776));
 AOI22xp5_ASAP7_75t_R g215608 (.A1(n_2069),
    .A2(n_3028),
    .B1(n_2329),
    .B2(n_2044),
    .Y(n_4775));
 AOI22xp33_ASAP7_75t_R g215609 (.A1(n_3701),
    .A2(n_1350),
    .B1(n_2143),
    .B2(n_1446),
    .Y(n_4774));
 AOI22xp33_ASAP7_75t_L g215610 (.A1(sa03[3]),
    .A2(n_1731),
    .B1(n_1967),
    .B2(n_2945),
    .Y(n_4773));
 AOI211xp5_ASAP7_75t_R g215611 (.A1(n_3098),
    .A2(n_3334),
    .B(n_3637),
    .C(n_3037),
    .Y(n_4772));
 AOI211xp5_ASAP7_75t_R g215612 (.A1(n_2938),
    .A2(n_2900),
    .B(n_3635),
    .C(n_3010),
    .Y(n_4771));
 OAI22xp5_ASAP7_75t_L g215613 (.A1(n_2045),
    .A2(n_3581),
    .B1(n_2107),
    .B2(n_1662),
    .Y(n_4770));
 OAI22xp33_ASAP7_75t_R g215614 (.A1(n_1573),
    .A2(n_2996),
    .B1(n_2316),
    .B2(n_2056),
    .Y(n_4769));
 OAI22xp33_ASAP7_75t_R g215615 (.A1(n_1749),
    .A2(n_1565),
    .B1(n_2619),
    .B2(n_1560),
    .Y(n_4768));
 AOI22xp33_ASAP7_75t_R g215616 (.A1(n_3079),
    .A2(sa33[3]),
    .B1(n_2416),
    .B2(n_8189),
    .Y(n_4767));
 OAI32xp33_ASAP7_75t_R g215617 (.A1(n_2424),
    .A2(n_2786),
    .A3(n_2313),
    .B1(n_2011),
    .B2(n_2073),
    .Y(n_4766));
 OAI211xp5_ASAP7_75t_R g215618 (.A1(n_2256),
    .A2(n_1637),
    .B(n_2823),
    .C(sa01[0]),
    .Y(n_4765));
 OAI22xp33_ASAP7_75t_L g215619 (.A1(n_1624),
    .A2(n_3367),
    .B1(n_1639),
    .B2(n_1719),
    .Y(n_4764));
 AOI211xp5_ASAP7_75t_L g215620 (.A1(n_1445),
    .A2(n_2271),
    .B(n_2821),
    .C(n_1870),
    .Y(n_4763));
 OAI22xp33_ASAP7_75t_L g215621 (.A1(n_1568),
    .A2(n_3499),
    .B1(n_1565),
    .B2(n_2545),
    .Y(n_4762));
 AOI211xp5_ASAP7_75t_R g215622 (.A1(n_2398),
    .A2(n_2242),
    .B(n_2856),
    .C(n_8213),
    .Y(n_4761));
 OAI22xp33_ASAP7_75t_R g215623 (.A1(n_2434),
    .A2(n_3501),
    .B1(n_2557),
    .B2(n_2399),
    .Y(n_4760));
 OAI32xp33_ASAP7_75t_L g215624 (.A1(n_2173),
    .A2(n_1397),
    .A3(n_1525),
    .B1(n_8181),
    .B2(n_2904),
    .Y(n_4759));
 AOI22xp33_ASAP7_75t_R g215625 (.A1(n_2413),
    .A2(n_3511),
    .B1(n_2544),
    .B2(n_8703),
    .Y(n_4758));
 OAI22xp5_ASAP7_75t_L g215626 (.A1(n_1656),
    .A2(n_3495),
    .B1(n_2592),
    .B2(n_1662),
    .Y(n_4757));
 AOI22xp33_ASAP7_75t_R g215627 (.A1(n_3492),
    .A2(n_2420),
    .B1(n_2550),
    .B2(n_2392),
    .Y(n_4756));
 AOI22xp33_ASAP7_75t_R g215628 (.A1(n_2065),
    .A2(n_2941),
    .B1(n_1554),
    .B2(n_2580),
    .Y(n_4755));
 AOI22xp33_ASAP7_75t_R g215629 (.A1(n_3083),
    .A2(n_1589),
    .B1(n_2332),
    .B2(n_1448),
    .Y(n_4754));
 AOI22xp33_ASAP7_75t_SL g215630 (.A1(n_1636),
    .A2(n_1722),
    .B1(n_2560),
    .B2(n_1645),
    .Y(n_4753));
 AOI211xp5_ASAP7_75t_R g215631 (.A1(n_2229),
    .A2(n_2046),
    .B(n_2797),
    .C(n_1509),
    .Y(n_4752));
 AOI22xp33_ASAP7_75t_R g215632 (.A1(n_1622),
    .A2(n_2934),
    .B1(n_2552),
    .B2(n_1445),
    .Y(n_4751));
 OAI321xp33_ASAP7_75t_R g215633 (.A1(n_2131),
    .A2(n_1496),
    .A3(n_1534),
    .B1(n_1967),
    .B2(n_2891),
    .C(n_1553),
    .Y(n_4750));
 AOI22xp5_ASAP7_75t_R g215634 (.A1(n_2893),
    .A2(n_2390),
    .B1(n_2606),
    .B2(n_2058),
    .Y(n_4749));
 AOI21xp5_ASAP7_75t_R g215635 (.A1(n_3420),
    .A2(n_1343),
    .B(n_2773),
    .Y(n_4748));
 OAI22xp33_ASAP7_75t_R g215636 (.A1(n_2541),
    .A2(n_3379),
    .B1(n_2238),
    .B2(n_2844),
    .Y(n_4747));
 OAI221xp5_ASAP7_75t_R g215637 (.A1(n_3241),
    .A2(n_2083),
    .B1(n_1548),
    .B2(n_1852),
    .C(n_2627),
    .Y(n_4746));
 AOI22xp33_ASAP7_75t_L g215638 (.A1(n_1622),
    .A2(n_2943),
    .B1(n_1475),
    .B2(n_1435),
    .Y(n_4745));
 AOI32xp33_ASAP7_75t_R g215639 (.A1(n_2604),
    .A2(n_1687),
    .A3(sa23[3]),
    .B1(n_3305),
    .B2(n_1983),
    .Y(n_4744));
 AOI32xp33_ASAP7_75t_SL g215640 (.A1(n_2048),
    .A2(n_1595),
    .A3(n_2020),
    .B1(n_1366),
    .B2(n_2228),
    .Y(n_4743));
 OAI22xp5_ASAP7_75t_R g215641 (.A1(n_3029),
    .A2(n_1647),
    .B1(n_1580),
    .B2(n_3030),
    .Y(n_4742));
 AO22x1_ASAP7_75t_R g215642 (.A1(sa20[3]),
    .A2(n_3124),
    .B1(n_1867),
    .B2(n_3294),
    .Y(n_4741));
 AOI32xp33_ASAP7_75t_R g215643 (.A1(n_1683),
    .A2(n_2547),
    .A3(sa22[3]),
    .B1(n_3279),
    .B2(n_1985),
    .Y(n_4740));
 AOI32xp33_ASAP7_75t_L g215644 (.A1(n_2044),
    .A2(n_2095),
    .A3(n_1480),
    .B1(n_1576),
    .B2(n_2227),
    .Y(n_4739));
 AOI32xp33_ASAP7_75t_R g215645 (.A1(n_2559),
    .A2(n_1682),
    .A3(n_1984),
    .B1(n_3307),
    .B2(n_8181),
    .Y(n_4738));
 AOI221xp5_ASAP7_75t_L g215646 (.A1(n_2817),
    .A2(n_1356),
    .B1(n_1545),
    .B2(n_1503),
    .C(n_2631),
    .Y(n_4737));
 AOI22xp33_ASAP7_75t_SL g215647 (.A1(n_1625),
    .A2(n_2991),
    .B1(n_3175),
    .B2(n_2079),
    .Y(n_4736));
 OAI22xp33_ASAP7_75t_R g215648 (.A1(n_3570),
    .A2(n_1967),
    .B1(n_1556),
    .B2(n_1425),
    .Y(n_4735));
 AOI32xp33_ASAP7_75t_L g215649 (.A1(n_2055),
    .A2(n_2192),
    .A3(n_1477),
    .B1(n_2965),
    .B2(n_2410),
    .Y(n_4734));
 AOI221xp5_ASAP7_75t_R g215650 (.A1(n_2054),
    .A2(sa22[4]),
    .B1(n_2782),
    .B2(n_2082),
    .C(n_2204),
    .Y(n_4733));
 AOI32xp33_ASAP7_75t_L g215651 (.A1(n_1677),
    .A2(n_2574),
    .A3(sa21[3]),
    .B1(n_2834),
    .B2(n_1975),
    .Y(n_4732));
 AOI221xp5_ASAP7_75t_L g215652 (.A1(n_1435),
    .A2(n_1375),
    .B1(n_2789),
    .B2(n_1391),
    .C(n_2188),
    .Y(n_4731));
 OAI22xp33_ASAP7_75t_R g215653 (.A1(n_1669),
    .A2(n_2912),
    .B1(n_2564),
    .B2(n_1637),
    .Y(n_4730));
 OAI32xp33_ASAP7_75t_R g215654 (.A1(n_8178),
    .A2(n_2594),
    .A3(n_2487),
    .B1(n_3289),
    .B2(n_1972),
    .Y(n_4729));
 AOI22xp5_ASAP7_75t_L g215655 (.A1(n_1343),
    .A2(n_3542),
    .B1(n_8894),
    .B2(n_2051),
    .Y(n_4728));
 AOI32xp33_ASAP7_75t_R g215656 (.A1(n_2564),
    .A2(n_1670),
    .A3(sa01[3]),
    .B1(n_2825),
    .B2(n_1859),
    .Y(n_4727));
 AOI22xp33_ASAP7_75t_R g215657 (.A1(n_1860),
    .A2(n_3562),
    .B1(n_8212),
    .B2(n_1421),
    .Y(n_4726));
 AO32x1_ASAP7_75t_R g215658 (.A1(n_1559),
    .A2(n_2205),
    .A3(n_1992),
    .B1(n_2090),
    .B2(n_2249),
    .Y(n_4725));
 AOI22xp33_ASAP7_75t_R g215659 (.A1(n_3566),
    .A2(n_1519),
    .B1(n_2392),
    .B2(n_1505),
    .Y(n_4724));
 OAI22xp33_ASAP7_75t_R g215660 (.A1(n_3536),
    .A2(n_1467),
    .B1(n_2419),
    .B2(n_1853),
    .Y(n_4723));
 OAI32xp33_ASAP7_75t_L g215661 (.A1(n_2546),
    .A2(n_2495),
    .A3(n_1507),
    .B1(n_1343),
    .B2(n_2845),
    .Y(n_4722));
 AOI221xp5_ASAP7_75t_R g215662 (.A1(n_1559),
    .A2(n_8899),
    .B1(n_2783),
    .B2(n_1412),
    .C(n_2250),
    .Y(n_4721));
 OAI32xp33_ASAP7_75t_R g215663 (.A1(n_2580),
    .A2(n_2445),
    .A3(n_1967),
    .B1(sa03[3]),
    .B2(n_3314),
    .Y(n_4720));
 AOI22xp33_ASAP7_75t_R g215664 (.A1(n_1497),
    .A2(n_2960),
    .B1(n_2130),
    .B2(n_1554),
    .Y(n_4719));
 AOI221xp5_ASAP7_75t_R g215665 (.A1(n_1419),
    .A2(n_1851),
    .B1(n_1577),
    .B2(n_2793),
    .C(n_2164),
    .Y(n_4718));
 AOI22xp33_ASAP7_75t_R g215666 (.A1(n_2087),
    .A2(n_2811),
    .B1(n_1385),
    .B2(n_1448),
    .Y(n_4717));
 AOI22xp33_ASAP7_75t_R g215667 (.A1(n_1366),
    .A2(n_1732),
    .B1(n_1425),
    .B2(n_1438),
    .Y(n_4716));
 AOI22xp33_ASAP7_75t_R g215668 (.A1(sa30[6]),
    .A2(n_3053),
    .B1(n_2169),
    .B2(n_1641),
    .Y(n_4715));
 AOI22xp33_ASAP7_75t_R g215669 (.A1(n_1934),
    .A2(n_3052),
    .B1(n_2174),
    .B2(n_2392),
    .Y(n_4714));
 OAI22xp33_ASAP7_75t_R g215670 (.A1(n_3049),
    .A2(n_1499),
    .B1(n_2052),
    .B2(n_2158),
    .Y(n_4713));
 AOI22xp33_ASAP7_75t_R g215671 (.A1(n_1455),
    .A2(n_3063),
    .B1(n_1609),
    .B2(n_8703),
    .Y(n_4712));
 OAI22xp33_ASAP7_75t_R g215672 (.A1(n_2395),
    .A2(n_3372),
    .B1(n_2645),
    .B2(n_2041),
    .Y(n_4711));
 AOI22xp33_ASAP7_75t_L g215673 (.A1(n_1377),
    .A2(n_2734),
    .B1(n_2095),
    .B2(n_1659),
    .Y(n_4710));
 OAI22xp5_ASAP7_75t_L g215674 (.A1(n_1651),
    .A2(n_3496),
    .B1(n_3555),
    .B2(n_2063),
    .Y(n_4709));
 OAI22xp33_ASAP7_75t_R g215675 (.A1(n_2961),
    .A2(n_3372),
    .B1(n_3273),
    .B2(n_2041),
    .Y(n_4708));
 AOI22xp5_ASAP7_75t_L g215676 (.A1(n_1507),
    .A2(n_3386),
    .B1(n_1343),
    .B2(n_3425),
    .Y(n_5108));
 AOI22xp5_ASAP7_75t_L g215677 (.A1(n_8178),
    .A2(n_3322),
    .B1(n_1972),
    .B2(n_3450),
    .Y(n_5107));
 OAI22xp5_ASAP7_75t_R g215678 (.A1(sa22[3]),
    .A2(n_3370),
    .B1(n_1985),
    .B2(n_3423),
    .Y(n_5106));
 AOI22xp5_ASAP7_75t_R g215679 (.A1(n_8177),
    .A2(n_3368),
    .B1(sa30[3]),
    .B2(n_3414),
    .Y(n_5105));
 OAI22xp33_ASAP7_75t_R g215680 (.A1(sa33[3]),
    .A2(n_3357),
    .B1(n_1979),
    .B2(n_3546),
    .Y(n_5104));
 AO22x1_ASAP7_75t_L g215681 (.A1(n_1975),
    .A2(n_3356),
    .B1(sa21[3]),
    .B2(n_3519),
    .Y(n_5103));
 AOI22xp5_ASAP7_75t_R g215682 (.A1(n_8181),
    .A2(n_3347),
    .B1(n_1984),
    .B2(n_3516),
    .Y(n_5101));
 AOI22xp33_ASAP7_75t_L g215683 (.A1(n_1867),
    .A2(n_3348),
    .B1(sa20[3]),
    .B2(n_3453),
    .Y(n_5100));
 OAI22xp5_ASAP7_75t_R g215684 (.A1(sa23[3]),
    .A2(n_3355),
    .B1(n_1983),
    .B2(n_3455),
    .Y(n_5099));
 OAI22xp5_ASAP7_75t_L g215685 (.A1(n_1986),
    .A2(n_3560),
    .B1(sa11[3]),
    .B2(n_3337),
    .Y(n_5098));
 OAI22xp5_ASAP7_75t_L g215686 (.A1(n_8210),
    .A2(n_2887),
    .B1(n_1860),
    .B2(n_3319),
    .Y(n_1789));
 AOI22xp5_ASAP7_75t_R g215687 (.A1(n_1519),
    .A2(n_1752),
    .B1(n_1518),
    .B2(n_3332),
    .Y(n_5097));
 AOI22xp5_ASAP7_75t_R g215688 (.A1(sa00[3]),
    .A2(n_3592),
    .B1(n_1467),
    .B2(n_1743),
    .Y(n_5096));
 AOI21xp5_ASAP7_75t_R g215689 (.A1(n_3297),
    .A2(n_2496),
    .B(n_2074),
    .Y(n_5095));
 OAI21xp5_ASAP7_75t_R g215690 (.A1(n_2504),
    .A2(n_2829),
    .B(n_1586),
    .Y(n_5093));
 NAND2xp33_ASAP7_75t_R g215691 (.A(n_2064),
    .B(n_4706),
    .Y(n_4707));
 OAI21xp5_ASAP7_75t_R g215692 (.A1(n_2507),
    .A2(n_2838),
    .B(n_1570),
    .Y(n_5091));
 OAI21xp5_ASAP7_75t_R g215693 (.A1(n_2520),
    .A2(n_2844),
    .B(n_1576),
    .Y(n_5089));
 AOI21xp33_ASAP7_75t_R g215694 (.A1(n_2534),
    .A2(n_3361),
    .B(n_2081),
    .Y(n_5088));
 OAI21xp5_ASAP7_75t_L g215695 (.A1(n_2511),
    .A2(n_2848),
    .B(n_2089),
    .Y(n_5087));
 AOI22xp33_ASAP7_75t_R g215696 (.A1(sa01[3]),
    .A2(n_3449),
    .B1(n_1859),
    .B2(n_3317),
    .Y(n_5086));
 AOI21xp33_ASAP7_75t_R g215697 (.A1(n_2525),
    .A2(n_3312),
    .B(n_1337),
    .Y(n_5085));
 AOI21xp33_ASAP7_75t_R g215698 (.A1(n_1715),
    .A2(n_2537),
    .B(n_2091),
    .Y(n_5084));
 OAI21xp5_ASAP7_75t_L g215699 (.A1(n_2532),
    .A2(n_2858),
    .B(n_2084),
    .Y(n_5083));
 AOI21xp33_ASAP7_75t_R g215700 (.A1(n_2831),
    .A2(n_1691),
    .B(n_1588),
    .Y(n_5082));
 NOR3xp33_ASAP7_75t_L g215701 (.A(n_2911),
    .B(n_2825),
    .C(n_2057),
    .Y(n_5080));
 OAI21xp5_ASAP7_75t_R g215702 (.A1(n_2572),
    .A2(n_2850),
    .B(n_1577),
    .Y(n_5078));
 NAND3xp33_ASAP7_75t_R g215703 (.A(n_3278),
    .B(n_2054),
    .C(n_3447),
    .Y(n_5077));
 OAI21xp5_ASAP7_75t_R g215704 (.A1(n_2825),
    .A2(n_2911),
    .B(n_1667),
    .Y(n_5076));
 AOI22xp5_ASAP7_75t_R g215705 (.A1(n_1512),
    .A2(n_3533),
    .B1(n_1971),
    .B2(n_3325),
    .Y(n_5075));
 OAI21xp5_ASAP7_75t_L g215706 (.A1(n_3279),
    .A2(n_3446),
    .B(n_2427),
    .Y(n_5073));
 NAND3xp33_ASAP7_75t_SL g215707 (.A(n_4291),
    .B(n_3262),
    .C(n_2414),
    .Y(n_5072));
 OAI21xp5_ASAP7_75t_R g215708 (.A1(n_8200),
    .A2(n_1710),
    .B(n_2192),
    .Y(n_5070));
 NAND2xp5_ASAP7_75t_L g215709 (.A(n_2759),
    .B(n_4343),
    .Y(n_5069));
 AOI21xp5_ASAP7_75t_R g215710 (.A1(n_2817),
    .A2(n_1503),
    .B(n_2120),
    .Y(n_5068));
 AO21x1_ASAP7_75t_SL g215711 (.A1(n_1375),
    .A2(n_2789),
    .B(n_2214),
    .Y(n_5066));
 OAI22xp33_ASAP7_75t_R g215712 (.A1(n_1967),
    .A2(n_3482),
    .B1(sa03[3]),
    .B2(n_3374),
    .Y(n_5065));
 NOR2xp33_ASAP7_75t_L g215713 (.A(n_2758),
    .B(n_4337),
    .Y(n_5064));
 AOI21xp5_ASAP7_75t_L g215714 (.A1(n_1385),
    .A2(n_2809),
    .B(n_2170),
    .Y(n_5063));
 OAI21xp33_ASAP7_75t_R g215715 (.A1(n_1852),
    .A2(n_3241),
    .B(n_2103),
    .Y(n_5061));
 AOI21xp5_ASAP7_75t_R g215716 (.A1(n_8899),
    .A2(n_2783),
    .B(n_2206),
    .Y(n_1788));
 OAI21xp33_ASAP7_75t_R g215717 (.A1(n_1950),
    .A2(n_3271),
    .B(n_1606),
    .Y(n_5059));
 OAI21xp5_ASAP7_75t_R g215718 (.A1(n_8212),
    .A2(n_2803),
    .B(n_1605),
    .Y(n_5057));
 AO21x1_ASAP7_75t_L g215719 (.A1(sa22[4]),
    .A2(n_2782),
    .B(n_1602),
    .Y(n_5055));
 AOI21xp33_ASAP7_75t_R g215720 (.A1(sa23[4]),
    .A2(n_3266),
    .B(n_2160),
    .Y(n_5053));
 NOR2xp33_ASAP7_75t_L g215721 (.A(n_2760),
    .B(n_4356),
    .Y(n_5051));
 OAI21xp5_ASAP7_75t_L g215722 (.A1(n_1505),
    .A2(n_1726),
    .B(n_2178),
    .Y(n_5049));
 OAI21xp5_ASAP7_75t_SL g215723 (.A1(n_3372),
    .A2(n_2437),
    .B(n_1972),
    .Y(n_5048));
 INVxp67_ASAP7_75t_R g215724 (.A(n_4701),
    .Y(n_4702));
 INVxp33_ASAP7_75t_R g215725 (.A(n_4697),
    .Y(n_4698));
 INVxp67_ASAP7_75t_R g215726 (.A(n_4694),
    .Y(n_4695));
 INVxp33_ASAP7_75t_R g215727 (.A(n_4692),
    .Y(n_4693));
 INVxp33_ASAP7_75t_R g215728 (.A(n_4685),
    .Y(n_4686));
 INVxp67_ASAP7_75t_R g215729 (.A(n_4683),
    .Y(n_4684));
 INVxp33_ASAP7_75t_R g215730 (.A(n_4676),
    .Y(n_4677));
 INVxp33_ASAP7_75t_R g215731 (.A(n_4674),
    .Y(n_4675));
 INVxp33_ASAP7_75t_R g215732 (.A(n_4670),
    .Y(n_4671));
 INVxp67_ASAP7_75t_R g215733 (.A(n_4657),
    .Y(n_4658));
 INVxp33_ASAP7_75t_R g215734 (.A(n_4655),
    .Y(n_4656));
 INVxp67_ASAP7_75t_R g215735 (.A(n_4652),
    .Y(n_4653));
 INVxp67_ASAP7_75t_L g215737 (.A(n_4648),
    .Y(n_4649));
 INVxp33_ASAP7_75t_R g215738 (.A(n_4645),
    .Y(n_4646));
 INVxp67_ASAP7_75t_R g215739 (.A(n_4643),
    .Y(n_4644));
 INVxp33_ASAP7_75t_R g215740 (.A(n_4633),
    .Y(n_4634));
 INVxp67_ASAP7_75t_L g215741 (.A(n_4631),
    .Y(n_4632));
 INVxp67_ASAP7_75t_R g215742 (.A(n_4629),
    .Y(n_4630));
 INVxp33_ASAP7_75t_R g215743 (.A(n_4625),
    .Y(n_4626));
 INVxp67_ASAP7_75t_R g215744 (.A(n_4623),
    .Y(n_4624));
 INVx1_ASAP7_75t_R g215746 (.A(n_1340),
    .Y(n_4620));
 INVxp33_ASAP7_75t_R g215747 (.A(n_4618),
    .Y(n_4619));
 INVxp67_ASAP7_75t_R g215748 (.A(n_4615),
    .Y(n_4616));
 INVxp67_ASAP7_75t_R g215749 (.A(n_4613),
    .Y(n_4614));
 INVxp67_ASAP7_75t_L g215750 (.A(n_4604),
    .Y(n_4605));
 INVxp33_ASAP7_75t_R g215751 (.A(n_4598),
    .Y(n_4599));
 INVxp33_ASAP7_75t_R g215752 (.A(n_4596),
    .Y(n_4597));
 INVx1_ASAP7_75t_R g215753 (.A(n_4594),
    .Y(n_4595));
 INVxp67_ASAP7_75t_R g215754 (.A(n_4590),
    .Y(n_4591));
 INVxp33_ASAP7_75t_R g215755 (.A(n_4587),
    .Y(n_4588));
 INVxp67_ASAP7_75t_R g215756 (.A(n_4585),
    .Y(n_4586));
 INVxp67_ASAP7_75t_R g215757 (.A(n_4583),
    .Y(n_4584));
 INVxp67_ASAP7_75t_L g215758 (.A(n_4579),
    .Y(n_4580));
 INVxp33_ASAP7_75t_R g215759 (.A(n_4577),
    .Y(n_4578));
 INVxp67_ASAP7_75t_R g215761 (.A(n_4572),
    .Y(n_4573));
 INVxp67_ASAP7_75t_R g215762 (.A(n_4567),
    .Y(n_4568));
 INVxp33_ASAP7_75t_R g215763 (.A(n_4564),
    .Y(n_4565));
 INVxp67_ASAP7_75t_R g215764 (.A(n_4561),
    .Y(n_4562));
 INVxp33_ASAP7_75t_R g215765 (.A(n_4558),
    .Y(n_4559));
 INVxp33_ASAP7_75t_R g215766 (.A(n_4550),
    .Y(n_4551));
 INVxp33_ASAP7_75t_R g215767 (.A(n_4547),
    .Y(n_4548));
 INVxp67_ASAP7_75t_R g215768 (.A(n_4543),
    .Y(n_4544));
 INVxp67_ASAP7_75t_L g215769 (.A(n_4540),
    .Y(n_4541));
 INVxp67_ASAP7_75t_L g215770 (.A(n_4534),
    .Y(n_4535));
 INVxp33_ASAP7_75t_R g215771 (.A(n_4527),
    .Y(n_4528));
 INVxp33_ASAP7_75t_R g215772 (.A(n_4517),
    .Y(n_4518));
 INVxp67_ASAP7_75t_R g215773 (.A(n_4514),
    .Y(n_4515));
 INVx1_ASAP7_75t_L g215774 (.A(n_4513),
    .Y(n_4512));
 INVx1_ASAP7_75t_L g215775 (.A(n_4510),
    .Y(n_4511));
 INVxp67_ASAP7_75t_L g215776 (.A(n_4506),
    .Y(n_4507));
 INVxp33_ASAP7_75t_R g215777 (.A(n_4504),
    .Y(n_4505));
 INVxp33_ASAP7_75t_R g215778 (.A(n_4503),
    .Y(n_4502));
 INVxp67_ASAP7_75t_R g215779 (.A(n_4499),
    .Y(n_4500));
 INVxp67_ASAP7_75t_R g215780 (.A(n_4489),
    .Y(n_4490));
 INVxp67_ASAP7_75t_R g215781 (.A(n_4485),
    .Y(n_4486));
 INVxp67_ASAP7_75t_L g215782 (.A(n_4481),
    .Y(n_4480));
 INVxp33_ASAP7_75t_R g215784 (.A(n_4478),
    .Y(n_4479));
 INVxp67_ASAP7_75t_L g215785 (.A(n_4476),
    .Y(n_4477));
 INVxp33_ASAP7_75t_R g215786 (.A(n_4473),
    .Y(n_4474));
 INVxp67_ASAP7_75t_L g215788 (.A(n_4470),
    .Y(n_4471));
 INVxp33_ASAP7_75t_R g215789 (.A(n_4468),
    .Y(n_4469));
 INVxp67_ASAP7_75t_R g215792 (.A(n_4464),
    .Y(n_4465));
 INVxp67_ASAP7_75t_R g215793 (.A(n_4461),
    .Y(n_4462));
 INVx1_ASAP7_75t_L g215794 (.A(n_4459),
    .Y(n_4460));
 INVxp67_ASAP7_75t_R g215795 (.A(n_4458),
    .Y(n_4457));
 INVxp67_ASAP7_75t_L g215796 (.A(n_4455),
    .Y(n_4456));
 INVxp67_ASAP7_75t_R g215797 (.A(n_4453),
    .Y(n_4454));
 INVxp33_ASAP7_75t_R g215798 (.A(n_4451),
    .Y(n_4452));
 INVxp33_ASAP7_75t_R g215799 (.A(n_4445),
    .Y(n_4446));
 INVxp33_ASAP7_75t_R g215800 (.A(n_4443),
    .Y(n_4444));
 INVxp33_ASAP7_75t_R g215801 (.A(n_4441),
    .Y(n_4442));
 INVxp67_ASAP7_75t_L g215803 (.A(n_1782),
    .Y(n_4440));
 INVxp67_ASAP7_75t_R g215804 (.A(n_4437),
    .Y(n_4438));
 INVxp67_ASAP7_75t_R g215805 (.A(n_4436),
    .Y(n_4435));
 INVxp67_ASAP7_75t_R g215806 (.A(n_4432),
    .Y(n_4433));
 INVxp67_ASAP7_75t_R g215807 (.A(n_4430),
    .Y(n_4431));
 INVxp33_ASAP7_75t_R g215808 (.A(n_4425),
    .Y(n_4427));
 INVx1_ASAP7_75t_L g215810 (.A(n_4420),
    .Y(n_4421));
 INVxp33_ASAP7_75t_R g215811 (.A(n_4419),
    .Y(n_4418));
 INVxp67_ASAP7_75t_R g215812 (.A(n_4413),
    .Y(n_4414));
 INVxp67_ASAP7_75t_R g215813 (.A(n_4411),
    .Y(n_4412));
 INVxp67_ASAP7_75t_R g215814 (.A(n_4405),
    .Y(n_4406));
 INVxp67_ASAP7_75t_L g215815 (.A(n_4400),
    .Y(n_4401));
 INVxp33_ASAP7_75t_R g215816 (.A(n_4398),
    .Y(n_4397));
 INVxp33_ASAP7_75t_R g215817 (.A(n_4394),
    .Y(n_4395));
 INVxp67_ASAP7_75t_R g215818 (.A(n_4390),
    .Y(n_4389));
 INVxp67_ASAP7_75t_R g215819 (.A(n_4387),
    .Y(n_4388));
 INVxp33_ASAP7_75t_R g215820 (.A(n_4385),
    .Y(n_4386));
 INVxp67_ASAP7_75t_R g215821 (.A(n_4383),
    .Y(n_4384));
 INVxp33_ASAP7_75t_R g215823 (.A(n_4376),
    .Y(n_4377));
 INVxp67_ASAP7_75t_R g215824 (.A(n_4375),
    .Y(n_4374));
 INVxp33_ASAP7_75t_R g215825 (.A(n_4371),
    .Y(n_4372));
 INVxp67_ASAP7_75t_R g215826 (.A(n_4369),
    .Y(n_4370));
 INVxp67_ASAP7_75t_SL g215828 (.A(n_4368),
    .Y(n_4367));
 INVx1_ASAP7_75t_L g215829 (.A(n_4366),
    .Y(n_4365));
 INVx1_ASAP7_75t_R g215830 (.A(n_4364),
    .Y(n_4363));
 INVx1_ASAP7_75t_L g215831 (.A(n_4362),
    .Y(n_4361));
 INVxp67_ASAP7_75t_L g215832 (.A(n_4359),
    .Y(n_4358));
 INVxp33_ASAP7_75t_R g215833 (.A(n_4356),
    .Y(n_4357));
 INVxp67_ASAP7_75t_L g215834 (.A(n_4354),
    .Y(n_4353));
 INVx1_ASAP7_75t_L g215835 (.A(n_4352),
    .Y(n_4351));
 INVx1_ASAP7_75t_L g215836 (.A(n_4350),
    .Y(n_4349));
 INVx1_ASAP7_75t_R g215837 (.A(n_4347),
    .Y(n_4346));
 INVxp67_ASAP7_75t_L g215838 (.A(n_4343),
    .Y(n_4344));
 INVxp67_ASAP7_75t_L g215840 (.A(n_1780),
    .Y(n_4342));
 INVxp67_ASAP7_75t_R g215841 (.A(n_4340),
    .Y(n_4341));
 INVx1_ASAP7_75t_L g215842 (.A(n_4339),
    .Y(n_4340));
 INVx1_ASAP7_75t_SL g215843 (.A(n_4338),
    .Y(n_4337));
 INVx1_ASAP7_75t_R g215844 (.A(n_4336),
    .Y(n_4335));
 INVx1_ASAP7_75t_L g215846 (.A(n_4334),
    .Y(n_1779));
 INVx1_ASAP7_75t_L g215847 (.A(n_4333),
    .Y(n_4334));
 INVxp67_ASAP7_75t_R g215848 (.A(n_4332),
    .Y(n_4331));
 INVx1_ASAP7_75t_L g215852 (.A(n_1777),
    .Y(n_1778));
 INVxp67_ASAP7_75t_R g215853 (.A(n_4330),
    .Y(n_4329));
 INVx1_ASAP7_75t_L g215854 (.A(n_4328),
    .Y(n_4327));
 INVx2_ASAP7_75t_L g215855 (.A(n_4326),
    .Y(n_4325));
 INVx1_ASAP7_75t_R g215858 (.A(n_4324),
    .Y(n_1776));
 INVx2_ASAP7_75t_L g215859 (.A(n_4323),
    .Y(n_4322));
 INVxp67_ASAP7_75t_R g215860 (.A(n_4318),
    .Y(n_4321));
 INVx1_ASAP7_75t_L g215861 (.A(n_4319),
    .Y(n_4320));
 BUFx3_ASAP7_75t_SL g215863 (.A(n_4318),
    .Y(n_4319));
 INVx1_ASAP7_75t_L g215864 (.A(n_4317),
    .Y(n_4316));
 INVxp67_ASAP7_75t_L g215865 (.A(n_4315),
    .Y(n_4314));
 INVx1_ASAP7_75t_L g215866 (.A(n_4313),
    .Y(n_4312));
 INVx1_ASAP7_75t_R g215868 (.A(n_4310),
    .Y(n_4311));
 INVx1_ASAP7_75t_L g215869 (.A(n_1775),
    .Y(n_4310));
 INVxp33_ASAP7_75t_R g215870 (.A(n_4309),
    .Y(n_4308));
 INVx1_ASAP7_75t_L g215872 (.A(n_4307),
    .Y(n_4306));
 INVxp67_ASAP7_75t_R g215873 (.A(n_4305),
    .Y(n_4304));
 INVx2_ASAP7_75t_L g215874 (.A(n_4302),
    .Y(n_4301));
 INVx1_ASAP7_75t_SL g215875 (.A(n_4300),
    .Y(n_4299));
 INVx2_ASAP7_75t_SL g215876 (.A(n_4298),
    .Y(n_4297));
 INVx2_ASAP7_75t_L g215877 (.A(n_4296),
    .Y(n_4295));
 INVxp67_ASAP7_75t_R g215878 (.A(n_4294),
    .Y(n_4293));
 INVx1_ASAP7_75t_L g215879 (.A(n_4292),
    .Y(n_4291));
 INVx1_ASAP7_75t_SL g215881 (.A(n_4290),
    .Y(n_4289));
 INVx2_ASAP7_75t_L g215882 (.A(n_4288),
    .Y(n_4287));
 INVx1_ASAP7_75t_L g215883 (.A(n_4286),
    .Y(n_4285));
 INVxp67_ASAP7_75t_R g215884 (.A(n_4284),
    .Y(n_4283));
 INVx1_ASAP7_75t_L g215885 (.A(n_4282),
    .Y(n_4281));
 INVx2_ASAP7_75t_L g215886 (.A(n_4280),
    .Y(n_4279));
 INVx2_ASAP7_75t_L g215887 (.A(n_4278),
    .Y(n_4277));
 NAND2xp5_ASAP7_75t_R g215888 (.A(n_1550),
    .B(n_3484),
    .Y(n_4276));
 AND2x2_ASAP7_75t_R g215889 (.A(n_2707),
    .B(n_3110),
    .Y(n_4275));
 NOR2xp33_ASAP7_75t_R g215890 (.A(n_3142),
    .B(n_3686),
    .Y(n_4274));
 NAND2xp33_ASAP7_75t_R g215891 (.A(n_3477),
    .B(n_3011),
    .Y(n_4273));
 NOR2xp33_ASAP7_75t_L g215892 (.A(n_3689),
    .B(n_1553),
    .Y(n_4272));
 NOR2xp33_ASAP7_75t_R g215893 (.A(n_3349),
    .B(n_3463),
    .Y(n_4271));
 NOR2xp33_ASAP7_75t_SL g215894 (.A(n_3159),
    .B(n_3658),
    .Y(n_4270));
 NOR2xp33_ASAP7_75t_SL g215895 (.A(n_3173),
    .B(n_3651),
    .Y(n_4269));
 AND2x2_ASAP7_75t_R g215896 (.A(n_2645),
    .B(n_2940),
    .Y(n_4268));
 NOR2xp33_ASAP7_75t_R g215897 (.A(n_3616),
    .B(n_1389),
    .Y(n_4267));
 NOR2xp33_ASAP7_75t_R g215898 (.A(n_2141),
    .B(n_3424),
    .Y(n_4266));
 NAND2xp33_ASAP7_75t_R g215899 (.A(n_2128),
    .B(n_3432),
    .Y(n_4265));
 NOR2xp33_ASAP7_75t_R g215900 (.A(n_2887),
    .B(n_2068),
    .Y(n_4264));
 NAND2xp5_ASAP7_75t_L g215901 (.A(n_1456),
    .B(n_1753),
    .Y(n_4263));
 NAND2xp5_ASAP7_75t_L g215902 (.A(n_3291),
    .B(n_2509),
    .Y(n_4706));
 NOR2xp33_ASAP7_75t_R g215903 (.A(n_2143),
    .B(n_2885),
    .Y(n_4262));
 NOR2xp33_ASAP7_75t_R g215904 (.A(n_2992),
    .B(n_2911),
    .Y(n_4261));
 OAI21xp33_ASAP7_75t_R g215905 (.A1(n_2489),
    .A2(n_2590),
    .B(sa00[3]),
    .Y(n_4260));
 OAI21xp5_ASAP7_75t_L g215906 (.A1(n_2472),
    .A2(n_2591),
    .B(sa11[3]),
    .Y(n_4259));
 AND2x2_ASAP7_75t_R g215907 (.A(n_3574),
    .B(n_2421),
    .Y(n_4258));
 NOR2xp33_ASAP7_75t_R g215908 (.A(n_1860),
    .B(n_3301),
    .Y(n_4257));
 NOR2xp33_ASAP7_75t_R g215909 (.A(n_2045),
    .B(n_1755),
    .Y(n_4256));
 NOR2xp33_ASAP7_75t_R g215910 (.A(n_2096),
    .B(n_3551),
    .Y(n_4255));
 OAI21xp33_ASAP7_75t_R g215911 (.A1(n_2158),
    .A2(n_2449),
    .B(n_1411),
    .Y(n_4254));
 NOR2xp33_ASAP7_75t_R g215912 (.A(n_2513),
    .B(n_3071),
    .Y(n_4253));
 NOR2xp33_ASAP7_75t_R g215913 (.A(n_3434),
    .B(n_3517),
    .Y(n_4252));
 NAND2xp5_ASAP7_75t_L g215914 (.A(n_3017),
    .B(n_2167),
    .Y(n_4251));
 NAND2xp33_ASAP7_75t_R g215915 (.A(n_2169),
    .B(n_2883),
    .Y(n_4250));
 NAND2xp33_ASAP7_75t_R g215916 (.A(n_1721),
    .B(n_2692),
    .Y(n_4249));
 NOR2xp33_ASAP7_75t_L g215917 (.A(n_2535),
    .B(n_3045),
    .Y(n_4248));
 NAND2xp5_ASAP7_75t_R g215918 (.A(n_1406),
    .B(n_1742),
    .Y(n_4247));
 NOR2xp33_ASAP7_75t_L g215919 (.A(n_2240),
    .B(n_2879),
    .Y(n_4246));
 NAND2xp33_ASAP7_75t_R g215920 (.A(n_2817),
    .B(n_2938),
    .Y(n_4245));
 NAND2xp33_ASAP7_75t_R g215921 (.A(n_2785),
    .B(n_2574),
    .Y(n_4244));
 NAND2xp33_ASAP7_75t_R g215922 (.A(n_3347),
    .B(n_1633),
    .Y(n_4243));
 NOR2xp33_ASAP7_75t_R g215923 (.A(n_2838),
    .B(n_2932),
    .Y(n_4242));
 NAND2xp33_ASAP7_75t_R g215924 (.A(n_3302),
    .B(n_2557),
    .Y(n_4241));
 NOR2xp33_ASAP7_75t_R g215925 (.A(n_2126),
    .B(n_2877),
    .Y(n_4240));
 NAND2xp33_ASAP7_75t_R g215926 (.A(n_2543),
    .B(n_3243),
    .Y(n_4239));
 NOR2xp33_ASAP7_75t_R g215927 (.A(n_2548),
    .B(n_3279),
    .Y(n_4238));
 NOR2xp33_ASAP7_75t_R g215928 (.A(n_2570),
    .B(n_2839),
    .Y(n_4237));
 NAND2xp5_ASAP7_75t_L g215929 (.A(n_3579),
    .B(n_3199),
    .Y(n_4236));
 AND2x2_ASAP7_75t_L g215930 (.A(n_3212),
    .B(n_1572),
    .Y(n_4235));
 NOR2xp33_ASAP7_75t_L g215931 (.A(n_3198),
    .B(n_2091),
    .Y(n_4234));
 NOR2xp33_ASAP7_75t_R g215932 (.A(n_3441),
    .B(n_3293),
    .Y(n_4233));
 NOR2xp33_ASAP7_75t_R g215933 (.A(n_2063),
    .B(n_3155),
    .Y(n_4232));
 NOR2xp33_ASAP7_75t_R g215934 (.A(n_2222),
    .B(n_2909),
    .Y(n_4231));
 NAND2xp33_ASAP7_75t_R g215935 (.A(n_1497),
    .B(n_2848),
    .Y(n_4230));
 NOR2xp33_ASAP7_75t_R g215936 (.A(n_2594),
    .B(n_3288),
    .Y(n_4229));
 NOR2xp33_ASAP7_75t_R g215937 (.A(n_2074),
    .B(n_3728),
    .Y(n_4228));
 AND2x2_ASAP7_75t_R g215938 (.A(n_2090),
    .B(n_3606),
    .Y(n_4227));
 NOR2xp33_ASAP7_75t_R g215939 (.A(n_2088),
    .B(n_3182),
    .Y(n_4226));
 AND2x2_ASAP7_75t_L g215940 (.A(n_1424),
    .B(n_3611),
    .Y(n_4225));
 NOR2xp33_ASAP7_75t_L g215941 (.A(n_2858),
    .B(n_3032),
    .Y(n_4224));
 NOR2xp33_ASAP7_75t_R g215942 (.A(n_2453),
    .B(n_3207),
    .Y(n_4223));
 NAND2xp33_ASAP7_75t_R g215943 (.A(n_3380),
    .B(n_2917),
    .Y(n_4222));
 NOR2xp33_ASAP7_75t_R g215944 (.A(n_2438),
    .B(n_3111),
    .Y(n_4221));
 NAND2xp33_ASAP7_75t_R g215945 (.A(n_1659),
    .B(n_1755),
    .Y(n_4705));
 OR2x2_ASAP7_75t_SL g215946 (.A(n_2419),
    .B(n_3487),
    .Y(n_4704));
 NAND2xp5_ASAP7_75t_R g215947 (.A(n_2060),
    .B(n_1752),
    .Y(n_4703));
 NOR2xp67_ASAP7_75t_L g215948 (.A(n_2080),
    .B(n_1752),
    .Y(n_4701));
 OR2x2_ASAP7_75t_L g215949 (.A(n_3323),
    .B(n_3526),
    .Y(n_4700));
 NAND2xp5_ASAP7_75t_R g215950 (.A(n_2425),
    .B(n_3700),
    .Y(n_4699));
 NAND2xp5_ASAP7_75t_R g215951 (.A(n_3474),
    .B(n_3597),
    .Y(n_4697));
 NAND2xp5_ASAP7_75t_R g215952 (.A(n_3393),
    .B(n_2509),
    .Y(n_4696));
 NAND2xp5_ASAP7_75t_R g215953 (.A(n_3326),
    .B(n_3532),
    .Y(n_4694));
 NAND2xp33_ASAP7_75t_R g215954 (.A(n_3314),
    .B(n_2444),
    .Y(n_4692));
 NOR2xp33_ASAP7_75t_SL g215955 (.A(n_3633),
    .B(n_2063),
    .Y(n_4691));
 NAND2xp33_ASAP7_75t_R g215956 (.A(n_1641),
    .B(n_3534),
    .Y(n_4690));
 NAND2xp5_ASAP7_75t_L g215957 (.A(n_1664),
    .B(n_3599),
    .Y(n_4689));
 NOR2xp67_ASAP7_75t_R g215958 (.A(n_2393),
    .B(n_3497),
    .Y(n_4688));
 NOR2xp33_ASAP7_75t_L g215959 (.A(n_3628),
    .B(n_1342),
    .Y(n_4687));
 NAND2xp5_ASAP7_75t_R g215960 (.A(n_3528),
    .B(n_8719),
    .Y(n_4685));
 NAND2xp5_ASAP7_75t_R g215961 (.A(n_3393),
    .B(n_3533),
    .Y(n_4683));
 NOR2xp33_ASAP7_75t_SL g215962 (.A(n_3490),
    .B(n_3079),
    .Y(n_4682));
 NOR2xp33_ASAP7_75t_R g215963 (.A(n_2052),
    .B(n_3527),
    .Y(n_4681));
 NAND2xp5_ASAP7_75t_R g215964 (.A(n_2397),
    .B(n_3491),
    .Y(n_4680));
 NOR2xp33_ASAP7_75t_L g215965 (.A(n_3569),
    .B(n_3489),
    .Y(n_4679));
 NOR2xp33_ASAP7_75t_L g215966 (.A(n_3564),
    .B(n_3514),
    .Y(n_4678));
 NAND2xp5_ASAP7_75t_R g215967 (.A(n_1682),
    .B(n_3306),
    .Y(n_4676));
 NOR2xp33_ASAP7_75t_L g215968 (.A(n_2507),
    .B(n_3366),
    .Y(n_4674));
 NOR2xp33_ASAP7_75t_L g215969 (.A(n_2399),
    .B(n_3488),
    .Y(n_4673));
 NOR2xp33_ASAP7_75t_R g215970 (.A(sa02[1]),
    .B(n_3111),
    .Y(n_4220));
 OAI21xp33_ASAP7_75t_R g215971 (.A1(n_2001),
    .A2(n_2504),
    .B(n_1615),
    .Y(n_4672));
 NAND2xp5_ASAP7_75t_R g215972 (.A(n_1663),
    .B(n_3322),
    .Y(n_4670));
 NOR2xp33_ASAP7_75t_L g215973 (.A(n_3261),
    .B(n_3461),
    .Y(n_4669));
 NOR2x1_ASAP7_75t_SL g215974 (.A(n_3288),
    .B(n_3461),
    .Y(n_4668));
 NOR2xp33_ASAP7_75t_R g215975 (.A(n_2447),
    .B(n_2825),
    .Y(n_4667));
 AND2x2_ASAP7_75t_L g215976 (.A(n_2394),
    .B(n_3485),
    .Y(n_4666));
 NOR2xp67_ASAP7_75t_SL g215977 (.A(n_3305),
    .B(n_3459),
    .Y(n_4665));
 NAND2xp5_ASAP7_75t_L g215978 (.A(n_3458),
    .B(n_3304),
    .Y(n_4664));
 NAND2xp5_ASAP7_75t_L g215979 (.A(n_2401),
    .B(n_3731),
    .Y(n_4663));
 NOR2xp33_ASAP7_75t_SL g215980 (.A(n_3535),
    .B(n_3036),
    .Y(n_4662));
 NAND2xp5_ASAP7_75t_R g215981 (.A(sa10[4]),
    .B(n_3273),
    .Y(n_4661));
 NAND2xp33_ASAP7_75t_L g215982 (.A(n_3429),
    .B(n_2211),
    .Y(n_4660));
 AND2x2_ASAP7_75t_SL g215983 (.A(n_1758),
    .B(n_1755),
    .Y(n_4659));
 NAND2xp5_ASAP7_75t_L g215984 (.A(n_2132),
    .B(n_3415),
    .Y(n_4657));
 NAND2xp5_ASAP7_75t_L g215985 (.A(n_3486),
    .B(n_3536),
    .Y(n_4655));
 NAND2xp5_ASAP7_75t_SL g215986 (.A(n_2387),
    .B(n_3586),
    .Y(n_4654));
 NOR2xp33_ASAP7_75t_L g215987 (.A(n_2489),
    .B(n_3298),
    .Y(n_4652));
 NOR2xp33_ASAP7_75t_L g215988 (.A(n_3566),
    .B(n_3497),
    .Y(n_1787));
 NAND2xp5_ASAP7_75t_L g215989 (.A(sa12[4]),
    .B(n_3274),
    .Y(n_4651));
 NAND2xp33_ASAP7_75t_R g215990 (.A(n_2130),
    .B(n_3686),
    .Y(n_4650));
 NOR2xp33_ASAP7_75t_L g215991 (.A(n_2513),
    .B(n_2860),
    .Y(n_4648));
 NOR2xp33_ASAP7_75t_L g215992 (.A(n_3529),
    .B(n_3641),
    .Y(n_4647));
 NOR2xp33_ASAP7_75t_L g215993 (.A(n_1342),
    .B(n_3591),
    .Y(n_4645));
 NOR2xp33_ASAP7_75t_L g215994 (.A(n_2088),
    .B(n_3483),
    .Y(n_4643));
 NAND2xp5_ASAP7_75t_L g215995 (.A(n_1657),
    .B(n_3580),
    .Y(n_4642));
 NOR2xp33_ASAP7_75t_SL g215996 (.A(n_1575),
    .B(n_3560),
    .Y(n_4641));
 NOR2xp33_ASAP7_75t_R g215997 (.A(n_2513),
    .B(n_2872),
    .Y(n_4640));
 NOR2x1_ASAP7_75t_L g215998 (.A(n_3527),
    .B(n_3542),
    .Y(n_4639));
 NAND2xp33_ASAP7_75t_R g215999 (.A(n_2494),
    .B(n_2845),
    .Y(n_4638));
 NAND2xp5_ASAP7_75t_R g216000 (.A(n_3432),
    .B(n_2122),
    .Y(n_4637));
 NOR2xp33_ASAP7_75t_L g216001 (.A(n_3295),
    .B(n_3504),
    .Y(n_4636));
 NAND2xp33_ASAP7_75t_R g216002 (.A(n_2519),
    .B(n_3380),
    .Y(n_4635));
 NAND2xp5_ASAP7_75t_L g216003 (.A(n_3491),
    .B(n_3552),
    .Y(n_4633));
 NAND2xp5_ASAP7_75t_R g216004 (.A(n_3499),
    .B(n_1730),
    .Y(n_4631));
 NOR2xp67_ASAP7_75t_SL g216005 (.A(n_2846),
    .B(n_3498),
    .Y(n_4629));
 NAND2xp5_ASAP7_75t_L g216006 (.A(n_3308),
    .B(n_3512),
    .Y(n_4628));
 NOR2xp33_ASAP7_75t_R g216007 (.A(n_2141),
    .B(n_3687),
    .Y(n_4627));
 NAND3xp33_ASAP7_75t_R g216008 (.A(n_2410),
    .B(n_2585),
    .C(n_1477),
    .Y(n_4625));
 NAND2xp5_ASAP7_75t_L g216009 (.A(n_3447),
    .B(n_3253),
    .Y(n_4623));
 NOR2xp33_ASAP7_75t_L g216010 (.A(n_3562),
    .B(n_3488),
    .Y(n_1786));
 NOR2xp33_ASAP7_75t_SL g216011 (.A(n_3301),
    .B(n_3500),
    .Y(n_4622));
 NAND2xp33_ASAP7_75t_SL g216012 (.A(n_3501),
    .B(n_3247),
    .Y(n_4621));
 NAND2xp5_ASAP7_75t_R g216014 (.A(n_2536),
    .B(n_2827),
    .Y(n_4618));
 NAND2xp5_ASAP7_75t_R g216015 (.A(n_2814),
    .B(n_1387),
    .Y(n_4617));
 NAND2xp33_ASAP7_75t_R g216016 (.A(n_1952),
    .B(n_2815),
    .Y(n_4219));
 NOR2xp33_ASAP7_75t_L g216017 (.A(n_3299),
    .B(n_3504),
    .Y(n_4615));
 NAND2xp5_ASAP7_75t_L g216018 (.A(n_2077),
    .B(n_3533),
    .Y(n_4613));
 NOR2xp33_ASAP7_75t_L g216019 (.A(n_2063),
    .B(n_3533),
    .Y(n_4612));
 NAND2xp5_ASAP7_75t_L g216020 (.A(n_3685),
    .B(n_3485),
    .Y(n_4611));
 AND2x2_ASAP7_75t_R g216021 (.A(n_2100),
    .B(n_3678),
    .Y(n_4610));
 NAND2xp33_ASAP7_75t_R g216022 (.A(n_3627),
    .B(n_2127),
    .Y(n_4609));
 NAND2xp5_ASAP7_75t_SL g216023 (.A(n_1425),
    .B(n_1732),
    .Y(n_4608));
 NOR2xp33_ASAP7_75t_L g216024 (.A(n_1582),
    .B(n_3555),
    .Y(n_4607));
 NAND2xp33_ASAP7_75t_R g216025 (.A(n_2157),
    .B(n_3660),
    .Y(n_4606));
 NOR2xp33_ASAP7_75t_L g216026 (.A(n_3244),
    .B(n_3511),
    .Y(n_4604));
 NAND2xp33_ASAP7_75t_R g216027 (.A(n_3387),
    .B(n_2527),
    .Y(n_4603));
 NOR2xp33_ASAP7_75t_R g216028 (.A(n_3525),
    .B(n_3282),
    .Y(n_4218));
 NOR2xp67_ASAP7_75t_L g216029 (.A(n_3492),
    .B(n_3311),
    .Y(n_4602));
 AND2x2_ASAP7_75t_SL g216030 (.A(n_2060),
    .B(n_3573),
    .Y(n_4601));
 NOR2xp33_ASAP7_75t_R g216031 (.A(n_3693),
    .B(n_3463),
    .Y(n_4600));
 NAND2xp33_ASAP7_75t_R g216032 (.A(n_1683),
    .B(n_3278),
    .Y(n_4598));
 NAND2xp33_ASAP7_75t_R g216033 (.A(n_3287),
    .B(n_2537),
    .Y(n_4596));
 NAND2xp5_ASAP7_75t_L g216034 (.A(n_2456),
    .B(n_3396),
    .Y(n_4594));
 NAND2xp33_ASAP7_75t_R g216035 (.A(n_2525),
    .B(n_3329),
    .Y(n_4593));
 NAND2xp5_ASAP7_75t_R g216036 (.A(n_3281),
    .B(n_2534),
    .Y(n_4592));
 NOR2xp67_ASAP7_75t_SL g216037 (.A(n_3492),
    .B(n_3259),
    .Y(n_4590));
 NOR2xp33_ASAP7_75t_R g216038 (.A(n_1503),
    .B(n_2817),
    .Y(n_4217));
 NOR2xp33_ASAP7_75t_R g216039 (.A(n_3471),
    .B(n_3277),
    .Y(n_4589));
 NAND2xp33_ASAP7_75t_R g216040 (.A(n_3396),
    .B(n_1689),
    .Y(n_4587));
 NAND2xp5_ASAP7_75t_R g216041 (.A(n_3692),
    .B(n_3468),
    .Y(n_4585));
 NOR2xp33_ASAP7_75t_L g216042 (.A(n_3315),
    .B(n_2941),
    .Y(n_4583));
 NOR2xp33_ASAP7_75t_L g216043 (.A(n_1368),
    .B(n_2792),
    .Y(n_4582));
 NAND2xp33_ASAP7_75t_R g216044 (.A(n_1368),
    .B(n_2792),
    .Y(n_4216));
 NAND2xp5_ASAP7_75t_R g216045 (.A(n_3495),
    .B(n_2805),
    .Y(n_4581));
 NOR2xp67_ASAP7_75t_L g216046 (.A(n_2842),
    .B(n_3494),
    .Y(n_4579));
 NAND2xp33_ASAP7_75t_R g216047 (.A(n_1745),
    .B(n_3260),
    .Y(n_4577));
 OR2x2_ASAP7_75t_L g216048 (.A(n_3476),
    .B(n_2856),
    .Y(n_4576));
 NOR2xp33_ASAP7_75t_L g216049 (.A(n_2057),
    .B(n_3448),
    .Y(n_4575));
 NAND2xp5_ASAP7_75t_L g216050 (.A(n_1622),
    .B(n_3719),
    .Y(n_4574));
 NOR2xp33_ASAP7_75t_L g216051 (.A(n_1588),
    .B(n_3449),
    .Y(n_1785));
 NOR2xp67_ASAP7_75t_L g216052 (.A(n_3307),
    .B(n_1722),
    .Y(n_4572));
 NOR2xp33_ASAP7_75t_L g216053 (.A(n_2919),
    .B(n_2780),
    .Y(n_4571));
 NAND2xp5_ASAP7_75t_R g216054 (.A(n_1413),
    .B(n_3369),
    .Y(n_4215));
 NOR2xp33_ASAP7_75t_L g216055 (.A(n_2799),
    .B(n_2941),
    .Y(n_4570));
 NOR2xp33_ASAP7_75t_L g216056 (.A(n_2935),
    .B(n_2834),
    .Y(n_4569));
 NOR2xp67_ASAP7_75t_SL g216057 (.A(n_2853),
    .B(n_2934),
    .Y(n_4567));
 NOR2xp33_ASAP7_75t_L g216058 (.A(n_2935),
    .B(n_2786),
    .Y(n_4566));
 NOR2xp33_ASAP7_75t_R g216059 (.A(n_2173),
    .B(n_3619),
    .Y(n_4564));
 NOR2x1_ASAP7_75t_R g216060 (.A(n_2778),
    .B(n_2934),
    .Y(n_4563));
 NOR2xp33_ASAP7_75t_R g216061 (.A(n_1672),
    .B(n_2853),
    .Y(n_4561));
 OR2x2_ASAP7_75t_R g216062 (.A(n_2187),
    .B(n_3629),
    .Y(n_4560));
 NAND2xp5_ASAP7_75t_L g216063 (.A(n_2851),
    .B(n_1691),
    .Y(n_4558));
 NAND2xp5_ASAP7_75t_R g216064 (.A(n_2142),
    .B(n_3635),
    .Y(n_4557));
 NAND2xp5_ASAP7_75t_R g216065 (.A(n_2389),
    .B(n_3474),
    .Y(n_4556));
 NOR2xp33_ASAP7_75t_R g216066 (.A(n_2168),
    .B(n_3620),
    .Y(n_4555));
 NOR2xp33_ASAP7_75t_R g216067 (.A(n_2532),
    .B(n_3417),
    .Y(n_4554));
 NAND2xp5_ASAP7_75t_L g216068 (.A(n_2807),
    .B(n_2939),
    .Y(n_4553));
 NAND2xp5_ASAP7_75t_L g216069 (.A(n_2820),
    .B(n_1748),
    .Y(n_4552));
 NAND2xp33_ASAP7_75t_R g216070 (.A(n_2001),
    .B(n_3215),
    .Y(n_4214));
 NOR2xp33_ASAP7_75t_R g216071 (.A(n_2472),
    .B(n_2842),
    .Y(n_4550));
 NAND2xp5_ASAP7_75t_R g216072 (.A(n_2431),
    .B(n_3695),
    .Y(n_4549));
 NAND2xp5_ASAP7_75t_R g216073 (.A(n_1348),
    .B(n_3386),
    .Y(n_4547));
 NOR2xp33_ASAP7_75t_R g216074 (.A(n_2465),
    .B(n_3301),
    .Y(n_4546));
 NAND2xp33_ASAP7_75t_R g216075 (.A(n_2128),
    .B(n_3637),
    .Y(n_4213));
 NOR2xp33_ASAP7_75t_R g216076 (.A(n_2864),
    .B(n_2572),
    .Y(n_4545));
 NAND2xp5_ASAP7_75t_R g216077 (.A(n_1670),
    .B(n_1734),
    .Y(n_4543));
 NAND2xp33_ASAP7_75t_R g216078 (.A(n_2065),
    .B(n_3539),
    .Y(n_4542));
 NOR2xp33_ASAP7_75t_L g216079 (.A(n_2423),
    .B(n_3708),
    .Y(n_4540));
 NOR2xp33_ASAP7_75t_L g216080 (.A(n_2832),
    .B(n_3503),
    .Y(n_4539));
 NOR2xp33_ASAP7_75t_L g216081 (.A(n_3490),
    .B(n_1357),
    .Y(n_4212));
 NAND2xp5_ASAP7_75t_R g216082 (.A(n_1446),
    .B(n_3356),
    .Y(n_4211));
 NOR2xp33_ASAP7_75t_L g216083 (.A(n_1601),
    .B(n_3424),
    .Y(n_4538));
 NAND2xp5_ASAP7_75t_L g216084 (.A(n_1627),
    .B(n_3435),
    .Y(n_4537));
 NOR2xp33_ASAP7_75t_SL g216085 (.A(n_2073),
    .B(n_3519),
    .Y(n_4536));
 NOR2xp67_ASAP7_75t_L g216086 (.A(n_1644),
    .B(n_3514),
    .Y(n_4534));
 NOR2xp33_ASAP7_75t_R g216087 (.A(n_1678),
    .B(n_3356),
    .Y(n_4533));
 NAND2xp5_ASAP7_75t_L g216088 (.A(n_3334),
    .B(n_2886),
    .Y(n_4532));
 OR2x2_ASAP7_75t_R g216089 (.A(n_1580),
    .B(n_3546),
    .Y(n_4531));
 NOR2xp33_ASAP7_75t_L g216090 (.A(n_1553),
    .B(n_3489),
    .Y(n_4530));
 NAND2xp5_ASAP7_75t_SL g216091 (.A(n_1569),
    .B(n_1757),
    .Y(n_4529));
 NOR2xp33_ASAP7_75t_L g216092 (.A(n_2433),
    .B(n_3316),
    .Y(n_4527));
 OR2x2_ASAP7_75t_L g216093 (.A(n_2056),
    .B(n_1756),
    .Y(n_4526));
 NOR3xp33_ASAP7_75t_R g216094 (.A(n_2428),
    .B(n_2501),
    .C(n_1470),
    .Y(n_4525));
 NOR2xp33_ASAP7_75t_SL g216095 (.A(n_2839),
    .B(n_2928),
    .Y(n_4524));
 NAND2xp33_ASAP7_75t_R g216096 (.A(n_2788),
    .B(n_2929),
    .Y(n_4523));
 NAND2xp5_ASAP7_75t_L g216097 (.A(n_2075),
    .B(n_2887),
    .Y(n_4522));
 NAND2xp33_ASAP7_75t_R g216098 (.A(n_1372),
    .B(n_3515),
    .Y(n_4210));
 NOR2xp33_ASAP7_75t_R g216099 (.A(n_2487),
    .B(n_3322),
    .Y(n_4521));
 NAND2xp5_ASAP7_75t_L g216100 (.A(n_1589),
    .B(n_3675),
    .Y(n_4520));
 NAND2xp5_ASAP7_75t_SL g216101 (.A(n_2494),
    .B(n_3385),
    .Y(n_4519));
 NAND2xp5_ASAP7_75t_R g216102 (.A(n_2139),
    .B(n_1750),
    .Y(n_4517));
 NAND2xp33_ASAP7_75t_R g216103 (.A(n_2840),
    .B(n_1680),
    .Y(n_4516));
 NOR2xp33_ASAP7_75t_SL g216104 (.A(n_2499),
    .B(n_3349),
    .Y(n_4514));
 NOR2x1_ASAP7_75t_L g216105 (.A(n_1681),
    .B(n_3347),
    .Y(n_4513));
 NAND2xp5_ASAP7_75t_L g216106 (.A(n_1683),
    .B(n_3370),
    .Y(n_4510));
 NAND2xp5_ASAP7_75t_L g216107 (.A(n_3516),
    .B(n_3416),
    .Y(n_4509));
 AND2x2_ASAP7_75t_L g216108 (.A(n_2444),
    .B(n_3374),
    .Y(n_4508));
 NOR2xp33_ASAP7_75t_L g216109 (.A(n_2586),
    .B(n_3298),
    .Y(n_4506));
 NOR2xp33_ASAP7_75t_SL g216110 (.A(n_2588),
    .B(n_2797),
    .Y(n_4504));
 NAND2xp33_ASAP7_75t_R g216111 (.A(n_2587),
    .B(n_3314),
    .Y(n_4503));
 NAND2xp5_ASAP7_75t_R g216112 (.A(n_3354),
    .B(n_1686),
    .Y(n_4501));
 NAND2xp5_ASAP7_75t_R g216113 (.A(n_1735),
    .B(n_2462),
    .Y(n_4499));
 AND2x2_ASAP7_75t_L g216114 (.A(n_2427),
    .B(n_3382),
    .Y(n_4498));
 NAND2xp5_ASAP7_75t_L g216115 (.A(n_2065),
    .B(n_3343),
    .Y(n_4497));
 NOR2xp33_ASAP7_75t_SL g216116 (.A(n_1676),
    .B(n_3332),
    .Y(n_4496));
 NAND2xp5_ASAP7_75t_L g216117 (.A(n_2420),
    .B(n_3390),
    .Y(n_4495));
 NOR2x1_ASAP7_75t_L g216118 (.A(n_1671),
    .B(n_3368),
    .Y(n_4494));
 NAND2xp5_ASAP7_75t_R g216119 (.A(n_2413),
    .B(n_1737),
    .Y(n_4493));
 NOR2xp33_ASAP7_75t_L g216120 (.A(n_2584),
    .B(n_2825),
    .Y(n_4492));
 NAND2xp5_ASAP7_75t_R g216121 (.A(n_2900),
    .B(n_3519),
    .Y(n_4491));
 NAND2xp5_ASAP7_75t_L g216122 (.A(n_2823),
    .B(n_2583),
    .Y(n_4489));
 NAND2xp5_ASAP7_75t_L g216123 (.A(n_3308),
    .B(n_2575),
    .Y(n_4488));
 AND2x2_ASAP7_75t_R g216124 (.A(n_2490),
    .B(n_1743),
    .Y(n_4487));
 NAND2xp5_ASAP7_75t_R g216125 (.A(n_1655),
    .B(n_1739),
    .Y(n_4485));
 NAND2xp5_ASAP7_75t_SL g216126 (.A(n_2435),
    .B(n_1740),
    .Y(n_4484));
 NAND2xp5_ASAP7_75t_R g216127 (.A(n_3546),
    .B(n_2865),
    .Y(n_4483));
 NAND2xp5_ASAP7_75t_R g216128 (.A(n_1741),
    .B(n_2466),
    .Y(n_4482));
 NAND2xp5_ASAP7_75t_L g216129 (.A(n_2410),
    .B(n_3376),
    .Y(n_4481));
 NOR2xp67_ASAP7_75t_SL g216130 (.A(n_1607),
    .B(n_3299),
    .Y(n_1784));
 AND2x2_ASAP7_75t_L g216131 (.A(n_2568),
    .B(n_3306),
    .Y(n_4478));
 NOR2xp33_ASAP7_75t_SL g216132 (.A(n_3476),
    .B(n_2806),
    .Y(n_4476));
 NAND2xp5_ASAP7_75t_R g216133 (.A(n_1559),
    .B(n_3358),
    .Y(n_4475));
 NAND2xp5_ASAP7_75t_L g216134 (.A(n_2051),
    .B(n_3358),
    .Y(n_4473));
 NOR2xp67_ASAP7_75t_L g216135 (.A(n_2115),
    .B(n_3421),
    .Y(n_4470));
 NAND2xp5_ASAP7_75t_R g216136 (.A(n_2400),
    .B(n_1740),
    .Y(n_4468));
 NAND2xp33_ASAP7_75t_R g216137 (.A(n_2067),
    .B(n_1740),
    .Y(n_4467));
 AND2x2_ASAP7_75t_R g216138 (.A(n_2553),
    .B(n_3310),
    .Y(n_4466));
 NOR2xp33_ASAP7_75t_L g216139 (.A(n_3338),
    .B(n_1583),
    .Y(n_1783));
 NAND2xp5_ASAP7_75t_L g216140 (.A(n_3262),
    .B(n_2575),
    .Y(n_4464));
 NOR2xp33_ASAP7_75t_SL g216141 (.A(n_2786),
    .B(n_3503),
    .Y(n_4463));
 NOR2xp33_ASAP7_75t_SL g216142 (.A(n_3417),
    .B(n_2486),
    .Y(n_4461));
 NAND2xp5_ASAP7_75t_R g216143 (.A(n_2471),
    .B(n_1736),
    .Y(n_4459));
 NAND2xp5_ASAP7_75t_R g216144 (.A(n_2464),
    .B(n_3319),
    .Y(n_4458));
 NOR2xp33_ASAP7_75t_R g216145 (.A(n_2567),
    .B(n_2856),
    .Y(n_4455));
 NOR2xp33_ASAP7_75t_L g216146 (.A(n_2586),
    .B(n_3245),
    .Y(n_4453));
 NOR2xp33_ASAP7_75t_R g216147 (.A(n_2562),
    .B(n_2842),
    .Y(n_4451));
 NOR2x1_ASAP7_75t_L g216148 (.A(n_2562),
    .B(n_3269),
    .Y(n_4450));
 NOR2x1_ASAP7_75t_L g216149 (.A(n_3366),
    .B(n_3592),
    .Y(n_4449));
 NAND2xp5_ASAP7_75t_R g216150 (.A(n_1431),
    .B(n_3390),
    .Y(n_4448));
 NOR2xp33_ASAP7_75t_L g216151 (.A(n_3303),
    .B(n_3526),
    .Y(n_4447));
 NAND2xp5_ASAP7_75t_R g216152 (.A(n_2854),
    .B(n_2556),
    .Y(n_4445));
 NOR2x1_ASAP7_75t_R g216153 (.A(n_2555),
    .B(n_2821),
    .Y(n_4443));
 NAND2xp5_ASAP7_75t_L g216154 (.A(n_1569),
    .B(n_3358),
    .Y(n_4441));
 NAND2xp5_ASAP7_75t_L g216155 (.A(n_3276),
    .B(n_2553),
    .Y(n_1782));
 NAND2xp5_ASAP7_75t_L g216156 (.A(n_2048),
    .B(n_3343),
    .Y(n_4439));
 NAND2xp5_ASAP7_75t_L g216157 (.A(n_2046),
    .B(n_3343),
    .Y(n_4437));
 NOR2xp67_ASAP7_75t_R g216158 (.A(n_2530),
    .B(n_2846),
    .Y(n_4436));
 NAND2xp5_ASAP7_75t_SL g216159 (.A(n_3254),
    .B(n_2529),
    .Y(n_4434));
 NAND2xp5_ASAP7_75t_R g216160 (.A(n_3380),
    .B(n_3560),
    .Y(n_4432));
 NAND2xp5_ASAP7_75t_R g216161 (.A(n_3532),
    .B(n_3300),
    .Y(n_4430));
 NAND2xp33_ASAP7_75t_R g216162 (.A(n_2514),
    .B(n_3324),
    .Y(n_4429));
 NOR2xp33_ASAP7_75t_L g216163 (.A(n_2515),
    .B(n_3305),
    .Y(n_4428));
 AND2x2_ASAP7_75t_SL g216164 (.A(n_2416),
    .B(n_3392),
    .Y(n_4425));
 NAND2xp5_ASAP7_75t_R g216165 (.A(n_2055),
    .B(n_3376),
    .Y(n_4424));
 NAND2xp5_ASAP7_75t_L g216166 (.A(n_3387),
    .B(n_3455),
    .Y(n_4423));
 NAND2xp5_ASAP7_75t_R g216167 (.A(n_1653),
    .B(n_3376),
    .Y(n_4422));
 NAND2xp5_ASAP7_75t_L g216168 (.A(n_2429),
    .B(n_1739),
    .Y(n_4420));
 NOR2xp33_ASAP7_75t_L g216169 (.A(n_2045),
    .B(n_1738),
    .Y(n_4419));
 NOR2xp33_ASAP7_75t_L g216170 (.A(n_2517),
    .B(n_3295),
    .Y(n_4417));
 NAND2xp5_ASAP7_75t_R g216171 (.A(n_3304),
    .B(n_2159),
    .Y(n_4416));
 NAND2xp5_ASAP7_75t_R g216172 (.A(n_1953),
    .B(n_3275),
    .Y(n_4415));
 NAND2xp5_ASAP7_75t_R g216173 (.A(n_3289),
    .B(n_2505),
    .Y(n_4413));
 NOR2xp33_ASAP7_75t_L g216174 (.A(n_2506),
    .B(n_3285),
    .Y(n_4411));
 NAND2xp5_ASAP7_75t_R g216175 (.A(n_2840),
    .B(n_2540),
    .Y(n_4410));
 NAND2xp5_ASAP7_75t_R g216176 (.A(n_1687),
    .B(n_1733),
    .Y(n_4409));
 NAND2xp5_ASAP7_75t_R g216177 (.A(n_1505),
    .B(n_1726),
    .Y(n_4408));
 NAND2xp5_ASAP7_75t_L g216178 (.A(n_2397),
    .B(n_3382),
    .Y(n_4407));
 NAND2xp5_ASAP7_75t_R g216179 (.A(n_3265),
    .B(n_1856),
    .Y(n_4405));
 NOR2x1_ASAP7_75t_R g216180 (.A(n_2539),
    .B(n_2818),
    .Y(n_4404));
 NOR2xp33_ASAP7_75t_L g216181 (.A(n_3471),
    .B(n_3259),
    .Y(n_4403));
 NOR2xp33_ASAP7_75t_R g216182 (.A(sa22[4]),
    .B(n_2782),
    .Y(n_4402));
 NOR2xp33_ASAP7_75t_L g216183 (.A(n_2577),
    .B(n_3454),
    .Y(n_4400));
 NOR2xp33_ASAP7_75t_R g216184 (.A(n_2577),
    .B(n_2871),
    .Y(n_4399));
 NAND2xp5_ASAP7_75t_R g216185 (.A(n_3396),
    .B(n_3483),
    .Y(n_4398));
 NAND2xp5_ASAP7_75t_R g216186 (.A(n_2488),
    .B(n_3289),
    .Y(n_4396));
 NAND2xp5_ASAP7_75t_SL g216187 (.A(n_2521),
    .B(n_3283),
    .Y(n_4394));
 NOR2xp33_ASAP7_75t_R g216188 (.A(n_2522),
    .B(n_3301),
    .Y(n_4393));
 NOR2xp33_ASAP7_75t_R g216189 (.A(n_2517),
    .B(n_3327),
    .Y(n_4392));
 NOR2xp33_ASAP7_75t_L g216190 (.A(n_2453),
    .B(n_3454),
    .Y(n_4391));
 NOR2xp33_ASAP7_75t_SL g216191 (.A(n_3327),
    .B(n_3454),
    .Y(n_4390));
 NOR2xp33_ASAP7_75t_L g216192 (.A(n_3453),
    .B(n_3454),
    .Y(n_4387));
 NAND2xp33_ASAP7_75t_R g216193 (.A(n_2803),
    .B(n_1359),
    .Y(n_4209));
 NOR2xp33_ASAP7_75t_R g216194 (.A(n_1702),
    .B(n_2797),
    .Y(n_4385));
 AND2x2_ASAP7_75t_L g216195 (.A(n_2536),
    .B(n_2900),
    .Y(n_4383));
 AND2x2_ASAP7_75t_L g216196 (.A(n_1949),
    .B(n_2790),
    .Y(n_4382));
 NOR2xp33_ASAP7_75t_SL g216197 (.A(n_3525),
    .B(n_3248),
    .Y(n_4381));
 NAND2xp5_ASAP7_75t_SL g216198 (.A(n_2835),
    .B(n_2523),
    .Y(n_1781));
 NAND2xp5_ASAP7_75t_SL g216199 (.A(n_1950),
    .B(n_3271),
    .Y(n_4380));
 NOR2xp33_ASAP7_75t_R g216200 (.A(n_1425),
    .B(n_1732),
    .Y(n_4208));
 NOR2xp33_ASAP7_75t_L g216201 (.A(sa32[4]),
    .B(n_2783),
    .Y(n_4379));
 NAND2xp5_ASAP7_75t_L g216202 (.A(n_2500),
    .B(n_3294),
    .Y(n_4378));
 NAND2xp5_ASAP7_75t_R g216203 (.A(n_2523),
    .B(n_2833),
    .Y(n_4376));
 NOR2x1_ASAP7_75t_L g216204 (.A(n_2501),
    .B(n_3256),
    .Y(n_4375));
 NAND2xp5_ASAP7_75t_R g216205 (.A(n_2502),
    .B(n_3278),
    .Y(n_4373));
 NOR2xp33_ASAP7_75t_L g216206 (.A(sa31[4]),
    .B(n_3242),
    .Y(n_4371));
 NAND2xp5_ASAP7_75t_SL g216207 (.A(n_1760),
    .B(n_2869),
    .Y(n_4369));
 NAND2x1_ASAP7_75t_SL g216208 (.A(n_2867),
    .B(n_3689),
    .Y(n_4368));
 NOR2x1_ASAP7_75t_SL g216209 (.A(n_3091),
    .B(n_2861),
    .Y(n_4366));
 NOR2xp33_ASAP7_75t_L g216210 (.A(n_2906),
    .B(n_3298),
    .Y(n_4364));
 NAND2x1_ASAP7_75t_SL g216211 (.A(n_3669),
    .B(n_1748),
    .Y(n_4362));
 NOR2x1_ASAP7_75t_L g216212 (.A(n_3307),
    .B(n_2889),
    .Y(n_4360));
 AND2x2_ASAP7_75t_SL g216213 (.A(n_3655),
    .B(n_3340),
    .Y(n_4359));
 NOR2x1_ASAP7_75t_L g216214 (.A(sa10[4]),
    .B(n_3273),
    .Y(n_4356));
 AND2x2_ASAP7_75t_L g216215 (.A(n_2895),
    .B(n_3308),
    .Y(n_4355));
 NOR2x1_ASAP7_75t_L g216216 (.A(n_2913),
    .B(n_3311),
    .Y(n_4354));
 AND2x2_ASAP7_75t_SL g216217 (.A(n_3654),
    .B(n_3406),
    .Y(n_4352));
 NAND2xp5_ASAP7_75t_L g216218 (.A(n_3644),
    .B(n_3502),
    .Y(n_4350));
 NAND2x1_ASAP7_75t_SL g216219 (.A(n_3639),
    .B(n_1746),
    .Y(n_4348));
 AND2x2_ASAP7_75t_SL g216220 (.A(n_1759),
    .B(n_3470),
    .Y(n_4347));
 NAND2xp5_ASAP7_75t_SL g216221 (.A(n_3617),
    .B(n_1745),
    .Y(n_4345));
 NAND2xp5_ASAP7_75t_L g216222 (.A(n_8200),
    .B(n_1710),
    .Y(n_4343));
 NAND2xp5_ASAP7_75t_SL g216223 (.A(n_3616),
    .B(n_3524),
    .Y(n_1780));
 NAND2xp5_ASAP7_75t_SL g216224 (.A(n_3612),
    .B(n_3532),
    .Y(n_4339));
 OR2x2_ASAP7_75t_SL g216225 (.A(n_1385),
    .B(n_2811),
    .Y(n_4338));
 NOR2x1_ASAP7_75t_L g216226 (.A(n_3614),
    .B(n_3526),
    .Y(n_4336));
 NAND2xp5_ASAP7_75t_SL g216227 (.A(n_1856),
    .B(n_3266),
    .Y(n_4333));
 AND2x2_ASAP7_75t_SL g216228 (.A(n_1425),
    .B(n_3267),
    .Y(n_4332));
 NAND2x1_ASAP7_75t_SL g216229 (.A(n_1852),
    .B(n_3242),
    .Y(n_1777));
 AND2x4_ASAP7_75t_SL g216230 (.A(n_1950),
    .B(n_3270),
    .Y(n_4330));
 NAND2xp5_ASAP7_75t_SL g216231 (.A(n_8200),
    .B(n_2794),
    .Y(n_4328));
 NAND2x1p5_ASAP7_75t_L g216232 (.A(n_8912),
    .B(n_2783),
    .Y(n_4326));
 NAND2xp5_ASAP7_75t_SL g216233 (.A(n_1855),
    .B(n_2782),
    .Y(n_4324));
 OR2x2_ASAP7_75t_SL g216234 (.A(n_1960),
    .B(n_3273),
    .Y(n_4323));
 NAND2x1_ASAP7_75t_SL g216235 (.A(sa31[4]),
    .B(n_3241),
    .Y(n_4318));
 NAND2x1p5_ASAP7_75t_SL g216236 (.A(n_2488),
    .B(n_3322),
    .Y(n_4317));
 AND2x2_ASAP7_75t_SL g216237 (.A(n_1345),
    .B(n_3317),
    .Y(n_4315));
 NOR2x1p5_ASAP7_75t_SL g216238 (.A(n_1950),
    .B(n_3270),
    .Y(n_4313));
 NAND2x1_ASAP7_75t_SL g216239 (.A(n_1853),
    .B(n_1710),
    .Y(n_1775));
 NOR2x2_ASAP7_75t_SL g216240 (.A(n_2817),
    .B(n_1944),
    .Y(n_4309));
 OR2x2_ASAP7_75t_SL g216241 (.A(n_1949),
    .B(n_2791),
    .Y(n_4307));
 OR2x2_ASAP7_75t_SL g216242 (.A(n_1856),
    .B(n_3266),
    .Y(n_4305));
 AND2x2_ASAP7_75t_SL g216243 (.A(n_1506),
    .B(n_3249),
    .Y(n_4303));
 AND2x2_ASAP7_75t_SL g216244 (.A(sa12[4]),
    .B(n_3275),
    .Y(n_4302));
 NAND2x1p5_ASAP7_75t_SL g216245 (.A(n_1675),
    .B(n_3332),
    .Y(n_4300));
 NAND2x1_ASAP7_75t_SL g216246 (.A(n_8189),
    .B(n_2793),
    .Y(n_4298));
 AND2x4_ASAP7_75t_SL g216247 (.A(n_2464),
    .B(n_3320),
    .Y(n_4296));
 OR2x2_ASAP7_75t_SL g216248 (.A(n_8189),
    .B(n_2793),
    .Y(n_4294));
 AND2x4_ASAP7_75t_L g216249 (.A(n_2462),
    .B(n_3325),
    .Y(n_4292));
 AND2x2_ASAP7_75t_SL g216250 (.A(n_1385),
    .B(n_2808),
    .Y(n_4290));
 NOR2x1_ASAP7_75t_SL g216251 (.A(n_2472),
    .B(n_1736),
    .Y(n_4288));
 NAND2x1_ASAP7_75t_SL g216252 (.A(n_1949),
    .B(n_2791),
    .Y(n_4286));
 OR2x2_ASAP7_75t_SL g216253 (.A(n_2782),
    .B(n_1855),
    .Y(n_4284));
 AND2x4_ASAP7_75t_SL g216254 (.A(n_1954),
    .B(n_2803),
    .Y(n_4282));
 NAND2x1_ASAP7_75t_SL g216255 (.A(n_8896),
    .B(n_2784),
    .Y(n_4280));
 AND2x2_ASAP7_75t_SL g216256 (.A(n_1387),
    .B(n_2815),
    .Y(n_4278));
 INVxp67_ASAP7_75t_R g216257 (.A(n_4206),
    .Y(n_4207));
 INVxp67_ASAP7_75t_R g216258 (.A(n_4201),
    .Y(n_4202));
 INVxp33_ASAP7_75t_R g216259 (.A(n_4197),
    .Y(n_4198));
 INVxp33_ASAP7_75t_R g216260 (.A(n_4190),
    .Y(n_4191));
 INVxp67_ASAP7_75t_L g216261 (.A(n_4188),
    .Y(n_4189));
 INVxp33_ASAP7_75t_R g216262 (.A(n_4184),
    .Y(n_4185));
 INVxp67_ASAP7_75t_R g216264 (.A(n_4175),
    .Y(n_4176));
 INVxp33_ASAP7_75t_R g216265 (.A(n_4173),
    .Y(n_4174));
 INVxp67_ASAP7_75t_R g216266 (.A(n_4171),
    .Y(n_4172));
 INVxp33_ASAP7_75t_R g216267 (.A(n_4169),
    .Y(n_4170));
 INVxp33_ASAP7_75t_R g216268 (.A(n_4164),
    .Y(n_4165));
 INVxp33_ASAP7_75t_R g216269 (.A(n_4160),
    .Y(n_4161));
 INVxp67_ASAP7_75t_L g216270 (.A(n_4158),
    .Y(n_4159));
 INVxp33_ASAP7_75t_R g216271 (.A(n_4152),
    .Y(n_4153));
 INVxp33_ASAP7_75t_R g216272 (.A(n_4147),
    .Y(n_4148));
 INVxp33_ASAP7_75t_R g216274 (.A(n_4144),
    .Y(n_4145));
 INVxp33_ASAP7_75t_R g216275 (.A(n_4142),
    .Y(n_4143));
 INVxp33_ASAP7_75t_R g216276 (.A(n_4132),
    .Y(n_4133));
 INVxp33_ASAP7_75t_R g216277 (.A(n_4130),
    .Y(n_4131));
 INVxp67_ASAP7_75t_L g216278 (.A(n_4127),
    .Y(n_4128));
 INVxp67_ASAP7_75t_R g216279 (.A(n_4122),
    .Y(n_4123));
 INVxp67_ASAP7_75t_L g216280 (.A(n_4120),
    .Y(n_4121));
 INVxp67_ASAP7_75t_SL g216281 (.A(n_4112),
    .Y(n_4113));
 INVxp67_ASAP7_75t_L g216282 (.A(n_4109),
    .Y(n_4110));
 INVxp67_ASAP7_75t_R g216283 (.A(n_4107),
    .Y(n_4108));
 INVxp67_ASAP7_75t_L g216284 (.A(n_4099),
    .Y(n_4100));
 INVxp33_ASAP7_75t_R g216285 (.A(n_4096),
    .Y(n_4097));
 INVxp67_ASAP7_75t_R g216287 (.A(n_4094),
    .Y(n_4095));
 INVxp33_ASAP7_75t_R g216288 (.A(n_4091),
    .Y(n_4092));
 INVxp33_ASAP7_75t_R g216289 (.A(n_4085),
    .Y(n_4086));
 INVxp33_ASAP7_75t_R g216290 (.A(n_4083),
    .Y(n_4084));
 INVxp67_ASAP7_75t_R g216291 (.A(n_4081),
    .Y(n_4082));
 INVxp67_ASAP7_75t_L g216292 (.A(n_4077),
    .Y(n_4078));
 INVxp67_ASAP7_75t_R g216293 (.A(n_4075),
    .Y(n_4076));
 INVxp67_ASAP7_75t_R g216294 (.A(n_4072),
    .Y(n_4073));
 INVxp33_ASAP7_75t_R g216295 (.A(n_4070),
    .Y(n_4071));
 INVxp67_ASAP7_75t_L g216296 (.A(n_4068),
    .Y(n_4069));
 INVxp33_ASAP7_75t_R g216297 (.A(n_4063),
    .Y(n_4064));
 INVxp33_ASAP7_75t_R g216298 (.A(n_4060),
    .Y(n_4061));
 INVxp33_ASAP7_75t_R g216299 (.A(n_4054),
    .Y(n_4055));
 INVxp67_ASAP7_75t_R g216300 (.A(n_4049),
    .Y(n_4050));
 INVxp67_ASAP7_75t_R g216301 (.A(n_4046),
    .Y(n_4047));
 INVxp33_ASAP7_75t_R g216302 (.A(n_4039),
    .Y(n_4040));
 INVxp67_ASAP7_75t_L g216304 (.A(n_4034),
    .Y(n_4035));
 INVxp33_ASAP7_75t_R g216305 (.A(n_4031),
    .Y(n_4032));
 INVxp33_ASAP7_75t_R g216306 (.A(n_4027),
    .Y(n_4028));
 INVxp67_ASAP7_75t_SL g216307 (.A(n_4023),
    .Y(n_4024));
 INVxp67_ASAP7_75t_L g216309 (.A(n_4020),
    .Y(n_4021));
 INVxp67_ASAP7_75t_R g216310 (.A(n_4018),
    .Y(n_4019));
 INVxp67_ASAP7_75t_L g216311 (.A(n_4016),
    .Y(n_4017));
 INVxp33_ASAP7_75t_R g216313 (.A(n_4012),
    .Y(n_4013));
 INVxp33_ASAP7_75t_R g216314 (.A(n_4011),
    .Y(n_4010));
 INVxp67_ASAP7_75t_R g216315 (.A(n_4008),
    .Y(n_4009));
 INVxp67_ASAP7_75t_R g216316 (.A(n_4005),
    .Y(n_4004));
 INVxp67_ASAP7_75t_R g216317 (.A(n_4003),
    .Y(n_4002));
 INVx1_ASAP7_75t_L g216318 (.A(n_4000),
    .Y(n_4001));
 INVxp67_ASAP7_75t_L g216319 (.A(n_3998),
    .Y(n_3999));
 INVxp67_ASAP7_75t_R g216320 (.A(n_3994),
    .Y(n_3995));
 INVxp33_ASAP7_75t_R g216321 (.A(n_3992),
    .Y(n_3993));
 INVxp67_ASAP7_75t_L g216322 (.A(n_3989),
    .Y(n_3990));
 INVx1_ASAP7_75t_SL g216323 (.A(n_3988),
    .Y(n_3989));
 HB1xp67_ASAP7_75t_L g216324 (.A(n_3984),
    .Y(n_3985));
 INVxp67_ASAP7_75t_R g216325 (.A(n_3982),
    .Y(n_3983));
 INVxp67_ASAP7_75t_L g216326 (.A(n_3981),
    .Y(n_3980));
 INVxp67_ASAP7_75t_L g216327 (.A(n_3977),
    .Y(n_3978));
 INVx1_ASAP7_75t_SL g216329 (.A(n_3974),
    .Y(n_3975));
 INVxp33_ASAP7_75t_R g216330 (.A(n_3972),
    .Y(n_3973));
 INVxp67_ASAP7_75t_L g216331 (.A(n_3971),
    .Y(n_3970));
 INVxp67_ASAP7_75t_R g216332 (.A(n_3968),
    .Y(n_3969));
 INVxp67_ASAP7_75t_R g216333 (.A(n_3966),
    .Y(n_3967));
 INVxp67_ASAP7_75t_SL g216334 (.A(n_3964),
    .Y(n_3965));
 INVxp33_ASAP7_75t_R g216335 (.A(n_3961),
    .Y(n_3962));
 INVxp33_ASAP7_75t_R g216336 (.A(n_3959),
    .Y(n_3960));
 INVxp67_ASAP7_75t_R g216337 (.A(n_3957),
    .Y(n_3958));
 INVxp67_ASAP7_75t_L g216338 (.A(n_3954),
    .Y(n_3955));
 INVxp33_ASAP7_75t_R g216339 (.A(n_3952),
    .Y(n_3953));
 INVxp33_ASAP7_75t_R g216340 (.A(n_3949),
    .Y(n_3950));
 INVxp67_ASAP7_75t_SL g216341 (.A(n_3948),
    .Y(n_3947));
 INVx1_ASAP7_75t_L g216342 (.A(n_3942),
    .Y(n_3943));
 INVxp33_ASAP7_75t_R g216343 (.A(n_3938),
    .Y(n_3939));
 INVxp67_ASAP7_75t_R g216344 (.A(n_3936),
    .Y(n_3937));
 INVxp33_ASAP7_75t_R g216345 (.A(n_3933),
    .Y(n_3934));
 INVx1_ASAP7_75t_L g216346 (.A(n_3931),
    .Y(n_3932));
 INVxp33_ASAP7_75t_R g216347 (.A(n_3928),
    .Y(n_3929));
 INVxp67_ASAP7_75t_R g216348 (.A(n_3922),
    .Y(n_3923));
 INVxp33_ASAP7_75t_R g216350 (.A(n_1767),
    .Y(n_3920));
 INVxp67_ASAP7_75t_R g216352 (.A(n_3918),
    .Y(n_3917));
 INVxp67_ASAP7_75t_R g216354 (.A(n_3916),
    .Y(n_3915));
 INVxp67_ASAP7_75t_R g216355 (.A(n_3914),
    .Y(n_3913));
 INVxp67_ASAP7_75t_L g216356 (.A(n_3911),
    .Y(n_3910));
 INVxp67_ASAP7_75t_R g216357 (.A(n_3909),
    .Y(n_3908));
 INVxp67_ASAP7_75t_R g216358 (.A(n_3906),
    .Y(n_3907));
 INVxp67_ASAP7_75t_R g216359 (.A(n_3904),
    .Y(n_3903));
 INVxp67_ASAP7_75t_R g216360 (.A(n_3902),
    .Y(n_3901));
 INVxp67_ASAP7_75t_R g216361 (.A(n_3900),
    .Y(n_3899));
 INVx1_ASAP7_75t_L g216363 (.A(n_3895),
    .Y(n_3896));
 INVx1_ASAP7_75t_SL g216364 (.A(n_3892),
    .Y(n_3893));
 INVx1_ASAP7_75t_L g216365 (.A(n_3890),
    .Y(n_3891));
 INVxp33_ASAP7_75t_R g216366 (.A(n_3888),
    .Y(n_3889));
 INVx1_ASAP7_75t_L g216367 (.A(n_3887),
    .Y(n_3886));
 INVx1_ASAP7_75t_L g216369 (.A(n_1763),
    .Y(n_1764));
 INVxp67_ASAP7_75t_R g216371 (.A(n_3884),
    .Y(n_3883));
 INVx1_ASAP7_75t_SL g216372 (.A(n_3882),
    .Y(n_3881));
 INVx1_ASAP7_75t_L g216373 (.A(n_3879),
    .Y(n_3878));
 INVxp67_ASAP7_75t_L g216375 (.A(n_3874),
    .Y(n_1762));
 INVxp33_ASAP7_75t_R g216376 (.A(n_3872),
    .Y(n_3873));
 INVx1_ASAP7_75t_L g216377 (.A(n_3870),
    .Y(n_3871));
 INVxp67_ASAP7_75t_R g216378 (.A(n_3868),
    .Y(n_3869));
 INVxp33_ASAP7_75t_L g216379 (.A(n_3866),
    .Y(n_3867));
 HB1xp67_ASAP7_75t_L g216380 (.A(n_3864),
    .Y(n_3865));
 INVx1_ASAP7_75t_L g216381 (.A(n_3863),
    .Y(n_3862));
 INVx1_ASAP7_75t_L g216382 (.A(n_3860),
    .Y(n_3859));
 INVx1_ASAP7_75t_L g216383 (.A(n_3858),
    .Y(n_3857));
 INVxp67_ASAP7_75t_L g216384 (.A(n_3856),
    .Y(n_3855));
 INVx1_ASAP7_75t_SL g216385 (.A(n_3854),
    .Y(n_3853));
 INVx1_ASAP7_75t_R g216388 (.A(n_1761),
    .Y(n_3852));
 INVxp67_ASAP7_75t_R g216389 (.A(n_3851),
    .Y(n_3850));
 INVx1_ASAP7_75t_R g216390 (.A(n_3848),
    .Y(n_3849));
 INVx1_ASAP7_75t_SL g216391 (.A(n_3847),
    .Y(n_3846));
 INVx2_ASAP7_75t_R g216392 (.A(n_3845),
    .Y(n_3844));
 OAI21xp33_ASAP7_75t_L g216393 (.A1(n_1358),
    .A2(n_2563),
    .B(n_3110),
    .Y(n_3843));
 NAND2xp33_ASAP7_75t_R g216394 (.A(n_2496),
    .B(n_2978),
    .Y(n_3842));
 AOI22xp33_ASAP7_75t_SL g216395 (.A1(n_2158),
    .A2(n_1561),
    .B1(n_2117),
    .B2(n_2345),
    .Y(n_3841));
 NAND2xp33_ASAP7_75t_R g216396 (.A(n_2065),
    .B(n_2960),
    .Y(n_3840));
 AOI22xp33_ASAP7_75t_R g216397 (.A1(n_2077),
    .A2(n_2282),
    .B1(n_2543),
    .B2(n_1454),
    .Y(n_3839));
 OAI21xp5_ASAP7_75t_R g216398 (.A1(n_2142),
    .A2(n_1543),
    .B(n_2762),
    .Y(n_3838));
 OAI22xp33_ASAP7_75t_R g216399 (.A1(n_1546),
    .A2(n_2172),
    .B1(n_1597),
    .B2(n_2352),
    .Y(n_3837));
 AOI22xp33_ASAP7_75t_R g216400 (.A1(n_2168),
    .A2(n_2042),
    .B1(n_1599),
    .B2(n_2349),
    .Y(n_3836));
 AOI22xp33_ASAP7_75t_R g216401 (.A1(n_1368),
    .A2(n_1577),
    .B1(n_1410),
    .B2(n_2572),
    .Y(n_3835));
 AOI22xp33_ASAP7_75t_R g216402 (.A1(n_1502),
    .A2(n_2072),
    .B1(n_1336),
    .B2(n_2535),
    .Y(n_3834));
 OAI22xp33_ASAP7_75t_R g216403 (.A1(n_1375),
    .A2(n_2078),
    .B1(n_1938),
    .B2(n_2512),
    .Y(n_3833));
 OR5x1_ASAP7_75t_R g216404 (.A(n_1928),
    .B(dcnt[3]),
    .C(dcnt[2]),
    .D(dcnt[1]),
    .E(ld),
    .Y(n_3832));
 AOI21xp33_ASAP7_75t_R g216405 (.A1(n_2440),
    .A2(n_2502),
    .B(n_2396),
    .Y(n_3831));
 OAI21xp33_ASAP7_75t_R g216406 (.A1(n_1526),
    .A2(n_1984),
    .B(n_3306),
    .Y(n_3830));
 OAI21xp33_ASAP7_75t_R g216407 (.A1(n_2437),
    .A2(n_2506),
    .B(n_2394),
    .Y(n_3829));
 NAND2xp33_ASAP7_75t_R g216408 (.A(n_3254),
    .B(n_3406),
    .Y(n_3828));
 AOI21xp5_ASAP7_75t_R g216409 (.A1(n_1467),
    .A2(n_1483),
    .B(n_3298),
    .Y(n_3827));
 OAI21xp33_ASAP7_75t_L g216410 (.A1(n_2437),
    .A2(n_2594),
    .B(n_1449),
    .Y(n_3826));
 OAI21xp33_ASAP7_75t_R g216411 (.A1(n_1499),
    .A2(n_2546),
    .B(n_3202),
    .Y(n_3825));
 AO21x1_ASAP7_75t_R g216412 (.A1(n_1395),
    .A2(n_2547),
    .B(n_3203),
    .Y(n_3824));
 OAI21xp33_ASAP7_75t_R g216413 (.A1(n_2019),
    .A2(n_1512),
    .B(n_3308),
    .Y(n_3823));
 AND3x1_ASAP7_75t_R g216414 (.A(n_1730),
    .B(n_1348),
    .C(n_2318),
    .Y(n_3822));
 OAI21xp33_ASAP7_75t_R g216415 (.A1(n_1839),
    .A2(n_2570),
    .B(n_3183),
    .Y(n_3821));
 AOI21xp33_ASAP7_75t_R g216416 (.A1(n_2100),
    .A2(n_2436),
    .B(n_1363),
    .Y(n_3820));
 AOI21xp33_ASAP7_75t_R g216417 (.A1(n_2107),
    .A2(n_2473),
    .B(n_2045),
    .Y(n_3819));
 AOI21xp33_ASAP7_75t_L g216418 (.A1(n_1675),
    .A2(n_2178),
    .B(n_1584),
    .Y(n_3818));
 NAND2xp33_ASAP7_75t_R g216419 (.A(n_2483),
    .B(n_2792),
    .Y(n_3817));
 NAND2xp33_ASAP7_75t_R g216420 (.A(n_2781),
    .B(n_2440),
    .Y(n_3816));
 OAI21xp33_ASAP7_75t_R g216421 (.A1(n_1410),
    .A2(n_2126),
    .B(n_1380),
    .Y(n_3815));
 OAI31xp33_ASAP7_75t_R g216422 (.A1(n_2126),
    .A2(n_1839),
    .A3(n_2014),
    .B(n_2415),
    .Y(n_3814));
 AOI21xp33_ASAP7_75t_R g216423 (.A1(n_2172),
    .A2(n_1933),
    .B(n_2040),
    .Y(n_3813));
 NAND2xp33_ASAP7_75t_R g216424 (.A(n_2410),
    .B(n_3058),
    .Y(n_3812));
 NAND2xp33_ASAP7_75t_R g216425 (.A(n_2796),
    .B(n_2867),
    .Y(n_3811));
 AOI21xp33_ASAP7_75t_R g216426 (.A1(n_1677),
    .A2(n_1596),
    .B(n_2073),
    .Y(n_3810));
 OAI21xp33_ASAP7_75t_L g216427 (.A1(n_2068),
    .A2(n_2558),
    .B(n_2962),
    .Y(n_3809));
 OAI21xp33_ASAP7_75t_R g216428 (.A1(n_1560),
    .A2(n_2546),
    .B(n_2994),
    .Y(n_3808));
 AOI21xp33_ASAP7_75t_R g216429 (.A1(n_1682),
    .A2(n_2103),
    .B(n_2083),
    .Y(n_3807));
 AOI21xp33_ASAP7_75t_R g216430 (.A1(n_2101),
    .A2(n_1680),
    .B(n_1580),
    .Y(n_3806));
 NAND2xp5_ASAP7_75t_L g216431 (.A(n_2414),
    .B(n_3063),
    .Y(n_3805));
 AND2x2_ASAP7_75t_L g216432 (.A(n_3053),
    .B(n_1625),
    .Y(n_3804));
 NAND2xp33_ASAP7_75t_R g216433 (.A(n_1717),
    .B(n_2779),
    .Y(n_3803));
 AOI21xp33_ASAP7_75t_R g216434 (.A1(n_2076),
    .A2(n_2543),
    .B(n_3026),
    .Y(n_3802));
 AOI21xp5_ASAP7_75t_SL g216435 (.A1(n_2060),
    .A2(n_2549),
    .B(n_1723),
    .Y(n_3801));
 OA21x2_ASAP7_75t_L g216436 (.A1(n_2552),
    .A2(n_2043),
    .B(n_2957),
    .Y(n_3800));
 AOI21xp5_ASAP7_75t_L g216437 (.A1(n_2559),
    .A2(n_2040),
    .B(n_3038),
    .Y(n_3799));
 AOI21xp33_ASAP7_75t_R g216438 (.A1(n_2579),
    .A2(n_1439),
    .B(n_3019),
    .Y(n_3798));
 AOI21xp33_ASAP7_75t_R g216439 (.A1(n_2512),
    .A2(n_2215),
    .B(n_1623),
    .Y(n_3797));
 NAND2xp5_ASAP7_75t_R g216440 (.A(n_1633),
    .B(n_3055),
    .Y(n_3796));
 NOR2xp33_ASAP7_75t_R g216441 (.A(n_1656),
    .B(n_3023),
    .Y(n_3795));
 NAND2xp33_ASAP7_75t_R g216442 (.A(n_2404),
    .B(n_3020),
    .Y(n_3794));
 AOI21xp33_ASAP7_75t_R g216443 (.A1(n_1844),
    .A2(n_1600),
    .B(n_2054),
    .Y(n_3793));
 AOI21xp33_ASAP7_75t_L g216444 (.A1(n_1670),
    .A2(n_2171),
    .B(n_1590),
    .Y(n_3792));
 OAI21xp33_ASAP7_75t_R g216445 (.A1(n_2120),
    .A2(n_2535),
    .B(n_1446),
    .Y(n_3791));
 NAND2xp33_ASAP7_75t_R g216446 (.A(n_2216),
    .B(n_1718),
    .Y(n_3790));
 AOI21xp33_ASAP7_75t_R g216447 (.A1(n_2110),
    .A2(n_2525),
    .B(n_2430),
    .Y(n_3789));
 OAI21xp33_ASAP7_75t_R g216448 (.A1(n_1454),
    .A2(n_2133),
    .B(n_1583),
    .Y(n_3788));
 OAI21xp33_ASAP7_75t_R g216449 (.A1(n_1377),
    .A2(n_2108),
    .B(n_1450),
    .Y(n_3787));
 OAI21xp33_ASAP7_75t_R g216450 (.A1(n_2199),
    .A2(n_1346),
    .B(n_1380),
    .Y(n_3786));
 AOI21xp33_ASAP7_75t_R g216451 (.A1(n_2536),
    .A2(n_2011),
    .B(n_1629),
    .Y(n_3785));
 OAI21xp33_ASAP7_75t_R g216452 (.A1(n_2280),
    .A2(n_1429),
    .B(n_3060),
    .Y(n_3784));
 OAI21xp33_ASAP7_75t_R g216453 (.A1(n_2434),
    .A2(n_2293),
    .B(n_2180),
    .Y(n_3783));
 OAI21xp33_ASAP7_75t_R g216454 (.A1(n_2327),
    .A2(n_1637),
    .B(n_2992),
    .Y(n_3782));
 OAI21xp33_ASAP7_75t_L g216455 (.A1(sa10[7]),
    .A2(n_2526),
    .B(n_1449),
    .Y(n_3781));
 OAI21xp33_ASAP7_75t_R g216456 (.A1(n_2313),
    .A2(n_1629),
    .B(n_2953),
    .Y(n_3780));
 AOI21xp33_ASAP7_75t_R g216457 (.A1(n_2249),
    .A2(n_1498),
    .B(n_1412),
    .Y(n_3779));
 OAI21xp33_ASAP7_75t_R g216458 (.A1(n_2574),
    .A2(n_2424),
    .B(sa21[0]),
    .Y(n_3778));
 AOI21xp33_ASAP7_75t_R g216459 (.A1(n_1559),
    .A2(n_2117),
    .B(n_1980),
    .Y(n_3777));
 NOR2xp33_ASAP7_75t_R g216460 (.A(n_3313),
    .B(n_3285),
    .Y(n_3776));
 AOI21xp33_ASAP7_75t_R g216461 (.A1(n_1419),
    .A2(n_2199),
    .B(sa33[0]),
    .Y(n_3775));
 OAI21xp33_ASAP7_75t_R g216462 (.A1(n_2537),
    .A2(n_1560),
    .B(n_1981),
    .Y(n_3774));
 NOR2xp33_ASAP7_75t_R g216463 (.A(n_2260),
    .B(n_3201),
    .Y(n_3773));
 AOI21xp33_ASAP7_75t_R g216464 (.A1(n_2543),
    .A2(n_2462),
    .B(n_1971),
    .Y(n_3772));
 AOI21xp33_ASAP7_75t_R g216465 (.A1(n_2569),
    .A2(n_1680),
    .B(n_1979),
    .Y(n_3771));
 OAI21xp33_ASAP7_75t_R g216466 (.A1(n_2231),
    .A2(n_1429),
    .B(n_1966),
    .Y(n_3770));
 OAI21xp33_ASAP7_75t_R g216467 (.A1(n_2304),
    .A2(n_1647),
    .B(n_2264),
    .Y(n_3769));
 NAND2xp33_ASAP7_75t_R g216468 (.A(n_2239),
    .B(n_3195),
    .Y(n_3768));
 OAI21xp33_ASAP7_75t_R g216469 (.A1(n_1496),
    .A2(n_2587),
    .B(n_1553),
    .Y(n_3767));
 OAI21xp33_ASAP7_75t_R g216470 (.A1(n_1611),
    .A2(n_2419),
    .B(sa00[0]),
    .Y(n_3766));
 AO21x1_ASAP7_75t_SL g216471 (.A1(sa11[3]),
    .A2(n_2227),
    .B(n_3206),
    .Y(n_3765));
 OAI21xp33_ASAP7_75t_R g216472 (.A1(n_8178),
    .A2(n_2437),
    .B(n_2346),
    .Y(n_3764));
 OAI21xp33_ASAP7_75t_R g216473 (.A1(n_1967),
    .A2(n_2457),
    .B(n_2338),
    .Y(n_3763));
 OA21x2_ASAP7_75t_R g216474 (.A1(n_8210),
    .A2(n_2438),
    .B(n_2380),
    .Y(n_3762));
 AOI21xp33_ASAP7_75t_R g216475 (.A1(n_2442),
    .A2(sa01[3]),
    .B(n_2342),
    .Y(n_3761));
 OAI21xp33_ASAP7_75t_R g216476 (.A1(n_2571),
    .A2(n_2061),
    .B(n_1540),
    .Y(n_3760));
 AOI21xp33_ASAP7_75t_R g216477 (.A1(n_2450),
    .A2(n_1519),
    .B(n_2373),
    .Y(n_3759));
 OA21x2_ASAP7_75t_R g216478 (.A1(n_1979),
    .A2(n_2484),
    .B(n_2382),
    .Y(n_3758));
 OA21x2_ASAP7_75t_R g216479 (.A1(n_1975),
    .A2(n_2476),
    .B(n_2377),
    .Y(n_3757));
 OA21x2_ASAP7_75t_R g216480 (.A1(n_1867),
    .A2(n_2453),
    .B(n_2379),
    .Y(n_3756));
 AOI21xp33_ASAP7_75t_R g216481 (.A1(sa22[3]),
    .A2(n_2440),
    .B(n_2336),
    .Y(n_3755));
 AOI21xp5_ASAP7_75t_L g216482 (.A1(n_1975),
    .A2(n_1502),
    .B(n_3517),
    .Y(n_3754));
 NOR3xp33_ASAP7_75t_L g216483 (.A(n_3255),
    .B(n_2546),
    .C(n_1343),
    .Y(n_3753));
 AOI21xp33_ASAP7_75t_R g216484 (.A1(n_1689),
    .A2(n_1534),
    .B(n_1558),
    .Y(n_3752));
 NOR3xp33_ASAP7_75t_R g216485 (.A(n_2797),
    .B(n_2580),
    .C(sa03[3]),
    .Y(n_3751));
 OAI21xp33_ASAP7_75t_R g216486 (.A1(sa10[7]),
    .A2(n_2594),
    .B(n_2394),
    .Y(n_3750));
 OAI21xp33_ASAP7_75t_R g216487 (.A1(n_1536),
    .A2(n_2548),
    .B(n_2397),
    .Y(n_3749));
 AO21x1_ASAP7_75t_R g216488 (.A1(n_2729),
    .A2(n_1689),
    .B(n_1496),
    .Y(n_3748));
 OAI21xp33_ASAP7_75t_R g216489 (.A1(n_1491),
    .A2(n_2546),
    .B(n_1566),
    .Y(n_3747));
 OAI21xp33_ASAP7_75t_R g216490 (.A1(n_1483),
    .A2(n_2590),
    .B(n_1653),
    .Y(n_3746));
 OAI21xp33_ASAP7_75t_R g216491 (.A1(n_1525),
    .A2(n_2560),
    .B(n_1645),
    .Y(n_3745));
 AOI21xp33_ASAP7_75t_R g216492 (.A1(n_2543),
    .A2(n_2019),
    .B(n_8691),
    .Y(n_3744));
 AOI21xp33_ASAP7_75t_L g216493 (.A1(n_2551),
    .A2(n_1485),
    .B(n_1639),
    .Y(n_3743));
 OAI21xp33_ASAP7_75t_R g216494 (.A1(sa02[7]),
    .A2(n_2558),
    .B(n_1422),
    .Y(n_3742));
 OAI21xp33_ASAP7_75t_R g216495 (.A1(sa13[7]),
    .A2(n_2550),
    .B(n_1436),
    .Y(n_3741));
 AOI21xp33_ASAP7_75t_R g216496 (.A1(n_2521),
    .A2(n_1982),
    .B(n_2399),
    .Y(n_3740));
 NOR3xp33_ASAP7_75t_R g216497 (.A(n_2856),
    .B(n_2560),
    .C(n_1984),
    .Y(n_3739));
 OAI21xp33_ASAP7_75t_R g216498 (.A1(n_2128),
    .A2(n_2434),
    .B(n_8208),
    .Y(n_3738));
 NAND2xp5_ASAP7_75t_L g216499 (.A(n_2215),
    .B(n_2777),
    .Y(n_4206));
 NAND2xp33_ASAP7_75t_R g216500 (.A(n_2882),
    .B(n_2902),
    .Y(n_4205));
 NAND2xp5_ASAP7_75t_R g216501 (.A(n_2042),
    .B(n_3056),
    .Y(n_4204));
 AOI21xp5_ASAP7_75t_R g216502 (.A1(n_2505),
    .A2(n_2525),
    .B(n_1665),
    .Y(n_4203));
 AOI21xp5_ASAP7_75t_R g216503 (.A1(n_2531),
    .A2(n_2568),
    .B(n_1635),
    .Y(n_4201));
 OR2x2_ASAP7_75t_SL g216504 (.A(n_2045),
    .B(n_3023),
    .Y(n_4200));
 AOI21xp33_ASAP7_75t_R g216505 (.A1(n_2503),
    .A2(n_2136),
    .B(n_2393),
    .Y(n_4199));
 NAND2xp5_ASAP7_75t_L g216506 (.A(n_3406),
    .B(n_1728),
    .Y(n_3737));
 NAND2xp33_ASAP7_75t_R g216507 (.A(n_2439),
    .B(n_3334),
    .Y(n_4197));
 NAND2xp5_ASAP7_75t_L g216508 (.A(n_2875),
    .B(n_2136),
    .Y(n_4196));
 NOR2xp67_ASAP7_75t_L g216509 (.A(n_3438),
    .B(n_3424),
    .Y(n_4195));
 NAND2xp5_ASAP7_75t_L g216510 (.A(n_2054),
    .B(n_2997),
    .Y(n_4194));
 NOR2xp33_ASAP7_75t_L g216511 (.A(n_1676),
    .B(n_3311),
    .Y(n_4193));
 AOI21xp5_ASAP7_75t_R g216512 (.A1(n_2496),
    .A2(n_2122),
    .B(n_2399),
    .Y(n_4192));
 NOR2xp33_ASAP7_75t_L g216513 (.A(n_2057),
    .B(n_3041),
    .Y(n_4190));
 NAND2xp5_ASAP7_75t_L g216514 (.A(n_2875),
    .B(n_2914),
    .Y(n_4188));
 NOR2xp33_ASAP7_75t_L g216515 (.A(n_1599),
    .B(n_2884),
    .Y(n_4187));
 NAND2xp5_ASAP7_75t_R g216516 (.A(n_3432),
    .B(n_3419),
    .Y(n_4186));
 OAI21xp33_ASAP7_75t_R g216517 (.A1(n_2530),
    .A2(n_2538),
    .B(n_1569),
    .Y(n_4184));
 NAND2xp5_ASAP7_75t_R g216518 (.A(n_2082),
    .B(n_3423),
    .Y(n_4183));
 NOR2xp33_ASAP7_75t_R g216519 (.A(n_2053),
    .B(n_3423),
    .Y(n_4182));
 NAND2xp5_ASAP7_75t_R g216520 (.A(n_1542),
    .B(n_3003),
    .Y(n_4181));
 OAI21xp33_ASAP7_75t_R g216521 (.A1(n_1690),
    .A2(n_2584),
    .B(n_2431),
    .Y(n_4180));
 AND2x2_ASAP7_75t_L g216522 (.A(n_1559),
    .B(n_3076),
    .Y(n_4179));
 NAND2xp33_ASAP7_75t_SL g216523 (.A(n_3414),
    .B(n_2873),
    .Y(n_1774));
 OAI21xp33_ASAP7_75t_R g216524 (.A1(n_1593),
    .A2(n_2507),
    .B(n_1653),
    .Y(n_4178));
 AOI21xp5_ASAP7_75t_R g216525 (.A1(n_2509),
    .A2(n_2132),
    .B(n_8720),
    .Y(n_4177));
 NAND2xp5_ASAP7_75t_L g216526 (.A(n_2079),
    .B(n_3413),
    .Y(n_3736));
 NAND2xp5_ASAP7_75t_R g216527 (.A(n_2878),
    .B(n_2200),
    .Y(n_4175));
 NAND2xp5_ASAP7_75t_R g216528 (.A(n_2899),
    .B(n_2878),
    .Y(n_4173));
 AOI21xp33_ASAP7_75t_R g216529 (.A1(n_2556),
    .A2(n_2512),
    .B(n_1626),
    .Y(n_4171));
 NAND2xp5_ASAP7_75t_SL g216530 (.A(n_2462),
    .B(n_3308),
    .Y(n_4169));
 NAND2xp5_ASAP7_75t_R g216531 (.A(n_2394),
    .B(n_3260),
    .Y(n_4168));
 NOR2xp33_ASAP7_75t_L g216532 (.A(n_1749),
    .B(n_3421),
    .Y(n_4167));
 OAI21xp33_ASAP7_75t_R g216533 (.A1(n_2185),
    .A2(n_2511),
    .B(n_1554),
    .Y(n_4166));
 AOI21xp5_ASAP7_75t_R g216534 (.A1(n_2519),
    .A2(n_2561),
    .B(n_1656),
    .Y(n_4164));
 AOI21xp5_ASAP7_75t_R g216535 (.A1(n_2521),
    .A2(n_2496),
    .B(n_2434),
    .Y(n_4163));
 NOR2xp33_ASAP7_75t_R g216536 (.A(n_2198),
    .B(n_3275),
    .Y(n_4162));
 NOR2xp33_ASAP7_75t_SL g216537 (.A(n_2091),
    .B(n_3425),
    .Y(n_4160));
 NAND2xp5_ASAP7_75t_R g216538 (.A(n_1559),
    .B(n_3425),
    .Y(n_4158));
 OAI21xp33_ASAP7_75t_R g216539 (.A1(n_1599),
    .A2(n_2513),
    .B(n_1445),
    .Y(n_4157));
 NAND2xp33_ASAP7_75t_L g216540 (.A(n_2429),
    .B(n_3219),
    .Y(n_3735));
 NOR2xp33_ASAP7_75t_L g216541 (.A(n_2041),
    .B(n_3451),
    .Y(n_4156));
 NAND2xp5_ASAP7_75t_R g216542 (.A(n_2092),
    .B(n_3451),
    .Y(n_4155));
 OAI21xp5_ASAP7_75t_R g216543 (.A1(n_2134),
    .A2(n_2535),
    .B(n_1350),
    .Y(n_4154));
 OAI21xp5_ASAP7_75t_L g216544 (.A1(n_2154),
    .A2(n_1690),
    .B(n_1638),
    .Y(n_4152));
 OAI21xp5_ASAP7_75t_R g216545 (.A1(n_2148),
    .A2(n_2532),
    .B(n_1645),
    .Y(n_4151));
 NAND2xp33_ASAP7_75t_R g216546 (.A(n_2835),
    .B(n_1677),
    .Y(n_4150));
 OAI21xp5_ASAP7_75t_R g216547 (.A1(n_2113),
    .A2(n_2538),
    .B(n_1566),
    .Y(n_4149));
 NAND2xp33_ASAP7_75t_R g216548 (.A(n_2820),
    .B(n_1622),
    .Y(n_4147));
 NAND2xp5_ASAP7_75t_SL g216549 (.A(n_2037),
    .B(n_1730),
    .Y(n_1773));
 NOR2xp33_ASAP7_75t_R g216550 (.A(n_1593),
    .B(n_2879),
    .Y(n_4146));
 NAND2xp5_ASAP7_75t_R g216551 (.A(n_2882),
    .B(n_2107),
    .Y(n_4144));
 OAI21xp33_ASAP7_75t_R g216552 (.A1(n_2200),
    .A2(n_2415),
    .B(n_2931),
    .Y(n_4142));
 NOR2xp33_ASAP7_75t_R g216553 (.A(n_1747),
    .B(n_3244),
    .Y(n_4141));
 AOI21xp5_ASAP7_75t_L g216554 (.A1(n_2534),
    .A2(n_1600),
    .B(n_2396),
    .Y(n_4140));
 NAND2xp5_ASAP7_75t_R g216555 (.A(n_1606),
    .B(n_3270),
    .Y(n_4139));
 NOR2xp33_ASAP7_75t_SL g216556 (.A(n_2177),
    .B(n_1726),
    .Y(n_4138));
 OAI21xp33_ASAP7_75t_R g216557 (.A1(n_2210),
    .A2(n_2526),
    .B(n_2394),
    .Y(n_4137));
 NOR2xp33_ASAP7_75t_L g216558 (.A(n_2134),
    .B(n_2885),
    .Y(n_4136));
 NAND2xp5_ASAP7_75t_R g216559 (.A(n_2159),
    .B(n_3266),
    .Y(n_4135));
 OAI21xp33_ASAP7_75t_R g216560 (.A1(n_2586),
    .A2(n_2507),
    .B(n_2410),
    .Y(n_4134));
 NOR2xp33_ASAP7_75t_L g216561 (.A(n_2871),
    .B(n_3327),
    .Y(n_4132));
 NAND2xp33_ASAP7_75t_R g216562 (.A(n_2791),
    .B(n_2215),
    .Y(n_4130));
 NAND2xp5_ASAP7_75t_R g216563 (.A(n_2429),
    .B(n_2805),
    .Y(n_4129));
 NAND2xp5_ASAP7_75t_SL g216564 (.A(n_2167),
    .B(n_2782),
    .Y(n_4127));
 NOR2xp33_ASAP7_75t_R g216565 (.A(n_2066),
    .B(n_2797),
    .Y(n_4126));
 NOR2x1_ASAP7_75t_R g216566 (.A(n_3277),
    .B(n_3293),
    .Y(n_4125));
 NAND2xp5_ASAP7_75t_L g216567 (.A(n_3243),
    .B(n_8703),
    .Y(n_4124));
 NAND2xp5_ASAP7_75t_L g216568 (.A(n_2205),
    .B(n_2783),
    .Y(n_4122));
 NOR2xp67_ASAP7_75t_SL g216569 (.A(n_1637),
    .B(n_1714),
    .Y(n_4120));
 NOR2xp33_ASAP7_75t_SL g216570 (.A(n_1558),
    .B(n_2799),
    .Y(n_4119));
 OAI21xp33_ASAP7_75t_R g216571 (.A1(n_2510),
    .A2(n_2576),
    .B(n_2413),
    .Y(n_4118));
 NOR2xp33_ASAP7_75t_R g216572 (.A(n_2154),
    .B(n_2909),
    .Y(n_4117));
 NOR2xp33_ASAP7_75t_R g216573 (.A(n_2104),
    .B(n_3241),
    .Y(n_3734));
 AOI21xp5_ASAP7_75t_R g216574 (.A1(n_2503),
    .A2(n_2553),
    .B(n_2423),
    .Y(n_4116));
 NAND2xp33_ASAP7_75t_R g216575 (.A(n_2893),
    .B(n_2910),
    .Y(n_4115));
 NAND2xp5_ASAP7_75t_R g216576 (.A(n_3334),
    .B(n_3283),
    .Y(n_4114));
 NAND2xp5_ASAP7_75t_L g216577 (.A(n_2880),
    .B(n_2883),
    .Y(n_4112));
 NAND2xp33_ASAP7_75t_R g216578 (.A(n_3363),
    .B(n_3324),
    .Y(n_4111));
 NOR2xp67_ASAP7_75t_L g216579 (.A(n_1654),
    .B(n_2780),
    .Y(n_4109));
 NAND2xp5_ASAP7_75t_L g216580 (.A(n_2900),
    .B(n_2475),
    .Y(n_4107));
 AOI21xp5_ASAP7_75t_R g216581 (.A1(n_1689),
    .A2(n_2587),
    .B(n_2066),
    .Y(n_4106));
 NAND2xp5_ASAP7_75t_R g216582 (.A(n_2954),
    .B(n_1419),
    .Y(n_4105));
 NOR2xp33_ASAP7_75t_L g216583 (.A(n_2102),
    .B(n_2792),
    .Y(n_4104));
 NAND2xp5_ASAP7_75t_R g216584 (.A(n_3254),
    .B(n_1715),
    .Y(n_4103));
 NAND2xp33_ASAP7_75t_R g216585 (.A(n_3257),
    .B(n_3361),
    .Y(n_4102));
 NOR2xp33_ASAP7_75t_L g216586 (.A(n_3290),
    .B(n_3263),
    .Y(n_4101));
 NAND2xp5_ASAP7_75t_L g216587 (.A(n_1445),
    .B(n_2777),
    .Y(n_4099));
 NAND2xp5_ASAP7_75t_L g216588 (.A(n_2788),
    .B(n_1451),
    .Y(n_4098));
 NAND2xp5_ASAP7_75t_R g216589 (.A(n_1750),
    .B(n_1751),
    .Y(n_4096));
 NAND2xp5_ASAP7_75t_R g216590 (.A(n_1713),
    .B(n_2912),
    .Y(n_1772));
 NAND2xp5_ASAP7_75t_R g216591 (.A(n_1439),
    .B(n_3556),
    .Y(n_4094));
 NAND2xp33_ASAP7_75t_L g216592 (.A(n_2854),
    .B(n_2385),
    .Y(n_4093));
 NOR2xp33_ASAP7_75t_R g216593 (.A(n_2829),
    .B(n_2080),
    .Y(n_4091));
 NAND2xp33_ASAP7_75t_R g216594 (.A(n_1423),
    .B(n_3297),
    .Y(n_4090));
 NOR2xp33_ASAP7_75t_R g216595 (.A(n_2078),
    .B(n_2860),
    .Y(n_4089));
 NAND2xp33_ASAP7_75t_R g216596 (.A(n_2820),
    .B(n_2859),
    .Y(n_4088));
 NOR2xp33_ASAP7_75t_R g216597 (.A(n_1337),
    .B(n_3313),
    .Y(n_4087));
 NAND2xp5_ASAP7_75t_R g216598 (.A(n_2090),
    .B(n_1715),
    .Y(n_4085));
 NAND2xp5_ASAP7_75t_L g216599 (.A(n_2896),
    .B(n_2890),
    .Y(n_4083));
 NOR2xp33_ASAP7_75t_L g216600 (.A(n_2858),
    .B(n_2856),
    .Y(n_4081));
 NOR2xp33_ASAP7_75t_L g216601 (.A(n_1575),
    .B(n_2844),
    .Y(n_4080));
 NOR2xp67_ASAP7_75t_L g216602 (.A(n_2083),
    .B(n_2858),
    .Y(n_4079));
 NOR2xp67_ASAP7_75t_SL g216603 (.A(n_2148),
    .B(n_2904),
    .Y(n_4077));
 NAND2xp5_ASAP7_75t_R g216604 (.A(n_3541),
    .B(n_1549),
    .Y(n_4075));
 NAND2xp5_ASAP7_75t_L g216605 (.A(n_2831),
    .B(n_1589),
    .Y(n_4074));
 NAND2xp5_ASAP7_75t_R g216606 (.A(n_2823),
    .B(n_2851),
    .Y(n_4072));
 NAND2xp5_ASAP7_75t_R g216607 (.A(n_2837),
    .B(n_1570),
    .Y(n_4070));
 NAND2xp5_ASAP7_75t_L g216608 (.A(n_2820),
    .B(n_2873),
    .Y(n_4068));
 NAND2xp5_ASAP7_75t_R g216609 (.A(n_2089),
    .B(n_2847),
    .Y(n_4067));
 NAND2xp5_ASAP7_75t_R g216610 (.A(n_1577),
    .B(n_2849),
    .Y(n_4066));
 NOR2xp33_ASAP7_75t_L g216611 (.A(n_3605),
    .B(n_1548),
    .Y(n_4065));
 NAND2xp5_ASAP7_75t_R g216612 (.A(n_2865),
    .B(n_2819),
    .Y(n_4063));
 NOR2xp33_ASAP7_75t_L g216613 (.A(n_3372),
    .B(n_3428),
    .Y(n_4062));
 NOR2xp33_ASAP7_75t_L g216614 (.A(n_2497),
    .B(n_3333),
    .Y(n_4060));
 NAND2xp33_ASAP7_75t_L g216615 (.A(n_2903),
    .B(n_2888),
    .Y(n_4059));
 NAND2xp5_ASAP7_75t_L g216616 (.A(n_2816),
    .B(n_2475),
    .Y(n_4058));
 NOR2xp33_ASAP7_75t_L g216617 (.A(n_1658),
    .B(n_3269),
    .Y(n_4057));
 NAND2xp5_ASAP7_75t_L g216618 (.A(n_3281),
    .B(n_2440),
    .Y(n_3733));
 NAND2xp33_ASAP7_75t_R g216619 (.A(n_2469),
    .B(n_3387),
    .Y(n_4056));
 NOR2xp33_ASAP7_75t_R g216620 (.A(n_2043),
    .B(n_2872),
    .Y(n_4054));
 AND2x2_ASAP7_75t_L g216621 (.A(n_2067),
    .B(n_3034),
    .Y(n_4053));
 NAND2xp5_ASAP7_75t_R g216622 (.A(n_3265),
    .B(n_2469),
    .Y(n_4052));
 NAND2xp5_ASAP7_75t_R g216623 (.A(n_3287),
    .B(n_2448),
    .Y(n_3732));
 NOR2xp33_ASAP7_75t_R g216624 (.A(n_2908),
    .B(n_3269),
    .Y(n_4051));
 NOR2xp33_ASAP7_75t_L g216625 (.A(n_2915),
    .B(n_2885),
    .Y(n_4049));
 NOR2xp33_ASAP7_75t_R g216626 (.A(n_1604),
    .B(n_3248),
    .Y(n_4048));
 NAND2xp5_ASAP7_75t_R g216627 (.A(n_2907),
    .B(n_2805),
    .Y(n_4046));
 NAND2xp5_ASAP7_75t_R g216628 (.A(n_2895),
    .B(n_3415),
    .Y(n_4045));
 AND2x2_ASAP7_75t_L g216629 (.A(n_2823),
    .B(n_2869),
    .Y(n_4044));
 NOR2xp33_ASAP7_75t_R g216630 (.A(n_2868),
    .B(n_1714),
    .Y(n_4043));
 NOR2xp33_ASAP7_75t_SL g216631 (.A(n_2866),
    .B(n_2801),
    .Y(n_4042));
 OAI21xp33_ASAP7_75t_R g216632 (.A1(n_2539),
    .A2(n_2572),
    .B(n_2404),
    .Y(n_4041));
 NAND2xp5_ASAP7_75t_L g216633 (.A(n_1603),
    .B(n_3243),
    .Y(n_4039));
 NAND2xp33_ASAP7_75t_R g216634 (.A(n_2105),
    .B(n_1718),
    .Y(n_4038));
 NAND2xp5_ASAP7_75t_R g216635 (.A(n_1718),
    .B(n_2863),
    .Y(n_4037));
 NAND2xp5_ASAP7_75t_SL g216636 (.A(n_2863),
    .B(n_2452),
    .Y(n_1771));
 NOR2xp33_ASAP7_75t_R g216637 (.A(n_2453),
    .B(n_3270),
    .Y(n_4036));
 NOR2xp33_ASAP7_75t_L g216638 (.A(n_2120),
    .B(n_2786),
    .Y(n_4034));
 OAI21xp5_ASAP7_75t_L g216639 (.A1(n_2524),
    .A2(n_2535),
    .B(n_2425),
    .Y(n_4033));
 AOI21xp33_ASAP7_75t_R g216640 (.A1(n_2502),
    .A2(n_2534),
    .B(n_2428),
    .Y(n_4031));
 NOR2xp33_ASAP7_75t_R g216641 (.A(n_2879),
    .B(n_2906),
    .Y(n_4030));
 NAND2xp5_ASAP7_75t_L g216642 (.A(n_2436),
    .B(n_3329),
    .Y(n_4029));
 NOR2xp33_ASAP7_75t_R g216643 (.A(n_2437),
    .B(n_3273),
    .Y(n_4027));
 NOR2xp67_ASAP7_75t_SL g216644 (.A(n_1602),
    .B(n_3252),
    .Y(n_4026));
 NAND2xp5_ASAP7_75t_R g216645 (.A(n_2110),
    .B(n_3260),
    .Y(n_4025));
 NAND2xp5_ASAP7_75t_SL g216646 (.A(n_2450),
    .B(n_2914),
    .Y(n_4023));
 NOR2x1_ASAP7_75t_L g216647 (.A(n_1588),
    .B(n_2825),
    .Y(n_1770));
 NOR2xp33_ASAP7_75t_L g216648 (.A(n_3309),
    .B(n_2063),
    .Y(n_4022));
 NAND2xp5_ASAP7_75t_L g216649 (.A(n_2072),
    .B(n_2835),
    .Y(n_4020));
 NOR2xp33_ASAP7_75t_L g216650 (.A(n_2088),
    .B(n_3315),
    .Y(n_4018));
 NAND2xp5_ASAP7_75t_L g216651 (.A(n_1581),
    .B(n_2840),
    .Y(n_4016));
 NAND2xp5_ASAP7_75t_L g216652 (.A(n_1586),
    .B(n_3310),
    .Y(n_1769));
 AND2x2_ASAP7_75t_SL g216653 (.A(n_2084),
    .B(n_3306),
    .Y(n_4015));
 NAND2xp5_ASAP7_75t_L g216654 (.A(n_2090),
    .B(n_2845),
    .Y(n_4014));
 NAND2xp5_ASAP7_75t_L g216655 (.A(n_2079),
    .B(n_2854),
    .Y(n_4012));
 NOR2xp33_ASAP7_75t_SL g216656 (.A(n_1575),
    .B(n_2842),
    .Y(n_4011));
 NOR2xp33_ASAP7_75t_SL g216657 (.A(n_2081),
    .B(n_3279),
    .Y(n_4008));
 NAND2xp5_ASAP7_75t_L g216658 (.A(n_2075),
    .B(n_3302),
    .Y(n_4007));
 NOR2x1_ASAP7_75t_SL g216659 (.A(n_2486),
    .B(n_2889),
    .Y(n_4006));
 NOR2x1_ASAP7_75t_R g216660 (.A(n_1342),
    .B(n_3298),
    .Y(n_4005));
 AND2x2_ASAP7_75t_L g216661 (.A(n_2900),
    .B(n_2833),
    .Y(n_4003));
 NOR2x1_ASAP7_75t_SL g216662 (.A(n_2482),
    .B(n_2894),
    .Y(n_4000));
 NOR2xp33_ASAP7_75t_SL g216663 (.A(n_3395),
    .B(n_2797),
    .Y(n_3998));
 NOR2xp67_ASAP7_75t_L g216664 (.A(n_2206),
    .B(n_1729),
    .Y(n_3997));
 NOR2xp33_ASAP7_75t_SL g216665 (.A(n_2185),
    .B(n_2891),
    .Y(n_3996));
 NOR2xp33_ASAP7_75t_L g216666 (.A(n_3417),
    .B(n_2856),
    .Y(n_3994));
 NAND2xp5_ASAP7_75t_L g216667 (.A(n_3284),
    .B(n_3329),
    .Y(n_3992));
 NOR2xp33_ASAP7_75t_SL g216668 (.A(n_2170),
    .B(n_1714),
    .Y(n_3991));
 NAND2xp5_ASAP7_75t_SL g216669 (.A(n_2467),
    .B(n_2905),
    .Y(n_3988));
 NAND2x1_ASAP7_75t_L g216670 (.A(n_2473),
    .B(n_2902),
    .Y(n_3987));
 NAND2xp5_ASAP7_75t_R g216671 (.A(n_3419),
    .B(n_2439),
    .Y(n_3986));
 NAND2xp5_ASAP7_75t_SL g216672 (.A(n_1595),
    .B(n_2798),
    .Y(n_3984));
 NAND2xp5_ASAP7_75t_L g216673 (.A(n_3324),
    .B(n_3387),
    .Y(n_3982));
 NOR2xp33_ASAP7_75t_SL g216674 (.A(n_2482),
    .B(n_3394),
    .Y(n_3981));
 NAND2xp5_ASAP7_75t_L g216675 (.A(n_2899),
    .B(n_2483),
    .Y(n_3979));
 NOR2xp67_ASAP7_75t_L g216676 (.A(n_2474),
    .B(n_3379),
    .Y(n_3977));
 NAND2xp5_ASAP7_75t_R g216677 (.A(n_2873),
    .B(n_2477),
    .Y(n_3976));
 NOR2xp67_ASAP7_75t_L g216678 (.A(n_2443),
    .B(n_2852),
    .Y(n_3974));
 AND2x2_ASAP7_75t_SL g216679 (.A(n_2435),
    .B(n_3283),
    .Y(n_3972));
 NAND2xp5_ASAP7_75t_L g216680 (.A(n_2420),
    .B(n_3276),
    .Y(n_3971));
 NAND2xp5_ASAP7_75t_L g216681 (.A(n_2865),
    .B(n_2483),
    .Y(n_3968));
 NAND2xp5_ASAP7_75t_SL g216682 (.A(n_3365),
    .B(n_2467),
    .Y(n_3966));
 NAND2xp5_ASAP7_75t_L g216683 (.A(n_2192),
    .B(n_2779),
    .Y(n_3964));
 NAND2xp5_ASAP7_75t_L g216684 (.A(n_1569),
    .B(n_2783),
    .Y(n_3963));
 NAND2xp5_ASAP7_75t_SL g216685 (.A(n_2178),
    .B(n_3258),
    .Y(n_3961));
 NAND2xp33_ASAP7_75t_R g216686 (.A(n_2401),
    .B(n_2819),
    .Y(n_3959));
 NOR2x1_ASAP7_75t_L g216687 (.A(n_3394),
    .B(n_3263),
    .Y(n_3957));
 AND2x2_ASAP7_75t_SL g216688 (.A(n_2385),
    .B(n_2789),
    .Y(n_3956));
 NAND2xp33_ASAP7_75t_R g216689 (.A(n_2427),
    .B(n_2782),
    .Y(n_3954));
 NOR2xp33_ASAP7_75t_R g216690 (.A(n_1632),
    .B(n_3241),
    .Y(n_3952));
 NOR2x1_ASAP7_75t_R g216691 (.A(n_2088),
    .B(n_2949),
    .Y(n_3951));
 NAND2xp5_ASAP7_75t_R g216692 (.A(n_2103),
    .B(n_2807),
    .Y(n_3949));
 NAND2xp5_ASAP7_75t_R g216693 (.A(n_3292),
    .B(n_2450),
    .Y(n_3948));
 NAND2xp5_ASAP7_75t_R g216694 (.A(n_2431),
    .B(n_2823),
    .Y(n_3946));
 NAND2xp5_ASAP7_75t_L g216695 (.A(n_2072),
    .B(n_3064),
    .Y(n_3945));
 NAND2x1_ASAP7_75t_L g216696 (.A(n_2095),
    .B(n_2805),
    .Y(n_3944));
 NAND2xp5_ASAP7_75t_SL g216697 (.A(n_2092),
    .B(n_2973),
    .Y(n_3942));
 AND2x2_ASAP7_75t_L g216698 (.A(n_2079),
    .B(n_3035),
    .Y(n_3941));
 AND2x2_ASAP7_75t_R g216699 (.A(n_1664),
    .B(n_3273),
    .Y(n_3940));
 NOR2xp67_ASAP7_75t_L g216700 (.A(n_1342),
    .B(n_2965),
    .Y(n_3938));
 NAND2xp5_ASAP7_75t_SL g216701 (.A(n_3361),
    .B(n_3253),
    .Y(n_3936));
 OR2x2_ASAP7_75t_R g216702 (.A(n_2946),
    .B(n_1580),
    .Y(n_3935));
 NAND2xp5_ASAP7_75t_L g216703 (.A(n_1589),
    .B(n_2959),
    .Y(n_3933));
 NAND2xp5_ASAP7_75t_L g216704 (.A(n_2075),
    .B(n_3039),
    .Y(n_3931));
 NOR2xp33_ASAP7_75t_SL g216705 (.A(n_1344),
    .B(n_3014),
    .Y(n_3930));
 NAND2xp5_ASAP7_75t_L g216706 (.A(n_3274),
    .B(n_2414),
    .Y(n_3928));
 NAND2xp5_ASAP7_75t_L g216707 (.A(n_2870),
    .B(n_3300),
    .Y(n_3927));
 AND2x2_ASAP7_75t_L g216708 (.A(n_2420),
    .B(n_1727),
    .Y(n_3926));
 NAND2xp5_ASAP7_75t_SL g216709 (.A(n_1585),
    .B(n_1725),
    .Y(n_3925));
 NOR2xp33_ASAP7_75t_L g216710 (.A(n_2063),
    .B(n_2999),
    .Y(n_3924));
 NAND2xp5_ASAP7_75t_L g216711 (.A(n_2084),
    .B(n_2955),
    .Y(n_3922));
 NOR2xp67_ASAP7_75t_L g216712 (.A(n_2081),
    .B(n_2982),
    .Y(n_3921));
 NOR3xp33_ASAP7_75t_L g216713 (.A(n_2249),
    .B(n_2091),
    .C(n_2495),
    .Y(n_1768));
 NAND2xp5_ASAP7_75t_R g216714 (.A(n_2788),
    .B(n_2101),
    .Y(n_1767));
 NOR2x1_ASAP7_75t_L g216715 (.A(n_3364),
    .B(n_3303),
    .Y(n_3919));
 AND2x2_ASAP7_75t_L g216716 (.A(n_2065),
    .B(n_1732),
    .Y(n_3918));
 AND2x2_ASAP7_75t_SL g216717 (.A(n_2435),
    .B(n_2802),
    .Y(n_1766));
 NAND2xp5_ASAP7_75t_L g216718 (.A(n_2431),
    .B(n_2811),
    .Y(n_3916));
 NAND2xp5_ASAP7_75t_L g216719 (.A(n_2425),
    .B(n_2817),
    .Y(n_3914));
 OAI21xp5_ASAP7_75t_L g216720 (.A1(sa23[1]),
    .A2(n_2470),
    .B(n_3324),
    .Y(n_3912));
 NOR2x1_ASAP7_75t_L g216721 (.A(n_3295),
    .B(n_2862),
    .Y(n_3911));
 NAND2xp5_ASAP7_75t_L g216722 (.A(n_2916),
    .B(n_2835),
    .Y(n_3909));
 OAI21xp5_ASAP7_75t_R g216723 (.A1(n_1522),
    .A2(n_2476),
    .B(n_2833),
    .Y(n_3906));
 NAND2xp5_ASAP7_75t_R g216724 (.A(n_2401),
    .B(n_2793),
    .Y(n_3905));
 AOI21xp5_ASAP7_75t_L g216725 (.A1(n_2477),
    .A2(n_1475),
    .B(n_2821),
    .Y(n_3904));
 NAND2xp5_ASAP7_75t_R g216726 (.A(n_1733),
    .B(n_1751),
    .Y(n_3902));
 AOI21xp5_ASAP7_75t_SL g216727 (.A1(n_2452),
    .A2(n_1862),
    .B(n_3327),
    .Y(n_3900));
 OAI21xp5_ASAP7_75t_L g216728 (.A1(sa12[1]),
    .A2(n_2482),
    .B(n_3262),
    .Y(n_1765));
 OAI21xp5_ASAP7_75t_L g216729 (.A1(sa10[1]),
    .A2(n_2437),
    .B(n_3284),
    .Y(n_3898));
 NOR2x1_ASAP7_75t_SL g216730 (.A(n_2853),
    .B(n_1720),
    .Y(n_3897));
 AOI21xp5_ASAP7_75t_SL g216731 (.A1(n_2485),
    .A2(n_1904),
    .B(n_2856),
    .Y(n_3895));
 OA21x2_ASAP7_75t_R g216732 (.A1(n_1470),
    .A2(n_2441),
    .B(n_3257),
    .Y(n_3894));
 AOI21xp5_ASAP7_75t_L g216733 (.A1(n_2448),
    .A2(n_1995),
    .B(n_3255),
    .Y(n_3892));
 NOR2xp33_ASAP7_75t_SL g216734 (.A(n_3288),
    .B(n_3372),
    .Y(n_3890));
 NOR2x1_ASAP7_75t_SL g216735 (.A(n_2846),
    .B(n_1749),
    .Y(n_3888));
 OAI21xp5_ASAP7_75t_L g216736 (.A1(sa02[1]),
    .A2(n_2438),
    .B(n_3283),
    .Y(n_3887));
 NOR2x1_ASAP7_75t_L g216737 (.A(n_2898),
    .B(n_2839),
    .Y(n_3885));
 NOR2xp67_ASAP7_75t_L g216738 (.A(n_3230),
    .B(n_2797),
    .Y(n_1763));
 AND2x2_ASAP7_75t_L g216739 (.A(n_3419),
    .B(n_3302),
    .Y(n_3884));
 NOR2x1p5_ASAP7_75t_SL g216740 (.A(n_3438),
    .B(n_3279),
    .Y(n_3882));
 NOR2x1_ASAP7_75t_SL g216741 (.A(n_2842),
    .B(n_2901),
    .Y(n_3880));
 AOI21xp5_ASAP7_75t_L g216742 (.A1(n_2483),
    .A2(n_8204),
    .B(n_2818),
    .Y(n_3879));
 OAI21xp5_ASAP7_75t_L g216743 (.A1(n_1473),
    .A2(n_2451),
    .B(n_3276),
    .Y(n_3877));
 OAI21xp5_ASAP7_75t_SL g216744 (.A1(n_1479),
    .A2(n_2474),
    .B(n_3268),
    .Y(n_3876));
 NOR2x1_ASAP7_75t_SL g216745 (.A(n_3224),
    .B(n_3245),
    .Y(n_3875));
 NAND2xp5_ASAP7_75t_L g216746 (.A(n_2410),
    .B(n_1711),
    .Y(n_3874));
 OAI21xp5_ASAP7_75t_L g216747 (.A1(n_1492),
    .A2(n_2443),
    .B(n_2823),
    .Y(n_3872));
 AND2x2_ASAP7_75t_SL g216748 (.A(n_2469),
    .B(n_1751),
    .Y(n_3870));
 OAI21xp5_ASAP7_75t_SL g216749 (.A1(n_8204),
    .A2(n_2102),
    .B(n_3344),
    .Y(n_3868));
 NOR2xp33_ASAP7_75t_L g216750 (.A(n_2897),
    .B(n_3315),
    .Y(n_3866));
 NOR2x1_ASAP7_75t_SL g216751 (.A(n_3228),
    .B(n_2908),
    .Y(n_3864));
 NOR2x1_ASAP7_75t_L g216752 (.A(n_2825),
    .B(n_2892),
    .Y(n_3863));
 NOR2x1_ASAP7_75t_SL g216753 (.A(n_3231),
    .B(n_3476),
    .Y(n_3861));
 NAND2x1_ASAP7_75t_SL g216754 (.A(n_1657),
    .B(n_2814),
    .Y(n_3860));
 NAND2xp5_ASAP7_75t_SL g216755 (.A(n_2475),
    .B(n_2916),
    .Y(n_3858));
 NAND2x1_ASAP7_75t_SL g216756 (.A(n_2442),
    .B(n_2893),
    .Y(n_3856));
 NAND2x1_ASAP7_75t_SL g216757 (.A(n_2448),
    .B(n_3427),
    .Y(n_3854));
 NAND2x1_ASAP7_75t_SL g216758 (.A(n_3437),
    .B(n_2440),
    .Y(n_1761));
 OR2x2_ASAP7_75t_SL g216759 (.A(n_2478),
    .B(n_1720),
    .Y(n_3851));
 NOR2x1_ASAP7_75t_SL g216760 (.A(n_2457),
    .B(n_2897),
    .Y(n_3848));
 NAND2xp5_ASAP7_75t_SL g216761 (.A(n_1705),
    .B(n_2740),
    .Y(n_3847));
 AND2x2_ASAP7_75t_SL g216762 (.A(n_1701),
    .B(n_2739),
    .Y(n_3845));
 INVxp67_ASAP7_75t_L g216763 (.A(n_3729),
    .Y(n_3730));
 INVxp33_ASAP7_75t_R g216764 (.A(n_3725),
    .Y(n_3726));
 INVxp33_ASAP7_75t_R g216765 (.A(n_3722),
    .Y(n_3723));
 INVxp67_ASAP7_75t_R g216766 (.A(n_3720),
    .Y(n_3721));
 INVxp67_ASAP7_75t_R g216767 (.A(n_3717),
    .Y(n_3718));
 INVxp67_ASAP7_75t_R g216768 (.A(n_3715),
    .Y(n_3716));
 INVxp33_ASAP7_75t_R g216769 (.A(n_3710),
    .Y(n_3711));
 INVxp67_ASAP7_75t_R g216770 (.A(n_3708),
    .Y(n_3709));
 INVxp33_ASAP7_75t_R g216771 (.A(n_3706),
    .Y(n_3707));
 INVxp33_ASAP7_75t_R g216772 (.A(n_3704),
    .Y(n_3705));
 INVxp33_ASAP7_75t_R g216773 (.A(n_3700),
    .Y(n_3701));
 INVxp33_ASAP7_75t_R g216775 (.A(n_3695),
    .Y(n_3696));
 INVxp33_ASAP7_75t_R g216776 (.A(n_3693),
    .Y(n_3694));
 INVxp67_ASAP7_75t_SL g216777 (.A(n_3682),
    .Y(n_3683));
 INVxp33_ASAP7_75t_R g216778 (.A(n_3676),
    .Y(n_3677));
 INVxp33_ASAP7_75t_R g216779 (.A(n_3671),
    .Y(n_3672));
 INVxp33_ASAP7_75t_R g216780 (.A(n_3669),
    .Y(n_3670));
 INVxp67_ASAP7_75t_L g216781 (.A(n_3665),
    .Y(n_3666));
 INVxp33_ASAP7_75t_R g216783 (.A(n_3651),
    .Y(n_3652));
 INVxp67_ASAP7_75t_R g216784 (.A(n_3648),
    .Y(n_3649));
 INVxp33_ASAP7_75t_R g216785 (.A(n_3644),
    .Y(n_3645));
 INVxp33_ASAP7_75t_R g216786 (.A(n_3642),
    .Y(n_3643));
 INVxp33_ASAP7_75t_R g216787 (.A(n_3639),
    .Y(n_3640));
 INVxp33_ASAP7_75t_R g216788 (.A(n_3633),
    .Y(n_3634));
 INVxp33_ASAP7_75t_R g216789 (.A(n_3625),
    .Y(n_3626));
 INVxp33_ASAP7_75t_R g216790 (.A(n_3623),
    .Y(n_3624));
 INVxp33_ASAP7_75t_R g216792 (.A(n_3614),
    .Y(n_3615));
 INVxp33_ASAP7_75t_R g216793 (.A(n_3609),
    .Y(n_3610));
 INVxp33_ASAP7_75t_R g216794 (.A(n_3607),
    .Y(n_3608));
 INVxp33_ASAP7_75t_R g216795 (.A(n_3603),
    .Y(n_3604));
 INVxp33_ASAP7_75t_R g216796 (.A(n_3600),
    .Y(n_3601));
 INVxp67_ASAP7_75t_L g216797 (.A(n_3597),
    .Y(n_3598));
 INVx1_ASAP7_75t_SL g216798 (.A(n_3591),
    .Y(n_3592));
 INVxp67_ASAP7_75t_L g216799 (.A(n_3587),
    .Y(n_3588));
 INVxp33_ASAP7_75t_R g216800 (.A(n_3585),
    .Y(n_3584));
 INVxp33_ASAP7_75t_R g216801 (.A(n_3582),
    .Y(n_3583));
 INVx1_ASAP7_75t_L g216802 (.A(n_3580),
    .Y(n_3581));
 INVxp33_ASAP7_75t_R g216806 (.A(n_3575),
    .Y(n_3576));
 HB1xp67_ASAP7_75t_L g216807 (.A(n_3573),
    .Y(n_3574));
 INVxp67_ASAP7_75t_R g216808 (.A(n_3572),
    .Y(n_3571));
 INVxp33_ASAP7_75t_R g216809 (.A(n_3569),
    .Y(n_3570));
 INVxp33_ASAP7_75t_R g216811 (.A(n_3566),
    .Y(n_3567));
 INVxp67_ASAP7_75t_R g216812 (.A(n_3565),
    .Y(n_3564));
 INVxp33_ASAP7_75t_R g216813 (.A(n_3562),
    .Y(n_3563));
 INVxp67_ASAP7_75t_R g216814 (.A(n_3558),
    .Y(n_3559));
 INVxp33_ASAP7_75t_R g216815 (.A(n_3552),
    .Y(n_3553));
 INVxp67_ASAP7_75t_R g216816 (.A(n_3550),
    .Y(n_3549));
 INVxp33_ASAP7_75t_R g216817 (.A(n_3543),
    .Y(n_3544));
 INVxp33_ASAP7_75t_R g216818 (.A(n_3539),
    .Y(n_3540));
 INVxp67_ASAP7_75t_R g216819 (.A(n_3538),
    .Y(n_3537));
 INVx1_ASAP7_75t_L g216820 (.A(n_3534),
    .Y(n_3535));
 INVx1_ASAP7_75t_R g216821 (.A(n_3530),
    .Y(n_3531));
 INVxp67_ASAP7_75t_R g216823 (.A(n_3528),
    .Y(n_3529));
 INVx1_ASAP7_75t_L g216824 (.A(n_3524),
    .Y(n_3525));
 INVxp67_ASAP7_75t_L g216825 (.A(n_3523),
    .Y(n_3522));
 INVx1_ASAP7_75t_R g216826 (.A(n_3521),
    .Y(n_3520));
 INVxp67_ASAP7_75t_R g216827 (.A(n_3517),
    .Y(n_3518));
 INVxp67_ASAP7_75t_R g216828 (.A(n_3516),
    .Y(n_3515));
 INVx1_ASAP7_75t_R g216829 (.A(n_3511),
    .Y(n_3512));
 INVxp67_ASAP7_75t_R g216830 (.A(n_3509),
    .Y(n_3510));
 INVxp33_ASAP7_75t_R g216831 (.A(n_3508),
    .Y(n_3507));
 INVxp67_ASAP7_75t_R g216833 (.A(n_3506),
    .Y(n_3505));
 INVxp67_ASAP7_75t_R g216834 (.A(n_3502),
    .Y(n_3503));
 INVxp67_ASAP7_75t_SL g216835 (.A(n_3501),
    .Y(n_3500));
 INVx1_ASAP7_75t_SL g216836 (.A(n_3499),
    .Y(n_3498));
 INVx1_ASAP7_75t_L g216838 (.A(n_1753),
    .Y(n_3496));
 INVxp67_ASAP7_75t_SL g216839 (.A(n_3495),
    .Y(n_3494));
 INVx1_ASAP7_75t_L g216840 (.A(n_3486),
    .Y(n_3487));
 INVxp33_ASAP7_75t_R g216841 (.A(n_3485),
    .Y(n_3484));
 INVxp33_ASAP7_75t_R g216842 (.A(n_3483),
    .Y(n_3482));
 INVxp67_ASAP7_75t_L g216843 (.A(n_3480),
    .Y(n_3481));
 INVxp67_ASAP7_75t_R g216844 (.A(n_3479),
    .Y(n_3478));
 INVxp67_ASAP7_75t_R g216845 (.A(n_3474),
    .Y(n_3475));
 INVxp67_ASAP7_75t_R g216846 (.A(n_3473),
    .Y(n_3472));
 INVxp67_ASAP7_75t_R g216847 (.A(n_3470),
    .Y(n_3471));
 INVxp33_ASAP7_75t_R g216848 (.A(n_3469),
    .Y(n_3468));
 INVxp33_ASAP7_75t_R g216849 (.A(n_3467),
    .Y(n_3466));
 INVxp67_ASAP7_75t_R g216850 (.A(n_3465),
    .Y(n_3464));
 INVxp33_ASAP7_75t_R g216851 (.A(n_3461),
    .Y(n_3460));
 INVxp67_ASAP7_75t_L g216852 (.A(n_3459),
    .Y(n_3458));
 INVxp33_ASAP7_75t_R g216853 (.A(n_3457),
    .Y(n_3456));
 INVx1_ASAP7_75t_L g216854 (.A(n_3451),
    .Y(n_3450));
 INVx1_ASAP7_75t_L g216855 (.A(n_3449),
    .Y(n_3448));
 INVxp67_ASAP7_75t_R g216856 (.A(n_3447),
    .Y(n_3446));
 INVxp67_ASAP7_75t_R g216857 (.A(n_3445),
    .Y(n_3444));
 INVxp67_ASAP7_75t_SL g216858 (.A(n_3443),
    .Y(n_3442));
 INVxp67_ASAP7_75t_R g216859 (.A(n_1752),
    .Y(n_3441));
 INVx1_ASAP7_75t_R g216861 (.A(n_3440),
    .Y(n_3439));
 INVx2_ASAP7_75t_SL g216862 (.A(n_3437),
    .Y(n_3438));
 INVxp33_ASAP7_75t_R g216863 (.A(n_1751),
    .Y(n_3436));
 INVx1_ASAP7_75t_R g216866 (.A(n_3435),
    .Y(n_3434));
 INVxp33_ASAP7_75t_R g216868 (.A(n_3432),
    .Y(n_3433));
 INVxp67_ASAP7_75t_R g216869 (.A(n_3431),
    .Y(n_3430));
 INVxp67_ASAP7_75t_R g216870 (.A(n_3429),
    .Y(n_3428));
 INVx2_ASAP7_75t_L g216872 (.A(n_3427),
    .Y(n_1749));
 INVxp33_ASAP7_75t_R g216874 (.A(n_3423),
    .Y(n_3422));
 INVx1_ASAP7_75t_R g216875 (.A(n_3421),
    .Y(n_3420));
 INVx2_ASAP7_75t_SL g216876 (.A(n_3419),
    .Y(n_3418));
 INVx1_ASAP7_75t_SL g216877 (.A(n_3416),
    .Y(n_3417));
 INVxp67_ASAP7_75t_L g216878 (.A(n_3414),
    .Y(n_3413));
 INVxp67_ASAP7_75t_R g216880 (.A(n_1748),
    .Y(n_3412));
 INVxp67_ASAP7_75t_R g216881 (.A(n_3411),
    .Y(n_3410));
 INVxp67_ASAP7_75t_R g216882 (.A(n_3409),
    .Y(n_3408));
 INVx2_ASAP7_75t_L g216883 (.A(n_3407),
    .Y(n_3406));
 INVxp67_ASAP7_75t_R g216884 (.A(n_3405),
    .Y(n_3404));
 INVx1_ASAP7_75t_L g216888 (.A(n_1746),
    .Y(n_1747));
 INVx1_ASAP7_75t_R g216889 (.A(n_3402),
    .Y(n_3403));
 INVx1_ASAP7_75t_L g216890 (.A(n_3401),
    .Y(n_3400));
 INVxp33_ASAP7_75t_R g216891 (.A(n_3399),
    .Y(n_3398));
 INVxp33_ASAP7_75t_R g216895 (.A(n_1745),
    .Y(n_1744));
 INVxp67_ASAP7_75t_L g216896 (.A(n_3396),
    .Y(n_3395));
 INVx1_ASAP7_75t_L g216897 (.A(n_3394),
    .Y(n_3393));
 INVxp33_ASAP7_75t_R g216898 (.A(n_3392),
    .Y(n_3391));
 INVxp67_ASAP7_75t_R g216899 (.A(n_3390),
    .Y(n_3389));
 INVxp33_ASAP7_75t_R g216900 (.A(n_3387),
    .Y(n_3388));
 INVx1_ASAP7_75t_L g216901 (.A(n_3386),
    .Y(n_3385));
 INVx1_ASAP7_75t_L g216902 (.A(n_3384),
    .Y(n_3383));
 INVx1_ASAP7_75t_R g216903 (.A(n_3382),
    .Y(n_3381));
 INVxp67_ASAP7_75t_L g216906 (.A(n_1743),
    .Y(n_1742));
 INVx1_ASAP7_75t_L g216907 (.A(n_3380),
    .Y(n_3379));
 INVxp67_ASAP7_75t_R g216908 (.A(n_3378),
    .Y(n_3377));
 INVxp33_ASAP7_75t_R g216909 (.A(n_3376),
    .Y(n_3375));
 INVx1_ASAP7_75t_L g216910 (.A(n_3374),
    .Y(n_3373));
 INVxp33_ASAP7_75t_R g216911 (.A(n_3372),
    .Y(n_3371));
 INVxp67_ASAP7_75t_L g216912 (.A(n_3370),
    .Y(n_3369));
 INVxp67_ASAP7_75t_SL g216913 (.A(n_3368),
    .Y(n_3367));
 INVxp67_ASAP7_75t_L g216914 (.A(n_3366),
    .Y(n_3365));
 INVxp67_ASAP7_75t_R g216915 (.A(n_3364),
    .Y(n_3363));
 INVx1_ASAP7_75t_R g216917 (.A(n_3360),
    .Y(n_3359));
 INVxp67_ASAP7_75t_R g216918 (.A(n_1741),
    .Y(n_3357));
 INVx1_ASAP7_75t_L g216925 (.A(n_3355),
    .Y(n_3354));
 INVxp67_ASAP7_75t_R g216926 (.A(n_3353),
    .Y(n_3352));
 INVxp33_ASAP7_75t_R g216927 (.A(n_3351),
    .Y(n_3350));
 INVxp67_ASAP7_75t_SL g216929 (.A(n_1738),
    .Y(n_1739));
 INVx1_ASAP7_75t_L g216932 (.A(n_3349),
    .Y(n_3348));
 INVxp33_ASAP7_75t_R g216933 (.A(n_3347),
    .Y(n_3346));
 INVx1_ASAP7_75t_L g216934 (.A(n_3344),
    .Y(n_3345));
 INVxp67_ASAP7_75t_L g216935 (.A(n_3341),
    .Y(n_3342));
 HB1xp67_ASAP7_75t_SL g216937 (.A(n_3340),
    .Y(n_3341));
 INVxp67_ASAP7_75t_L g216940 (.A(n_3338),
    .Y(n_1737));
 INVxp67_ASAP7_75t_R g216942 (.A(n_1736),
    .Y(n_3337));
 INVxp33_ASAP7_75t_R g216943 (.A(n_3336),
    .Y(n_3335));
 INVx1_ASAP7_75t_L g216944 (.A(n_3334),
    .Y(n_3333));
 INVxp33_ASAP7_75t_R g216945 (.A(n_3330),
    .Y(n_3331));
 BUFx2_ASAP7_75t_SL g216946 (.A(n_3332),
    .Y(n_3330));
 INVxp33_ASAP7_75t_R g216947 (.A(n_3329),
    .Y(n_3328));
 INVx1_ASAP7_75t_L g216948 (.A(n_3327),
    .Y(n_3326));
 INVx2_ASAP7_75t_SL g216949 (.A(n_1735),
    .Y(n_3325));
 INVxp67_ASAP7_75t_L g216953 (.A(n_3324),
    .Y(n_3323));
 INVx1_ASAP7_75t_R g216954 (.A(n_3322),
    .Y(n_3321));
 INVx1_ASAP7_75t_L g216955 (.A(n_3320),
    .Y(n_3319));
 INVx1_ASAP7_75t_L g216958 (.A(n_3317),
    .Y(n_1734));
 INVx2_ASAP7_75t_SL g216959 (.A(n_3316),
    .Y(n_3317));
 INVx1_ASAP7_75t_SL g216961 (.A(n_3315),
    .Y(n_3314));
 INVx1_ASAP7_75t_L g216962 (.A(n_3313),
    .Y(n_3312));
 INVx2_ASAP7_75t_SL g216963 (.A(n_3311),
    .Y(n_3310));
 INVx2_ASAP7_75t_L g216964 (.A(n_3309),
    .Y(n_3308));
 INVx2_ASAP7_75t_SL g216965 (.A(n_3307),
    .Y(n_3306));
 INVx1_ASAP7_75t_SL g216967 (.A(n_1733),
    .Y(n_3305));
 INVx1_ASAP7_75t_L g216969 (.A(n_3304),
    .Y(n_3303));
 INVx1_ASAP7_75t_SL g216970 (.A(n_3302),
    .Y(n_3301));
 INVx1_ASAP7_75t_SL g216971 (.A(n_3300),
    .Y(n_3299));
 INVxp67_ASAP7_75t_R g216973 (.A(n_3297),
    .Y(n_3296));
 INVx1_ASAP7_75t_SL g216974 (.A(n_3295),
    .Y(n_3294));
 INVxp67_ASAP7_75t_SL g216975 (.A(n_3293),
    .Y(n_3292));
 INVx1_ASAP7_75t_SL g216976 (.A(n_3291),
    .Y(n_3290));
 INVx2_ASAP7_75t_L g216977 (.A(n_3289),
    .Y(n_3288));
 INVxp33_ASAP7_75t_R g216978 (.A(n_3287),
    .Y(n_3286));
 INVx2_ASAP7_75t_SL g216979 (.A(n_3285),
    .Y(n_3284));
 INVx1_ASAP7_75t_L g216980 (.A(n_3283),
    .Y(n_3282));
 INVx1_ASAP7_75t_SL g216981 (.A(n_3281),
    .Y(n_3280));
 INVx1_ASAP7_75t_L g216982 (.A(n_3279),
    .Y(n_3278));
 INVx2_ASAP7_75t_L g216983 (.A(n_3277),
    .Y(n_3276));
 INVx1_ASAP7_75t_L g216984 (.A(n_3275),
    .Y(n_3274));
 INVxp33_ASAP7_75t_R g216985 (.A(n_3273),
    .Y(n_3272));
 INVx3_ASAP7_75t_SL g216986 (.A(n_3271),
    .Y(n_3270));
 INVx1_ASAP7_75t_SL g216987 (.A(n_3269),
    .Y(n_3268));
 INVx1_ASAP7_75t_L g216993 (.A(n_1732),
    .Y(n_1731));
 INVx2_ASAP7_75t_SL g216994 (.A(n_3267),
    .Y(n_1732));
 INVx1_ASAP7_75t_SL g216995 (.A(n_3266),
    .Y(n_3265));
 INVx1_ASAP7_75t_L g217000 (.A(n_1730),
    .Y(n_1729));
 HB1xp67_ASAP7_75t_L g217002 (.A(n_1730),
    .Y(n_1728));
 INVx1_ASAP7_75t_SL g217003 (.A(n_3263),
    .Y(n_3262));
 INVx2_ASAP7_75t_SL g217004 (.A(n_3261),
    .Y(n_3260));
 INVx2_ASAP7_75t_SL g217005 (.A(n_3259),
    .Y(n_3258));
 INVx1_ASAP7_75t_L g217006 (.A(n_3257),
    .Y(n_3256));
 INVx2_ASAP7_75t_L g217007 (.A(n_3255),
    .Y(n_3254));
 INVx1_ASAP7_75t_SL g217008 (.A(n_3253),
    .Y(n_3252));
 INVxp67_ASAP7_75t_L g217010 (.A(n_1727),
    .Y(n_3251));
 INVx1_ASAP7_75t_L g217012 (.A(n_3249),
    .Y(n_1727));
 INVxp67_ASAP7_75t_R g217014 (.A(n_1726),
    .Y(n_3250));
 BUFx2_ASAP7_75t_SL g217015 (.A(n_3249),
    .Y(n_1726));
 INVx1_ASAP7_75t_L g217016 (.A(n_3248),
    .Y(n_3247));
 INVx2_ASAP7_75t_SL g217017 (.A(n_3246),
    .Y(n_3245));
 INVx2_ASAP7_75t_SL g217018 (.A(n_3244),
    .Y(n_3243));
 INVx3_ASAP7_75t_SL g217019 (.A(n_3242),
    .Y(n_3241));
 NOR2xp33_ASAP7_75t_R g217020 (.A(sa23[7]),
    .B(n_2605),
    .Y(n_3240));
 NAND2xp33_ASAP7_75t_R g217021 (.A(n_8191),
    .B(n_2569),
    .Y(n_3239));
 NAND2xp33_ASAP7_75t_R g217022 (.A(n_2011),
    .B(n_2574),
    .Y(n_3238));
 NAND2xp33_ASAP7_75t_R g217023 (.A(n_2496),
    .B(sa02[7]),
    .Y(n_3237));
 NAND2xp33_ASAP7_75t_R g217024 (.A(n_2477),
    .B(sa30[3]),
    .Y(n_3236));
 NOR2xp33_ASAP7_75t_R g217025 (.A(n_1972),
    .B(n_2212),
    .Y(n_3235));
 NOR2xp33_ASAP7_75t_R g217026 (.A(sa01[3]),
    .B(n_2255),
    .Y(n_3234));
 NOR2xp33_ASAP7_75t_R g217027 (.A(n_1498),
    .B(n_2360),
    .Y(n_3233));
 NAND2xp33_ASAP7_75t_R g217028 (.A(n_1985),
    .B(n_1610),
    .Y(n_3232));
 NOR2xp33_ASAP7_75t_L g217029 (.A(n_1486),
    .B(n_2104),
    .Y(n_3231));
 NOR2xp67_ASAP7_75t_SL g217030 (.A(sa03[1]),
    .B(n_2457),
    .Y(n_3230));
 NOR2xp33_ASAP7_75t_R g217031 (.A(n_2124),
    .B(n_2676),
    .Y(n_3229));
 NOR2xp33_ASAP7_75t_R g217032 (.A(n_1894),
    .B(n_2096),
    .Y(n_3228));
 NOR2xp33_ASAP7_75t_R g217033 (.A(n_1884),
    .B(n_2244),
    .Y(n_3227));
 NAND2xp33_ASAP7_75t_R g217034 (.A(sa22[5]),
    .B(n_2259),
    .Y(n_3226));
 NOR2xp33_ASAP7_75t_R g217035 (.A(sa20[7]),
    .B(n_2577),
    .Y(n_3225));
 NOR2xp33_ASAP7_75t_R g217036 (.A(n_1478),
    .B(n_2468),
    .Y(n_3224));
 NOR2xp33_ASAP7_75t_L g217037 (.A(n_1905),
    .B(n_2539),
    .Y(n_3731));
 NAND2xp5_ASAP7_75t_R g217038 (.A(sa22[4]),
    .B(n_1601),
    .Y(n_3729));
 NOR2xp33_ASAP7_75t_R g217039 (.A(n_1954),
    .B(n_1619),
    .Y(n_3728));
 NAND2xp33_ASAP7_75t_R g217040 (.A(n_1491),
    .B(n_2537),
    .Y(n_3727));
 NAND2xp5_ASAP7_75t_L g217041 (.A(n_2485),
    .B(n_1682),
    .Y(n_3725));
 NAND2xp33_ASAP7_75t_R g217042 (.A(n_1525),
    .B(n_2531),
    .Y(n_3724));
 NOR2xp33_ASAP7_75t_R g217043 (.A(n_2489),
    .B(n_2468),
    .Y(n_3722));
 NOR2xp33_ASAP7_75t_R g217044 (.A(n_2013),
    .B(n_2577),
    .Y(n_3720));
 NAND2xp33_ASAP7_75t_R g217045 (.A(n_2585),
    .B(n_1477),
    .Y(n_3223));
 NOR2xp33_ASAP7_75t_SL g217046 (.A(n_1476),
    .B(n_2555),
    .Y(n_3719));
 NOR2xp33_ASAP7_75t_L g217047 (.A(n_2011),
    .B(n_2535),
    .Y(n_3717));
 NAND2xp5_ASAP7_75t_R g217048 (.A(n_2519),
    .B(n_2015),
    .Y(n_3715));
 NAND2xp5_ASAP7_75t_L g217049 (.A(n_1484),
    .B(n_2512),
    .Y(n_3714));
 NOR2xp33_ASAP7_75t_SL g217050 (.A(sa10[4]),
    .B(n_1618),
    .Y(n_3713));
 NOR2xp33_ASAP7_75t_R g217051 (.A(n_1965),
    .B(n_1582),
    .Y(n_3712));
 NAND2xp33_ASAP7_75t_R g217052 (.A(n_1483),
    .B(n_2508),
    .Y(n_3710));
 NAND2xp5_ASAP7_75t_L g217053 (.A(n_2553),
    .B(n_1880),
    .Y(n_3708));
 NOR2xp33_ASAP7_75t_R g217054 (.A(n_2019),
    .B(n_2510),
    .Y(n_3706));
 NOR2xp33_ASAP7_75t_R g217055 (.A(n_2495),
    .B(n_2449),
    .Y(n_3704));
 NOR2xp33_ASAP7_75t_R g217056 (.A(n_1688),
    .B(n_2470),
    .Y(n_3703));
 NOR2xp33_ASAP7_75t_R g217057 (.A(n_8188),
    .B(n_1369),
    .Y(n_3702));
 NOR2xp33_ASAP7_75t_L g217058 (.A(n_1522),
    .B(n_2524),
    .Y(n_3700));
 NOR2xp33_ASAP7_75t_R g217059 (.A(n_1470),
    .B(n_2501),
    .Y(n_3222));
 NAND2xp33_ASAP7_75t_R g217060 (.A(sa13[7]),
    .B(n_2503),
    .Y(n_3221));
 NOR2xp33_ASAP7_75t_R g217061 (.A(n_2447),
    .B(n_2443),
    .Y(n_3699));
 NAND2xp5_ASAP7_75t_R g217062 (.A(n_2456),
    .B(n_2444),
    .Y(n_3698));
 NOR2xp33_ASAP7_75t_R g217063 (.A(n_1466),
    .B(n_2517),
    .Y(n_3697));
 NAND2xp5_ASAP7_75t_L g217064 (.A(n_2171),
    .B(n_1492),
    .Y(n_1760));
 NOR2xp33_ASAP7_75t_L g217065 (.A(n_1492),
    .B(n_2584),
    .Y(n_3695));
 NOR2xp33_ASAP7_75t_R g217066 (.A(n_1862),
    .B(n_2182),
    .Y(n_3693));
 NAND2xp5_ASAP7_75t_R g217067 (.A(n_2208),
    .B(sa23[1]),
    .Y(n_3692));
 NOR2xp33_ASAP7_75t_R g217068 (.A(n_2499),
    .B(n_2453),
    .Y(n_3691));
 NAND2xp5_ASAP7_75t_R g217069 (.A(n_1478),
    .B(n_1652),
    .Y(n_3690));
 NAND2xp5_ASAP7_75t_SL g217070 (.A(sa03[1]),
    .B(n_1595),
    .Y(n_3689));
 NOR2xp33_ASAP7_75t_R g217071 (.A(n_1873),
    .B(n_2609),
    .Y(n_3688));
 NAND2xp5_ASAP7_75t_L g217072 (.A(n_1535),
    .B(n_2082),
    .Y(n_3687));
 NOR2xp33_ASAP7_75t_L g217073 (.A(n_1534),
    .B(n_2088),
    .Y(n_3686));
 NAND2xp5_ASAP7_75t_SL g217074 (.A(sa10[1]),
    .B(n_2212),
    .Y(n_3685));
 NAND2xp33_ASAP7_75t_R g217075 (.A(sa30[5]),
    .B(n_2189),
    .Y(n_3684));
 NOR2xp33_ASAP7_75t_SL g217076 (.A(n_2023),
    .B(n_1553),
    .Y(n_3682));
 NAND2xp33_ASAP7_75t_R g217077 (.A(sa02[1]),
    .B(n_2400),
    .Y(n_3681));
 NAND2xp33_ASAP7_75t_R g217078 (.A(sa30[5]),
    .B(n_2629),
    .Y(n_3680));
 NOR2xp33_ASAP7_75t_R g217079 (.A(sa23[7]),
    .B(n_2194),
    .Y(n_3679));
 NOR2xp33_ASAP7_75t_R g217080 (.A(sa10[7]),
    .B(n_1337),
    .Y(n_3678));
 NAND2xp33_ASAP7_75t_R g217081 (.A(n_1492),
    .B(n_2389),
    .Y(n_3676));
 NOR2xp67_ASAP7_75t_R g217082 (.A(sa01[7]),
    .B(n_2222),
    .Y(n_3675));
 NOR2xp33_ASAP7_75t_L g217083 (.A(n_1873),
    .B(n_2250),
    .Y(n_3674));
 NOR2xp33_ASAP7_75t_SL g217084 (.A(n_8202),
    .B(n_1698),
    .Y(n_3673));
 NAND2xp33_ASAP7_75t_R g217085 (.A(sa01[7]),
    .B(n_1691),
    .Y(n_3671));
 NAND2xp5_ASAP7_75t_L g217086 (.A(n_1476),
    .B(n_2215),
    .Y(n_3669));
 NOR2xp33_ASAP7_75t_R g217087 (.A(sa10[1]),
    .B(n_1551),
    .Y(n_3668));
 NAND2xp5_ASAP7_75t_L g217088 (.A(sa03[1]),
    .B(n_2046),
    .Y(n_3667));
 NOR2xp33_ASAP7_75t_SL g217089 (.A(n_1535),
    .B(n_2533),
    .Y(n_3665));
 NAND2xp5_ASAP7_75t_R g217090 (.A(sa10[7]),
    .B(n_2525),
    .Y(n_3664));
 NAND2xp5_ASAP7_75t_R g217091 (.A(n_1912),
    .B(n_2611),
    .Y(n_3663));
 NAND2xp5_ASAP7_75t_L g217092 (.A(sa21[5]),
    .B(n_2632),
    .Y(n_3662));
 NAND2xp33_ASAP7_75t_R g217093 (.A(n_1912),
    .B(n_1608),
    .Y(n_3661));
 NOR2xp33_ASAP7_75t_R g217094 (.A(n_1491),
    .B(n_2091),
    .Y(n_3660));
 NAND2xp33_ASAP7_75t_R g217095 (.A(n_1905),
    .B(n_1451),
    .Y(n_3220));
 NAND2xp33_ASAP7_75t_R g217096 (.A(n_1683),
    .B(n_2440),
    .Y(n_3659));
 AND2x2_ASAP7_75t_R g217097 (.A(n_1525),
    .B(n_2084),
    .Y(n_3658));
 NAND2xp33_ASAP7_75t_R g217098 (.A(n_1522),
    .B(n_1350),
    .Y(n_3657));
 NAND2xp5_ASAP7_75t_SL g217099 (.A(n_1876),
    .B(n_2166),
    .Y(n_3655));
 NAND2xp5_ASAP7_75t_L g217100 (.A(n_1524),
    .B(n_2205),
    .Y(n_3654));
 NAND2xp5_ASAP7_75t_L g217101 (.A(n_2015),
    .B(n_1576),
    .Y(n_3653));
 NOR2xp33_ASAP7_75t_L g217102 (.A(n_1482),
    .B(n_1342),
    .Y(n_3651));
 AND2x2_ASAP7_75t_R g217103 (.A(n_1904),
    .B(n_2040),
    .Y(n_3650));
 NAND2xp5_ASAP7_75t_R g217104 (.A(n_2051),
    .B(n_1524),
    .Y(n_3648));
 NAND2xp33_ASAP7_75t_R g217105 (.A(sa23[7]),
    .B(n_2527),
    .Y(n_3647));
 NOR2xp33_ASAP7_75t_SL g217106 (.A(n_8207),
    .B(n_2565),
    .Y(n_3646));
 NAND2xp5_ASAP7_75t_R g217107 (.A(n_2119),
    .B(n_1522),
    .Y(n_3644));
 AND2x2_ASAP7_75t_R g217108 (.A(sa12[7]),
    .B(n_2064),
    .Y(n_3642));
 NOR2xp33_ASAP7_75t_L g217109 (.A(n_1987),
    .B(n_2195),
    .Y(n_3641));
 NAND2xp5_ASAP7_75t_R g217110 (.A(sa12[1]),
    .B(n_2197),
    .Y(n_3639));
 NOR2xp33_ASAP7_75t_R g217111 (.A(sa23[4]),
    .B(n_2298),
    .Y(n_3638));
 NOR2xp33_ASAP7_75t_L g217112 (.A(sa02[7]),
    .B(n_2074),
    .Y(n_3637));
 NAND2xp33_ASAP7_75t_R g217113 (.A(n_2014),
    .B(n_2416),
    .Y(n_3636));
 NOR2xp33_ASAP7_75t_R g217114 (.A(sa21[7]),
    .B(n_2073),
    .Y(n_3635));
 NAND2xp5_ASAP7_75t_L g217115 (.A(n_2019),
    .B(n_1609),
    .Y(n_3633));
 NOR2xp33_ASAP7_75t_R g217116 (.A(sa20[7]),
    .B(n_2217),
    .Y(n_3632));
 NOR2xp33_ASAP7_75t_R g217117 (.A(n_1879),
    .B(n_1696),
    .Y(n_3631));
 NAND2xp5_ASAP7_75t_R g217118 (.A(sa02[7]),
    .B(n_2400),
    .Y(n_3630));
 NAND2xp5_ASAP7_75t_L g217119 (.A(n_1576),
    .B(n_1530),
    .Y(n_3629));
 NAND2xp5_ASAP7_75t_L g217120 (.A(n_1482),
    .B(n_2241),
    .Y(n_3628));
 NOR2xp33_ASAP7_75t_L g217121 (.A(n_2014),
    .B(n_1580),
    .Y(n_3627));
 NAND2xp5_ASAP7_75t_R g217122 (.A(n_1470),
    .B(n_2397),
    .Y(n_3625));
 NAND2xp5_ASAP7_75t_R g217123 (.A(sa23[4]),
    .B(n_2138),
    .Y(n_3623));
 NAND2xp33_ASAP7_75t_R g217124 (.A(sa23[5]),
    .B(n_2598),
    .Y(n_3622));
 NAND2xp33_ASAP7_75t_R g217125 (.A(n_1473),
    .B(n_1436),
    .Y(n_3621));
 NAND2xp5_ASAP7_75t_L g217126 (.A(n_1485),
    .B(n_2079),
    .Y(n_3620));
 NAND2xp5_ASAP7_75t_R g217127 (.A(n_1526),
    .B(n_2084),
    .Y(n_3619));
 NAND2xp33_ASAP7_75t_R g217128 (.A(n_2176),
    .B(n_1472),
    .Y(n_1759));
 NOR2xp33_ASAP7_75t_R g217129 (.A(n_1879),
    .B(n_2204),
    .Y(n_3618));
 NAND2xp5_ASAP7_75t_L g217130 (.A(sa10[1]),
    .B(n_2110),
    .Y(n_3617));
 NAND2xp5_ASAP7_75t_L g217131 (.A(n_1605),
    .B(sa02[1]),
    .Y(n_3616));
 NOR2xp33_ASAP7_75t_SL g217132 (.A(n_1513),
    .B(n_2160),
    .Y(n_3614));
 AND2x2_ASAP7_75t_R g217133 (.A(n_1476),
    .B(n_1445),
    .Y(n_3613));
 NAND2xp5_ASAP7_75t_R g217134 (.A(n_2218),
    .B(n_1466),
    .Y(n_3612));
 NAND2xp33_ASAP7_75t_R g217135 (.A(n_1855),
    .B(n_2294),
    .Y(n_3611));
 NAND2xp33_ASAP7_75t_R g217136 (.A(sa13[7]),
    .B(n_2392),
    .Y(n_3609));
 NOR2xp33_ASAP7_75t_R g217137 (.A(n_1884),
    .B(n_2602),
    .Y(n_3607));
 NAND2xp5_ASAP7_75t_R g217138 (.A(n_8912),
    .B(n_2317),
    .Y(n_3606));
 NOR2xp33_ASAP7_75t_L g217139 (.A(n_1706),
    .B(n_2532),
    .Y(n_3605));
 AND2x2_ASAP7_75t_R g217140 (.A(n_1506),
    .B(n_2137),
    .Y(n_3603));
 NAND2xp33_ASAP7_75t_R g217141 (.A(n_2067),
    .B(sa02[0]),
    .Y(n_3602));
 NAND2xp5_ASAP7_75t_R g217142 (.A(n_1709),
    .B(n_2578),
    .Y(n_3600));
 NOR2xp33_ASAP7_75t_SL g217143 (.A(sa10[1]),
    .B(n_2506),
    .Y(n_3599));
 NAND2xp5_ASAP7_75t_SL g217144 (.A(n_1492),
    .B(n_2255),
    .Y(n_3597));
 NAND2xp5_ASAP7_75t_R g217145 (.A(n_1510),
    .B(n_1439),
    .Y(n_3596));
 NAND2xp5_ASAP7_75t_R g217146 (.A(n_2033),
    .B(n_2273),
    .Y(n_3595));
 NOR2xp33_ASAP7_75t_L g217147 (.A(n_1517),
    .B(n_2515),
    .Y(n_3594));
 NOR2xp33_ASAP7_75t_L g217148 (.A(n_2644),
    .B(n_2437),
    .Y(n_3593));
 NOR2x1_ASAP7_75t_SL g217149 (.A(n_2489),
    .B(n_2507),
    .Y(n_3591));
 NOR2xp33_ASAP7_75t_L g217150 (.A(sa20[5]),
    .B(n_2283),
    .Y(n_3590));
 NOR2xp33_ASAP7_75t_L g217151 (.A(n_2642),
    .B(n_2528),
    .Y(n_3589));
 NAND2xp5_ASAP7_75t_L g217152 (.A(sa10[4]),
    .B(n_2210),
    .Y(n_3587));
 NOR2xp33_ASAP7_75t_L g217153 (.A(n_1487),
    .B(n_2567),
    .Y(n_3586));
 NAND2xp5_ASAP7_75t_R g217154 (.A(n_1873),
    .B(n_2267),
    .Y(n_3585));
 NAND2xp33_ASAP7_75t_R g217155 (.A(n_8209),
    .B(n_2239),
    .Y(n_3582));
 NOR2xp33_ASAP7_75t_SL g217156 (.A(n_1481),
    .B(n_2562),
    .Y(n_3580));
 NAND2xp5_ASAP7_75t_SL g217157 (.A(n_2226),
    .B(n_1479),
    .Y(n_1758));
 NOR2xp67_ASAP7_75t_L g217158 (.A(n_8183),
    .B(n_1700),
    .Y(n_3579));
 NOR2xp33_ASAP7_75t_SL g217159 (.A(n_1994),
    .B(n_2530),
    .Y(n_1757));
 NOR2xp33_ASAP7_75t_SL g217160 (.A(n_2201),
    .B(n_8207),
    .Y(n_3578));
 NAND2xp5_ASAP7_75t_R g217161 (.A(n_2022),
    .B(n_2277),
    .Y(n_3577));
 NOR2xp33_ASAP7_75t_SL g217162 (.A(n_2626),
    .B(n_1895),
    .Y(n_3575));
 NAND2xp5_ASAP7_75t_SL g217163 (.A(n_2503),
    .B(n_2651),
    .Y(n_3573));
 NAND2xp5_ASAP7_75t_SL g217164 (.A(n_1487),
    .B(n_1643),
    .Y(n_3572));
 NOR2xp33_ASAP7_75t_L g217165 (.A(n_2020),
    .B(n_2228),
    .Y(n_3569));
 NOR2xp33_ASAP7_75t_L g217166 (.A(n_1913),
    .B(n_2595),
    .Y(n_3568));
 NOR2xp67_ASAP7_75t_L g217167 (.A(n_2674),
    .B(n_2507),
    .Y(n_1756));
 AND2x2_ASAP7_75t_L g217168 (.A(n_1473),
    .B(n_2230),
    .Y(n_3566));
 NAND2xp5_ASAP7_75t_L g217169 (.A(n_2242),
    .B(n_1487),
    .Y(n_3565));
 NOR2xp33_ASAP7_75t_SL g217170 (.A(n_1982),
    .B(n_2235),
    .Y(n_3562));
 NAND2xp5_ASAP7_75t_R g217171 (.A(sa02[5]),
    .B(n_2224),
    .Y(n_3561));
 NOR2xp33_ASAP7_75t_SL g217172 (.A(n_2472),
    .B(n_2520),
    .Y(n_3560));
 NAND2xp5_ASAP7_75t_R g217173 (.A(n_8183),
    .B(n_2649),
    .Y(n_3558));
 NOR2xp33_ASAP7_75t_R g217174 (.A(sa22[5]),
    .B(n_2260),
    .Y(n_3557));
 NAND2xp5_ASAP7_75t_R g217175 (.A(n_1701),
    .B(n_1689),
    .Y(n_3556));
 NOR2x1_ASAP7_75t_R g217176 (.A(n_1707),
    .B(n_2510),
    .Y(n_3555));
 NAND2xp5_ASAP7_75t_R g217177 (.A(n_8202),
    .B(n_2258),
    .Y(n_3554));
 NAND2xp5_ASAP7_75t_R g217178 (.A(n_1470),
    .B(n_2247),
    .Y(n_3552));
 NAND2xp33_ASAP7_75t_R g217179 (.A(n_1479),
    .B(n_1659),
    .Y(n_3551));
 NAND2xp5_ASAP7_75t_R g217180 (.A(n_2022),
    .B(n_2601),
    .Y(n_3550));
 NOR2xp33_ASAP7_75t_R g217181 (.A(sa33[5]),
    .B(n_2265),
    .Y(n_3548));
 NAND2xp33_ASAP7_75t_R g217182 (.A(n_1471),
    .B(n_2054),
    .Y(n_3547));
 NAND2xp5_ASAP7_75t_L g217183 (.A(n_1905),
    .B(n_2540),
    .Y(n_3546));
 NAND2xp33_ASAP7_75t_R g217184 (.A(n_1493),
    .B(n_2058),
    .Y(n_3545));
 NAND2xp33_ASAP7_75t_R g217185 (.A(n_2245),
    .B(n_1884),
    .Y(n_3543));
 NOR2x1_ASAP7_75t_R g217186 (.A(n_1995),
    .B(n_2249),
    .Y(n_3542));
 NAND2xp5_ASAP7_75t_L g217187 (.A(n_2645),
    .B(n_2525),
    .Y(n_3541));
 NOR2xp33_ASAP7_75t_L g217188 (.A(sa03[1]),
    .B(n_2588),
    .Y(n_3539));
 NOR2xp33_ASAP7_75t_L g217189 (.A(n_1917),
    .B(n_2686),
    .Y(n_3538));
 NAND2xp5_ASAP7_75t_R g217190 (.A(n_1478),
    .B(n_2254),
    .Y(n_3536));
 NAND2xp5_ASAP7_75t_SL g217191 (.A(n_1475),
    .B(n_2269),
    .Y(n_3534));
 NOR2x1_ASAP7_75t_L g217192 (.A(n_2463),
    .B(n_2510),
    .Y(n_3533));
 NAND2x1_ASAP7_75t_SL g217193 (.A(n_1862),
    .B(n_2219),
    .Y(n_3532));
 NOR2xp67_ASAP7_75t_L g217194 (.A(n_1706),
    .B(n_2486),
    .Y(n_3530));
 NAND2xp5_ASAP7_75t_SL g217195 (.A(n_1480),
    .B(n_2227),
    .Y(n_1755));
 OR2x2_ASAP7_75t_L g217196 (.A(sa12[1]),
    .B(n_2196),
    .Y(n_3528));
 AND2x2_ASAP7_75t_SL g217197 (.A(n_1992),
    .B(n_2249),
    .Y(n_3527));
 AND2x2_ASAP7_75t_L g217198 (.A(n_1513),
    .B(n_2160),
    .Y(n_3526));
 NAND2xp5_ASAP7_75t_SL g217199 (.A(n_8212),
    .B(n_2123),
    .Y(n_3524));
 NAND2xp5_ASAP7_75t_R g217200 (.A(n_1701),
    .B(n_2456),
    .Y(n_3523));
 NAND2xp5_ASAP7_75t_SL g217201 (.A(n_1709),
    .B(n_2452),
    .Y(n_3521));
 OR2x2_ASAP7_75t_SL g217202 (.A(n_1523),
    .B(n_2524),
    .Y(n_3519));
 AND2x2_ASAP7_75t_SL g217203 (.A(n_1522),
    .B(n_2253),
    .Y(n_3517));
 NAND2xp5_ASAP7_75t_L g217204 (.A(n_1487),
    .B(n_2568),
    .Y(n_3516));
 AND2x2_ASAP7_75t_L g217205 (.A(n_1486),
    .B(n_2243),
    .Y(n_3514));
 NAND2xp5_ASAP7_75t_R g217206 (.A(n_2009),
    .B(n_2262),
    .Y(n_3513));
 AND2x2_ASAP7_75t_SL g217207 (.A(n_1953),
    .B(n_2319),
    .Y(n_3511));
 NOR2xp67_ASAP7_75t_L g217208 (.A(n_1895),
    .B(n_2614),
    .Y(n_3509));
 NAND2xp5_ASAP7_75t_R g217209 (.A(n_1884),
    .B(n_2152),
    .Y(n_3508));
 NOR2xp67_ASAP7_75t_L g217210 (.A(sa12[1]),
    .B(n_2576),
    .Y(n_1754));
 OR2x2_ASAP7_75t_L g217211 (.A(n_2650),
    .B(n_2451),
    .Y(n_3506));
 AND2x2_ASAP7_75t_L g217212 (.A(n_1950),
    .B(n_2286),
    .Y(n_3504));
 NAND2xp5_ASAP7_75t_L g217213 (.A(n_1523),
    .B(n_2121),
    .Y(n_3502));
 NAND2xp5_ASAP7_75t_SL g217214 (.A(n_8212),
    .B(n_1619),
    .Y(n_3501));
 NAND2x1_ASAP7_75t_SL g217215 (.A(n_8912),
    .B(n_2318),
    .Y(n_3499));
 AND2x2_ASAP7_75t_SL g217216 (.A(n_1880),
    .B(n_2231),
    .Y(n_3497));
 NAND2xp5_ASAP7_75t_L g217217 (.A(n_1708),
    .B(n_2481),
    .Y(n_1753));
 NAND2xp5_ASAP7_75t_L g217218 (.A(n_2287),
    .B(n_1952),
    .Y(n_3495));
 NOR2xp33_ASAP7_75t_SL g217219 (.A(sa23[5]),
    .B(n_2156),
    .Y(n_3493));
 AND2x2_ASAP7_75t_SL g217220 (.A(n_1505),
    .B(n_1615),
    .Y(n_3492));
 NAND2xp5_ASAP7_75t_L g217221 (.A(n_1469),
    .B(n_1610),
    .Y(n_3491));
 NOR2xp33_ASAP7_75t_SL g217222 (.A(n_2275),
    .B(n_1905),
    .Y(n_3490));
 AND2x2_ASAP7_75t_SL g217223 (.A(n_2020),
    .B(n_2228),
    .Y(n_3489));
 AND2x2_ASAP7_75t_SL g217224 (.A(n_1982),
    .B(n_2235),
    .Y(n_3488));
 NAND2xp5_ASAP7_75t_SL g217225 (.A(n_1477),
    .B(n_1611),
    .Y(n_3486));
 NAND2xp5_ASAP7_75t_L g217226 (.A(n_1871),
    .B(n_2213),
    .Y(n_3485));
 NOR2x1_ASAP7_75t_L g217227 (.A(n_2445),
    .B(n_2511),
    .Y(n_3483));
 NOR2xp33_ASAP7_75t_L g217228 (.A(n_2642),
    .B(n_2470),
    .Y(n_3480));
 NAND2xp5_ASAP7_75t_R g217229 (.A(sa20[5]),
    .B(n_2284),
    .Y(n_3479));
 NAND2xp33_ASAP7_75t_R g217230 (.A(n_8204),
    .B(n_2062),
    .Y(n_3477));
 NOR2x1p5_ASAP7_75t_L g217231 (.A(n_1487),
    .B(n_2103),
    .Y(n_3476));
 NAND2xp5_ASAP7_75t_L g217232 (.A(n_1493),
    .B(n_2256),
    .Y(n_3474));
 NAND2xp5_ASAP7_75t_R g217233 (.A(sa20[5]),
    .B(n_2656),
    .Y(n_3473));
 NAND2xp5_ASAP7_75t_SL g217234 (.A(n_1959),
    .B(n_2137),
    .Y(n_3470));
 AND2x2_ASAP7_75t_L g217235 (.A(n_1513),
    .B(n_2209),
    .Y(n_3469));
 NAND2xp5_ASAP7_75t_R g217236 (.A(n_8183),
    .B(n_2632),
    .Y(n_3467));
 NAND2xp5_ASAP7_75t_SL g217237 (.A(n_2467),
    .B(n_2675),
    .Y(n_3465));
 AND2x2_ASAP7_75t_R g217238 (.A(n_1862),
    .B(n_2182),
    .Y(n_3463));
 NOR2xp33_ASAP7_75t_L g217239 (.A(sa20[5]),
    .B(n_2233),
    .Y(n_3462));
 AND2x2_ASAP7_75t_L g217240 (.A(n_1960),
    .B(n_1618),
    .Y(n_3461));
 NOR2xp33_ASAP7_75t_L g217241 (.A(sa23[4]),
    .B(n_1617),
    .Y(n_3459));
 NAND2xp5_ASAP7_75t_L g217242 (.A(n_1895),
    .B(n_2627),
    .Y(n_3457));
 NAND2xp5_ASAP7_75t_SL g217243 (.A(sa23[1]),
    .B(n_2514),
    .Y(n_3455));
 AND2x2_ASAP7_75t_SL g217244 (.A(n_1862),
    .B(n_2517),
    .Y(n_3454));
 AND2x2_ASAP7_75t_R g217245 (.A(n_1466),
    .B(n_2518),
    .Y(n_3453));
 NAND2xp5_ASAP7_75t_L g217246 (.A(n_8197),
    .B(n_2601),
    .Y(n_3452));
 NOR2x1_ASAP7_75t_L g217247 (.A(n_1871),
    .B(n_2506),
    .Y(n_3451));
 NOR2xp67_ASAP7_75t_SL g217248 (.A(n_2447),
    .B(n_1690),
    .Y(n_3449));
 NAND2xp5_ASAP7_75t_SL g217249 (.A(n_1855),
    .B(n_2295),
    .Y(n_3447));
 NAND2xp5_ASAP7_75t_R g217250 (.A(n_2033),
    .B(n_2189),
    .Y(n_3445));
 NOR2xp33_ASAP7_75t_L g217251 (.A(n_1917),
    .B(n_2233),
    .Y(n_3443));
 NOR2x1_ASAP7_75t_SL g217252 (.A(n_1674),
    .B(n_2504),
    .Y(n_1752));
 NAND2xp5_ASAP7_75t_L g217253 (.A(n_1913),
    .B(n_2596),
    .Y(n_3440));
 NAND2xp5_ASAP7_75t_SL g217254 (.A(n_2162),
    .B(n_1855),
    .Y(n_3437));
 NAND2x1_ASAP7_75t_SL g217255 (.A(n_1856),
    .B(n_2139),
    .Y(n_1751));
 OR2x2_ASAP7_75t_SL g217256 (.A(n_1522),
    .B(n_2253),
    .Y(n_3435));
 OR2x2_ASAP7_75t_L g217257 (.A(n_1856),
    .B(n_1617),
    .Y(n_1750));
 NAND2xp5_ASAP7_75t_L g217258 (.A(n_1954),
    .B(n_1619),
    .Y(n_3432));
 NAND2xp5_ASAP7_75t_R g217259 (.A(n_8207),
    .B(n_2566),
    .Y(n_3431));
 NAND2xp5_ASAP7_75t_SL g217260 (.A(sa10[4]),
    .B(n_1618),
    .Y(n_3429));
 OR2x2_ASAP7_75t_SL g217261 (.A(n_8899),
    .B(n_2113),
    .Y(n_3427));
 NAND2xp5_ASAP7_75t_SL g217262 (.A(n_1994),
    .B(n_2529),
    .Y(n_3425));
 AND2x2_ASAP7_75t_SL g217263 (.A(sa22[4]),
    .B(n_2295),
    .Y(n_3424));
 AND2x2_ASAP7_75t_L g217264 (.A(n_1470),
    .B(n_2502),
    .Y(n_3423));
 AND2x2_ASAP7_75t_SL g217265 (.A(n_8896),
    .B(n_2318),
    .Y(n_3421));
 NAND2x1p5_ASAP7_75t_SL g217266 (.A(n_8212),
    .B(n_2122),
    .Y(n_3419));
 NAND2xp5_ASAP7_75t_SL g217267 (.A(n_1852),
    .B(n_2639),
    .Y(n_3416));
 NAND2xp5_ASAP7_75t_SL g217268 (.A(sa12[4]),
    .B(n_2319),
    .Y(n_3415));
 NAND2xp5_ASAP7_75t_SL g217269 (.A(n_1476),
    .B(n_2556),
    .Y(n_3414));
 NAND2x1_ASAP7_75t_SL g217270 (.A(n_1474),
    .B(n_2214),
    .Y(n_1748));
 NAND2xp5_ASAP7_75t_R g217271 (.A(n_2542),
    .B(n_8209),
    .Y(n_3411));
 NOR2xp33_ASAP7_75t_R g217272 (.A(sa33[5]),
    .B(n_2582),
    .Y(n_3409));
 AND2x2_ASAP7_75t_SL g217273 (.A(n_8912),
    .B(n_2118),
    .Y(n_3407));
 NAND2xp33_ASAP7_75t_R g217274 (.A(n_8190),
    .B(n_2611),
    .Y(n_3405));
 NAND2x1_ASAP7_75t_L g217275 (.A(n_1953),
    .B(n_2133),
    .Y(n_1746));
 NAND2xp5_ASAP7_75t_L g217276 (.A(n_1895),
    .B(n_2615),
    .Y(n_3402));
 NOR2xp33_ASAP7_75t_SL g217277 (.A(n_2609),
    .B(sa32[5]),
    .Y(n_3401));
 AND2x2_ASAP7_75t_R g217278 (.A(n_1884),
    .B(n_2603),
    .Y(n_3399));
 NAND2x1_ASAP7_75t_SL g217279 (.A(n_1871),
    .B(n_2111),
    .Y(n_1745));
 OR2x2_ASAP7_75t_SL g217280 (.A(sa03[4]),
    .B(n_1701),
    .Y(n_3396));
 AND2x4_ASAP7_75t_SL g217281 (.A(n_1987),
    .B(n_2576),
    .Y(n_3394));
 NOR2x1_ASAP7_75t_SL g217282 (.A(sa33[5]),
    .B(n_2164),
    .Y(n_3392));
 AND2x2_ASAP7_75t_L g217283 (.A(n_8207),
    .B(n_2202),
    .Y(n_3390));
 NAND2xp5_ASAP7_75t_SL g217284 (.A(n_1513),
    .B(n_2515),
    .Y(n_3387));
 AND2x2_ASAP7_75t_SL g217285 (.A(n_8908),
    .B(n_2619),
    .Y(n_3386));
 NOR2xp33_ASAP7_75t_SL g217286 (.A(sa20[5]),
    .B(n_2657),
    .Y(n_3384));
 NOR2x1_ASAP7_75t_L g217287 (.A(sa22[5]),
    .B(n_2204),
    .Y(n_3382));
 NAND2x1_ASAP7_75t_SL g217288 (.A(n_8200),
    .B(n_2675),
    .Y(n_1743));
 NAND2x1_ASAP7_75t_SL g217289 (.A(n_1480),
    .B(n_2562),
    .Y(n_3380));
 NOR2xp33_ASAP7_75t_SL g217290 (.A(sa00[5]),
    .B(n_2616),
    .Y(n_3378));
 AND2x2_ASAP7_75t_SL g217291 (.A(n_8202),
    .B(n_2184),
    .Y(n_3376));
 NAND2xp5_ASAP7_75t_L g217292 (.A(n_1948),
    .B(n_1701),
    .Y(n_3374));
 AND2x2_ASAP7_75t_SL g217293 (.A(n_1960),
    .B(n_2211),
    .Y(n_3372));
 NAND2x1_ASAP7_75t_SL g217294 (.A(n_1855),
    .B(n_1704),
    .Y(n_3370));
 AND2x2_ASAP7_75t_SL g217295 (.A(n_1949),
    .B(n_1699),
    .Y(n_3368));
 AND2x2_ASAP7_75t_SL g217296 (.A(n_1891),
    .B(n_2586),
    .Y(n_3366));
 AND2x2_ASAP7_75t_L g217297 (.A(n_1856),
    .B(n_1686),
    .Y(n_3364));
 NAND2x1_ASAP7_75t_SL g217298 (.A(n_1683),
    .B(n_1855),
    .Y(n_3361));
 NOR2xp33_ASAP7_75t_L g217299 (.A(sa22[5]),
    .B(n_1696),
    .Y(n_3360));
 AND2x2_ASAP7_75t_SL g217300 (.A(n_1873),
    .B(n_2251),
    .Y(n_3358));
 NAND2xp5_ASAP7_75t_SL g217301 (.A(n_8189),
    .B(n_1695),
    .Y(n_1741));
 AND2x2_ASAP7_75t_L g217302 (.A(n_1502),
    .B(n_2637),
    .Y(n_3356));
 NOR2x1p5_ASAP7_75t_SL g217303 (.A(sa02[5]),
    .B(n_2225),
    .Y(n_1740));
 AND2x2_ASAP7_75t_L g217304 (.A(n_1856),
    .B(n_2643),
    .Y(n_3355));
 AND2x2_ASAP7_75t_SL g217305 (.A(n_2033),
    .B(n_2629),
    .Y(n_3353));
 NAND2xp5_ASAP7_75t_L g217306 (.A(n_2009),
    .B(n_2598),
    .Y(n_3351));
 NAND2xp5_ASAP7_75t_L g217307 (.A(n_8209),
    .B(n_2191),
    .Y(n_1738));
 NOR2xp33_ASAP7_75t_SL g217308 (.A(n_1360),
    .B(n_2659),
    .Y(n_3349));
 AND2x2_ASAP7_75t_SL g217309 (.A(n_1852),
    .B(n_2640),
    .Y(n_3347));
 NAND2xp5_ASAP7_75t_L g217310 (.A(n_8204),
    .B(n_2102),
    .Y(n_3344));
 AND2x2_ASAP7_75t_SL g217311 (.A(n_8197),
    .B(n_2277),
    .Y(n_3343));
 NAND2xp5_ASAP7_75t_L g217312 (.A(n_1471),
    .B(n_2165),
    .Y(n_3340));
 NAND2xp5_ASAP7_75t_SL g217313 (.A(n_8190),
    .B(n_2236),
    .Y(n_3338));
 NAND2x1p5_ASAP7_75t_SL g217314 (.A(n_1952),
    .B(n_2633),
    .Y(n_1736));
 OR2x2_ASAP7_75t_L g217315 (.A(sa21[5]),
    .B(n_1700),
    .Y(n_3336));
 NAND2x1_ASAP7_75t_SL g217316 (.A(n_1982),
    .B(n_2522),
    .Y(n_3334));
 AND2x2_ASAP7_75t_SL g217317 (.A(n_1959),
    .B(n_2651),
    .Y(n_3332));
 NAND2x1p5_ASAP7_75t_SL g217318 (.A(n_1871),
    .B(n_2506),
    .Y(n_3329));
 AND2x2_ASAP7_75t_SL g217319 (.A(n_1466),
    .B(n_2453),
    .Y(n_3327));
 NAND2x1p5_ASAP7_75t_SL g217320 (.A(n_1953),
    .B(n_1708),
    .Y(n_1735));
 NAND2x1_ASAP7_75t_SL g217321 (.A(n_1517),
    .B(n_2470),
    .Y(n_3324));
 AND2x2_ASAP7_75t_SL g217322 (.A(n_1960),
    .B(n_2645),
    .Y(n_3322));
 AND2x2_ASAP7_75t_SL g217323 (.A(n_8212),
    .B(n_2618),
    .Y(n_3320));
 NAND2xp5_ASAP7_75t_SL g217324 (.A(n_1384),
    .B(n_2607),
    .Y(n_3316));
 AND2x2_ASAP7_75t_SL g217325 (.A(n_1425),
    .B(n_1701),
    .Y(n_3315));
 AND2x2_ASAP7_75t_L g217326 (.A(n_1960),
    .B(n_2488),
    .Y(n_3313));
 AND2x2_ASAP7_75t_SL g217327 (.A(n_1958),
    .B(n_2651),
    .Y(n_3311));
 AND2x2_ASAP7_75t_SL g217328 (.A(sa12[4]),
    .B(n_1708),
    .Y(n_3309));
 AND2x4_ASAP7_75t_SL g217329 (.A(sa31[4]),
    .B(n_2640),
    .Y(n_3307));
 NAND2xp5_ASAP7_75t_SL g217330 (.A(sa23[4]),
    .B(n_2643),
    .Y(n_1733));
 NAND2x1_ASAP7_75t_SL g217331 (.A(sa23[4]),
    .B(n_2139),
    .Y(n_3304));
 NAND2x1_ASAP7_75t_SL g217332 (.A(n_1954),
    .B(n_2618),
    .Y(n_3302));
 OR2x2_ASAP7_75t_SL g217333 (.A(n_1950),
    .B(n_2106),
    .Y(n_3300));
 AND2x4_ASAP7_75t_SL g217334 (.A(n_1853),
    .B(n_2675),
    .Y(n_3298));
 OR2x2_ASAP7_75t_SL g217335 (.A(n_1954),
    .B(n_2465),
    .Y(n_3297));
 AND2x2_ASAP7_75t_SL g217336 (.A(sa20[4]),
    .B(n_2658),
    .Y(n_3295));
 AND2x2_ASAP7_75t_SL g217337 (.A(n_1880),
    .B(n_2554),
    .Y(n_3293));
 NAND2xp5_ASAP7_75t_SL g217338 (.A(n_1953),
    .B(n_2462),
    .Y(n_3291));
 NAND2x1p5_ASAP7_75t_SL g217339 (.A(sa10[4]),
    .B(n_2645),
    .Y(n_3289));
 NAND2x1_ASAP7_75t_L g217340 (.A(n_1995),
    .B(n_2530),
    .Y(n_3287));
 AND2x2_ASAP7_75t_SL g217341 (.A(sa10[1]),
    .B(n_2437),
    .Y(n_3285));
 OR2x2_ASAP7_75t_SL g217342 (.A(n_1982),
    .B(n_2439),
    .Y(n_3283));
 NAND2x1p5_ASAP7_75t_SL g217343 (.A(n_1471),
    .B(n_2501),
    .Y(n_3281));
 AND2x2_ASAP7_75t_SL g217344 (.A(sa22[4]),
    .B(n_2635),
    .Y(n_3279));
 AND2x4_ASAP7_75t_SL g217345 (.A(n_1473),
    .B(n_2451),
    .Y(n_3277));
 OR2x2_ASAP7_75t_SL g217346 (.A(n_2463),
    .B(n_2655),
    .Y(n_3275));
 AND2x4_ASAP7_75t_SL g217347 (.A(n_2488),
    .B(n_2645),
    .Y(n_3273));
 NAND2x2_ASAP7_75t_SL g217348 (.A(n_2658),
    .B(n_2500),
    .Y(n_3271));
 AND2x2_ASAP7_75t_SL g217349 (.A(n_1481),
    .B(n_2474),
    .Y(n_3269));
 NAND2x1p5_ASAP7_75t_SL g217350 (.A(n_1701),
    .B(n_2444),
    .Y(n_3267));
 AND2x2_ASAP7_75t_SL g217351 (.A(n_1686),
    .B(n_2643),
    .Y(n_3266));
 NAND2x1_ASAP7_75t_SL g217352 (.A(sa32[4]),
    .B(n_2112),
    .Y(n_1730));
 AND2x4_ASAP7_75t_SL g217353 (.A(sa12[1]),
    .B(n_2482),
    .Y(n_3263));
 AND2x2_ASAP7_75t_SL g217354 (.A(sa10[4]),
    .B(n_2211),
    .Y(n_3261));
 AND2x2_ASAP7_75t_SL g217355 (.A(n_1958),
    .B(n_2136),
    .Y(n_3259));
 NAND2x1p5_ASAP7_75t_SL g217356 (.A(n_2441),
    .B(n_1470),
    .Y(n_3257));
 AND2x4_ASAP7_75t_SL g217357 (.A(n_1994),
    .B(n_2449),
    .Y(n_3255));
 OR2x2_ASAP7_75t_SL g217358 (.A(n_1855),
    .B(n_2161),
    .Y(n_3253));
 NAND2xp5_ASAP7_75t_SL g217359 (.A(n_2459),
    .B(n_2651),
    .Y(n_3249));
 AND2x4_ASAP7_75t_SL g217360 (.A(n_1954),
    .B(n_2122),
    .Y(n_3248));
 NAND2x1_ASAP7_75t_SL g217361 (.A(n_1890),
    .B(n_2468),
    .Y(n_3246));
 AND2x4_ASAP7_75t_SL g217362 (.A(sa12[4]),
    .B(n_2132),
    .Y(n_3244));
 AND2x2_ASAP7_75t_SL g217363 (.A(n_2479),
    .B(n_1338),
    .Y(n_3242));
 INVxp33_ASAP7_75t_R g217364 (.A(n_3217),
    .Y(n_3218));
 INVxp33_ASAP7_75t_R g217365 (.A(n_3213),
    .Y(n_3214));
 INVxp67_ASAP7_75t_R g217366 (.A(n_3199),
    .Y(n_3200));
 INVxp67_ASAP7_75t_L g217367 (.A(n_3191),
    .Y(n_3192));
 INVxp33_ASAP7_75t_R g217368 (.A(n_3187),
    .Y(n_3188));
 INVxp33_ASAP7_75t_R g217369 (.A(n_3180),
    .Y(n_3181));
 INVxp33_ASAP7_75t_R g217370 (.A(n_3177),
    .Y(n_3178));
 INVxp33_ASAP7_75t_R g217371 (.A(n_3175),
    .Y(n_3176));
 INVxp33_ASAP7_75t_R g217372 (.A(n_3173),
    .Y(n_3174));
 INVxp67_ASAP7_75t_R g217373 (.A(n_3171),
    .Y(n_3172));
 INVxp33_ASAP7_75t_R g217374 (.A(n_3165),
    .Y(n_3166));
 INVxp33_ASAP7_75t_R g217375 (.A(n_3161),
    .Y(n_3162));
 INVxp67_ASAP7_75t_R g217376 (.A(n_3152),
    .Y(n_3153));
 INVxp33_ASAP7_75t_R g217377 (.A(n_3150),
    .Y(n_3151));
 INVxp33_ASAP7_75t_R g217378 (.A(n_3147),
    .Y(n_3148));
 INVxp67_ASAP7_75t_R g217379 (.A(n_3144),
    .Y(n_3145));
 INVxp33_ASAP7_75t_R g217380 (.A(n_3139),
    .Y(n_3140));
 INVxp33_ASAP7_75t_R g217381 (.A(n_3137),
    .Y(n_3138));
 INVxp33_ASAP7_75t_R g217382 (.A(n_3132),
    .Y(n_3133));
 INVxp33_ASAP7_75t_R g217383 (.A(n_3130),
    .Y(n_3131));
 INVxp67_ASAP7_75t_R g217384 (.A(n_3125),
    .Y(n_3126));
 INVxp33_ASAP7_75t_R g217385 (.A(n_3122),
    .Y(n_3123));
 INVxp33_ASAP7_75t_R g217386 (.A(n_3119),
    .Y(n_3120));
 INVxp33_ASAP7_75t_R g217387 (.A(n_3113),
    .Y(n_3114));
 INVxp67_ASAP7_75t_R g217388 (.A(n_3108),
    .Y(n_3109));
 INVxp33_ASAP7_75t_R g217389 (.A(n_3106),
    .Y(n_3107));
 INVxp33_ASAP7_75t_R g217390 (.A(n_3104),
    .Y(n_3105));
 INVxp33_ASAP7_75t_R g217391 (.A(n_3101),
    .Y(n_3102));
 INVxp67_ASAP7_75t_R g217392 (.A(n_3099),
    .Y(n_3100));
 INVxp33_ASAP7_75t_R g217393 (.A(n_3095),
    .Y(n_3096));
 INVxp33_ASAP7_75t_R g217394 (.A(n_3091),
    .Y(n_3092));
 INVxp67_ASAP7_75t_R g217395 (.A(n_3087),
    .Y(n_3086));
 INVxp67_ASAP7_75t_R g217396 (.A(n_3083),
    .Y(n_3082));
 INVxp67_ASAP7_75t_R g217397 (.A(n_3080),
    .Y(n_3081));
 INVxp67_ASAP7_75t_L g217398 (.A(n_3074),
    .Y(n_3075));
 INVxp67_ASAP7_75t_R g217399 (.A(n_3072),
    .Y(n_3073));
 INVxp67_ASAP7_75t_R g217400 (.A(n_3070),
    .Y(n_3071));
 INVxp33_ASAP7_75t_R g217401 (.A(n_3067),
    .Y(n_3068));
 INVx1_ASAP7_75t_L g217402 (.A(n_3066),
    .Y(n_3065));
 INVxp67_ASAP7_75t_R g217404 (.A(n_3051),
    .Y(n_3052));
 INVxp67_ASAP7_75t_R g217405 (.A(n_3049),
    .Y(n_3050));
 INVxp33_ASAP7_75t_R g217406 (.A(n_3047),
    .Y(n_3048));
 INVxp67_ASAP7_75t_L g217407 (.A(n_3044),
    .Y(n_3043));
 INVxp33_ASAP7_75t_R g217408 (.A(n_3041),
    .Y(n_3042));
 INVxp33_ASAP7_75t_R g217409 (.A(n_3039),
    .Y(n_3040));
 INVxp33_ASAP7_75t_R g217410 (.A(n_3027),
    .Y(n_3028));
 INVxp33_ASAP7_75t_R g217411 (.A(n_3022),
    .Y(n_3021));
 INVxp67_ASAP7_75t_R g217412 (.A(n_3019),
    .Y(n_3018));
 INVxp33_ASAP7_75t_R g217413 (.A(n_3014),
    .Y(n_3013));
 INVxp67_ASAP7_75t_R g217414 (.A(n_3009),
    .Y(n_3010));
 INVx1_ASAP7_75t_L g217415 (.A(n_3006),
    .Y(n_3007));
 INVxp33_ASAP7_75t_R g217416 (.A(n_3005),
    .Y(n_3004));
 INVxp33_ASAP7_75t_R g217417 (.A(n_2999),
    .Y(n_3000));
 INVxp67_ASAP7_75t_R g217418 (.A(n_2997),
    .Y(n_2998));
 INVxp67_ASAP7_75t_R g217419 (.A(n_2995),
    .Y(n_2996));
 INVxp67_ASAP7_75t_L g217422 (.A(n_2989),
    .Y(n_2990));
 INVxp33_ASAP7_75t_R g217423 (.A(n_2985),
    .Y(n_2986));
 INVxp33_ASAP7_75t_R g217424 (.A(n_2982),
    .Y(n_2983));
 INVxp67_ASAP7_75t_R g217425 (.A(n_2980),
    .Y(n_2981));
 INVxp67_ASAP7_75t_R g217426 (.A(n_2977),
    .Y(n_2978));
 INVxp67_ASAP7_75t_R g217428 (.A(n_2975),
    .Y(n_2974));
 INVxp67_ASAP7_75t_R g217429 (.A(n_2971),
    .Y(n_2972));
 INVxp33_ASAP7_75t_R g217430 (.A(n_2969),
    .Y(n_2970));
 INVxp67_ASAP7_75t_R g217431 (.A(n_2968),
    .Y(n_2967));
 INVxp33_ASAP7_75t_R g217432 (.A(n_2965),
    .Y(n_2966));
 INVxp33_ASAP7_75t_R g217433 (.A(n_2963),
    .Y(n_2964));
 INVxp67_ASAP7_75t_R g217434 (.A(n_2959),
    .Y(n_2958));
 INVxp67_ASAP7_75t_R g217435 (.A(n_2951),
    .Y(n_2952));
 INVxp33_ASAP7_75t_R g217436 (.A(n_2949),
    .Y(n_2950));
 INVxp67_ASAP7_75t_R g217437 (.A(n_2947),
    .Y(n_2948));
 INVxp33_ASAP7_75t_R g217438 (.A(n_2945),
    .Y(n_2944));
 INVxp33_ASAP7_75t_R g217439 (.A(n_2941),
    .Y(n_2942));
 INVxp67_ASAP7_75t_R g217441 (.A(n_1722),
    .Y(n_2939));
 INVxp67_ASAP7_75t_SL g217444 (.A(n_2933),
    .Y(n_2932));
 INVxp67_ASAP7_75t_L g217445 (.A(n_2929),
    .Y(n_2928));
 INVxp33_ASAP7_75t_R g217446 (.A(n_2927),
    .Y(n_2926));
 INVx1_ASAP7_75t_R g217447 (.A(n_2924),
    .Y(n_2925));
 INVxp33_ASAP7_75t_R g217448 (.A(n_2922),
    .Y(n_2923));
 INVx1_ASAP7_75t_R g217449 (.A(n_2921),
    .Y(n_2920));
 INVx1_ASAP7_75t_L g217451 (.A(n_2916),
    .Y(n_2915));
 INVxp67_ASAP7_75t_SL g217452 (.A(n_2914),
    .Y(n_2913));
 INVx1_ASAP7_75t_SL g217453 (.A(n_2912),
    .Y(n_2911));
 INVxp67_ASAP7_75t_R g217454 (.A(n_2910),
    .Y(n_2909));
 INVxp67_ASAP7_75t_R g217455 (.A(n_2908),
    .Y(n_2907));
 INVx1_ASAP7_75t_R g217456 (.A(n_2905),
    .Y(n_2906));
 INVx1_ASAP7_75t_SL g217457 (.A(n_2903),
    .Y(n_2904));
 INVx1_ASAP7_75t_L g217458 (.A(n_2902),
    .Y(n_2901));
 INVxp67_ASAP7_75t_L g217459 (.A(n_2899),
    .Y(n_2898));
 INVx1_ASAP7_75t_R g217460 (.A(n_2897),
    .Y(n_2896));
 INVx1_ASAP7_75t_L g217461 (.A(n_2894),
    .Y(n_2895));
 INVx2_ASAP7_75t_L g217462 (.A(n_2893),
    .Y(n_2892));
 INVx1_ASAP7_75t_R g217463 (.A(n_2890),
    .Y(n_2891));
 INVxp67_ASAP7_75t_R g217464 (.A(n_2889),
    .Y(n_2888));
 INVx1_ASAP7_75t_L g217465 (.A(n_2887),
    .Y(n_2886));
 INVx1_ASAP7_75t_L g217466 (.A(n_2884),
    .Y(n_2883));
 INVxp67_ASAP7_75t_R g217467 (.A(n_2882),
    .Y(n_2881));
 INVxp67_ASAP7_75t_R g217470 (.A(n_2880),
    .Y(n_1719));
 INVxp67_ASAP7_75t_R g217471 (.A(n_1720),
    .Y(n_2880));
 INVxp33_ASAP7_75t_L g217472 (.A(n_2878),
    .Y(n_2877));
 INVxp33_ASAP7_75t_R g217474 (.A(n_1718),
    .Y(n_2876));
 INVxp67_ASAP7_75t_L g217476 (.A(n_2875),
    .Y(n_2874));
 INVx1_ASAP7_75t_L g217477 (.A(n_2873),
    .Y(n_2872));
 INVx1_ASAP7_75t_SL g217478 (.A(n_2871),
    .Y(n_2870));
 INVx1_ASAP7_75t_L g217479 (.A(n_2869),
    .Y(n_2868));
 INVxp67_ASAP7_75t_R g217480 (.A(n_2867),
    .Y(n_2866));
 INVx1_ASAP7_75t_L g217481 (.A(n_2864),
    .Y(n_2865));
 INVxp67_ASAP7_75t_SL g217482 (.A(n_2863),
    .Y(n_2862));
 INVx1_ASAP7_75t_SL g217485 (.A(n_1717),
    .Y(n_1716));
 INVx1_ASAP7_75t_L g217486 (.A(n_2861),
    .Y(n_1717));
 INVxp33_ASAP7_75t_R g217487 (.A(n_2860),
    .Y(n_2859));
 INVxp67_ASAP7_75t_R g217488 (.A(n_2858),
    .Y(n_2857));
 INVxp67_ASAP7_75t_R g217489 (.A(n_1715),
    .Y(n_2855));
 INVx2_ASAP7_75t_SL g217493 (.A(n_2854),
    .Y(n_2853));
 INVx2_ASAP7_75t_L g217494 (.A(n_2852),
    .Y(n_2851));
 INVxp67_ASAP7_75t_R g217495 (.A(n_2850),
    .Y(n_2849));
 INVx1_ASAP7_75t_L g217496 (.A(n_2848),
    .Y(n_2847));
 INVx2_ASAP7_75t_R g217497 (.A(n_2846),
    .Y(n_2845));
 INVxp67_ASAP7_75t_R g217498 (.A(n_2844),
    .Y(n_2843));
 INVxp33_ASAP7_75t_R g217499 (.A(n_2842),
    .Y(n_2841));
 INVx1_ASAP7_75t_L g217500 (.A(n_2840),
    .Y(n_2839));
 INVx1_ASAP7_75t_L g217501 (.A(n_2838),
    .Y(n_2837));
 INVx1_ASAP7_75t_SL g217503 (.A(n_2834),
    .Y(n_2835));
 INVxp67_ASAP7_75t_L g217506 (.A(n_2833),
    .Y(n_2832));
 INVx1_ASAP7_75t_R g217507 (.A(n_2831),
    .Y(n_2830));
 INVxp67_ASAP7_75t_R g217508 (.A(n_2829),
    .Y(n_2828));
 INVx1_ASAP7_75t_L g217509 (.A(n_2827),
    .Y(n_2826));
 INVxp33_ASAP7_75t_R g217510 (.A(n_2825),
    .Y(n_2824));
 INVxp67_ASAP7_75t_L g217511 (.A(n_2823),
    .Y(n_2822));
 INVx2_ASAP7_75t_SL g217512 (.A(n_2821),
    .Y(n_2820));
 INVx2_ASAP7_75t_L g217513 (.A(n_2819),
    .Y(n_2818));
 INVx1_ASAP7_75t_SL g217514 (.A(n_2817),
    .Y(n_2816));
 INVx2_ASAP7_75t_SL g217515 (.A(n_2815),
    .Y(n_2814));
 INVxp67_ASAP7_75t_R g217517 (.A(n_1714),
    .Y(n_2813));
 INVx2_ASAP7_75t_L g217520 (.A(n_1713),
    .Y(n_1714));
 INVx1_ASAP7_75t_R g217523 (.A(n_2811),
    .Y(n_1712));
 INVxp67_ASAP7_75t_L g217525 (.A(n_2808),
    .Y(n_2809));
 INVx2_ASAP7_75t_SL g217526 (.A(n_2811),
    .Y(n_2808));
 INVx1_ASAP7_75t_SL g217527 (.A(n_2807),
    .Y(n_2806));
 INVx1_ASAP7_75t_R g217528 (.A(n_2805),
    .Y(n_2804));
 INVx2_ASAP7_75t_SL g217529 (.A(n_2803),
    .Y(n_2802));
 INVx1_ASAP7_75t_L g217530 (.A(n_2800),
    .Y(n_2801));
 BUFx3_ASAP7_75t_SL g217535 (.A(n_2798),
    .Y(n_2800));
 INVx1_ASAP7_75t_L g217536 (.A(n_2798),
    .Y(n_2799));
 INVxp67_ASAP7_75t_R g217537 (.A(n_2797),
    .Y(n_2796));
 INVxp33_ASAP7_75t_R g217538 (.A(n_1711),
    .Y(n_2795));
 INVx2_ASAP7_75t_SL g217541 (.A(n_2794),
    .Y(n_1710));
 INVx1_ASAP7_75t_L g217542 (.A(n_1710),
    .Y(n_1711));
 INVx1_ASAP7_75t_SL g217544 (.A(n_2793),
    .Y(n_2792));
 INVx2_ASAP7_75t_L g217546 (.A(n_2790),
    .Y(n_2789));
 INVx2_ASAP7_75t_SL g217547 (.A(n_2791),
    .Y(n_2790));
 INVx1_ASAP7_75t_L g217550 (.A(n_2788),
    .Y(n_2787));
 INVx1_ASAP7_75t_R g217551 (.A(n_2786),
    .Y(n_2785));
 INVx5_ASAP7_75t_SL g217552 (.A(n_2784),
    .Y(n_2783));
 INVx1_ASAP7_75t_R g217553 (.A(n_2782),
    .Y(n_2781));
 INVx2_ASAP7_75t_SL g217554 (.A(n_2780),
    .Y(n_2779));
 INVx2_ASAP7_75t_L g217555 (.A(n_2778),
    .Y(n_2777));
 XNOR2xp5_ASAP7_75t_R g217556 (.A(w3[14]),
    .B(text_in_r[14]),
    .Y(n_2776));
 XNOR2xp5_ASAP7_75t_R g217557 (.A(w0[14]),
    .B(text_in_r[110]),
    .Y(n_2775));
 XNOR2xp5_ASAP7_75t_R g217558 (.A(w0[18]),
    .B(text_in_r[114]),
    .Y(n_2774));
 NOR3xp33_ASAP7_75t_R g217559 (.A(n_2158),
    .B(n_1499),
    .C(n_1491),
    .Y(n_2773));
 NAND2xp33_ASAP7_75t_R g217560 (.A(n_2173),
    .B(n_1633),
    .Y(n_2772));
 NAND2xp33_ASAP7_75t_R g217561 (.A(n_1603),
    .B(n_8690),
    .Y(n_2771));
 NOR2xp33_ASAP7_75t_R g217562 (.A(n_2173),
    .B(n_1642),
    .Y(n_2770));
 NAND2xp33_ASAP7_75t_R g217563 (.A(n_2168),
    .B(n_1625),
    .Y(n_2769));
 NOR2xp33_ASAP7_75t_R g217564 (.A(n_2231),
    .B(n_1369),
    .Y(n_2768));
 NAND2xp33_ASAP7_75t_R g217565 (.A(n_2141),
    .B(n_2427),
    .Y(n_2767));
 NOR2xp33_ASAP7_75t_R g217566 (.A(n_2187),
    .B(n_1662),
    .Y(n_2766));
 NAND2xp5_ASAP7_75t_R g217567 (.A(n_2235),
    .B(n_2075),
    .Y(n_2765));
 NAND2xp33_ASAP7_75t_R g217568 (.A(n_1601),
    .B(n_2353),
    .Y(n_2764));
 NAND2xp33_ASAP7_75t_R g217569 (.A(n_2253),
    .B(n_1545),
    .Y(n_2763));
 NAND2xp33_ASAP7_75t_L g217570 (.A(n_2134),
    .B(n_2347),
    .Y(n_2762));
 NAND2xp33_ASAP7_75t_R g217571 (.A(n_2394),
    .B(n_2212),
    .Y(n_2761));
 NAND2xp33_ASAP7_75t_R g217572 (.A(n_2436),
    .B(n_1552),
    .Y(n_2760));
 NOR2xp33_ASAP7_75t_R g217573 (.A(n_2056),
    .B(n_2468),
    .Y(n_2759));
 NAND2xp33_ASAP7_75t_R g217574 (.A(n_1448),
    .B(n_2442),
    .Y(n_2758));
 NAND2xp33_ASAP7_75t_R g217575 (.A(n_1592),
    .B(n_2467),
    .Y(n_2757));
 NAND2xp33_ASAP7_75t_R g217576 (.A(n_1678),
    .B(n_1446),
    .Y(n_2756));
 NAND2xp5_ASAP7_75t_L g217577 (.A(n_2445),
    .B(n_1432),
    .Y(n_2755));
 NAND2xp33_ASAP7_75t_R g217578 (.A(n_2447),
    .B(n_1668),
    .Y(n_2754));
 NAND2xp33_ASAP7_75t_L g217579 (.A(n_2523),
    .B(n_2475),
    .Y(n_2753));
 NAND2xp33_ASAP7_75t_R g217580 (.A(n_2519),
    .B(n_2107),
    .Y(n_3219));
 NAND2xp33_ASAP7_75t_R g217581 (.A(n_2484),
    .B(n_1647),
    .Y(n_2752));
 NAND2xp33_ASAP7_75t_R g217582 (.A(n_2552),
    .B(n_1623),
    .Y(n_2751));
 NAND2xp33_ASAP7_75t_R g217583 (.A(n_2548),
    .B(n_1398),
    .Y(n_2750));
 NAND2xp33_ASAP7_75t_R g217584 (.A(n_1673),
    .B(n_2215),
    .Y(n_2749));
 NAND2xp33_ASAP7_75t_R g217585 (.A(n_2508),
    .B(n_2192),
    .Y(n_2748));
 NOR2xp33_ASAP7_75t_R g217586 (.A(n_2104),
    .B(n_2532),
    .Y(n_2747));
 NOR2xp33_ASAP7_75t_L g217587 (.A(n_1498),
    .B(n_2158),
    .Y(n_2746));
 NOR2xp33_ASAP7_75t_R g217588 (.A(n_2550),
    .B(n_2393),
    .Y(n_2745));
 NAND2xp33_ASAP7_75t_R g217589 (.A(n_2550),
    .B(n_2420),
    .Y(n_2744));
 NOR2xp33_ASAP7_75t_R g217590 (.A(n_2170),
    .B(n_1690),
    .Y(n_2743));
 NOR2xp33_ASAP7_75t_R g217591 (.A(n_2102),
    .B(n_2572),
    .Y(n_2742));
 NOR2xp33_ASAP7_75t_L g217592 (.A(n_2590),
    .B(n_2419),
    .Y(n_2741));
 NOR2xp33_ASAP7_75t_L g217593 (.A(n_1941),
    .B(n_2460),
    .Y(n_2740));
 NOR2xp33_ASAP7_75t_L g217594 (.A(n_1427),
    .B(n_2445),
    .Y(n_2739));
 NAND2xp33_ASAP7_75t_R g217595 (.A(n_2634),
    .B(n_2044),
    .Y(n_2738));
 NAND2xp33_ASAP7_75t_R g217596 (.A(n_2135),
    .B(n_2475),
    .Y(n_3217));
 NOR2xp33_ASAP7_75t_R g217597 (.A(n_1506),
    .B(n_1615),
    .Y(n_3216));
 NOR2xp33_ASAP7_75t_R g217598 (.A(n_2175),
    .B(n_2080),
    .Y(n_3215));
 NOR2xp33_ASAP7_75t_SL g217599 (.A(n_1852),
    .B(n_2147),
    .Y(n_3213));
 NAND2xp5_ASAP7_75t_R g217600 (.A(n_8200),
    .B(n_1614),
    .Y(n_3212));
 NOR2xp33_ASAP7_75t_L g217601 (.A(n_1387),
    .B(n_1616),
    .Y(n_3211));
 NOR2xp33_ASAP7_75t_R g217602 (.A(sa31[4]),
    .B(n_2291),
    .Y(n_3210));
 NOR2xp33_ASAP7_75t_SL g217603 (.A(n_1567),
    .B(n_2302),
    .Y(n_3209));
 NOR2xp33_ASAP7_75t_L g217604 (.A(n_2281),
    .B(n_1651),
    .Y(n_3208));
 NOR2xp33_ASAP7_75t_R g217605 (.A(n_1360),
    .B(n_2286),
    .Y(n_3207));
 NOR2xp33_ASAP7_75t_SL g217606 (.A(n_2227),
    .B(n_2044),
    .Y(n_3206));
 NOR2xp33_ASAP7_75t_L g217607 (.A(n_2299),
    .B(n_2423),
    .Y(n_3205));
 NAND2xp5_ASAP7_75t_R g217608 (.A(n_1664),
    .B(n_2307),
    .Y(n_3204));
 NOR2xp33_ASAP7_75t_R g217609 (.A(n_2310),
    .B(n_2053),
    .Y(n_3203));
 NAND2xp5_ASAP7_75t_R g217610 (.A(n_2301),
    .B(n_1561),
    .Y(n_3202));
 NOR2xp33_ASAP7_75t_R g217611 (.A(n_2428),
    .B(n_2310),
    .Y(n_3201));
 NAND2xp5_ASAP7_75t_L g217612 (.A(n_1677),
    .B(n_2475),
    .Y(n_3199));
 NAND2xp5_ASAP7_75t_L g217613 (.A(n_8896),
    .B(n_2115),
    .Y(n_3198));
 NOR2xp33_ASAP7_75t_R g217614 (.A(n_1383),
    .B(n_2293),
    .Y(n_2737));
 NAND2xp33_ASAP7_75t_R g217615 (.A(n_2043),
    .B(n_2270),
    .Y(n_3197));
 NAND2xp5_ASAP7_75t_R g217616 (.A(n_2312),
    .B(n_2425),
    .Y(n_3196));
 NAND2xp5_ASAP7_75t_R g217617 (.A(n_2330),
    .B(n_1657),
    .Y(n_3195));
 NAND2xp5_ASAP7_75t_R g217618 (.A(n_2316),
    .B(n_1406),
    .Y(n_3194));
 NAND2xp5_ASAP7_75t_R g217619 (.A(n_2324),
    .B(n_2385),
    .Y(n_3193));
 NAND2xp5_ASAP7_75t_R g217620 (.A(n_2312),
    .B(n_1545),
    .Y(n_3191));
 NOR2xp33_ASAP7_75t_R g217621 (.A(n_2296),
    .B(n_1635),
    .Y(n_3190));
 NAND2xp33_ASAP7_75t_R g217622 (.A(n_2278),
    .B(n_8189),
    .Y(n_3189));
 NOR2xp33_ASAP7_75t_L g217623 (.A(n_2323),
    .B(n_2043),
    .Y(n_3187));
 NOR2xp33_ASAP7_75t_L g217624 (.A(n_1364),
    .B(n_2306),
    .Y(n_3186));
 NOR2xp33_ASAP7_75t_L g217625 (.A(n_1646),
    .B(n_2304),
    .Y(n_2736));
 NOR2xp33_ASAP7_75t_L g217626 (.A(n_1669),
    .B(n_2332),
    .Y(n_3185));
 NOR2xp33_ASAP7_75t_SL g217627 (.A(n_2111),
    .B(n_1665),
    .Y(n_3184));
 NAND2xp5_ASAP7_75t_R g217628 (.A(n_2303),
    .B(n_2062),
    .Y(n_3183));
 NOR2xp33_ASAP7_75t_R g217629 (.A(n_1425),
    .B(n_2325),
    .Y(n_3182));
 NOR2xp33_ASAP7_75t_R g217630 (.A(n_2332),
    .B(n_2057),
    .Y(n_3180));
 NOR2xp33_ASAP7_75t_R g217631 (.A(n_1375),
    .B(n_1620),
    .Y(n_3179));
 NAND2xp5_ASAP7_75t_R g217632 (.A(n_2136),
    .B(n_2450),
    .Y(n_3177));
 NOR2xp33_ASAP7_75t_R g217633 (.A(n_1949),
    .B(n_1598),
    .Y(n_3175));
 NOR2xp33_ASAP7_75t_SL g217634 (.A(n_2468),
    .B(n_2418),
    .Y(n_3173));
 NAND2xp5_ASAP7_75t_R g217635 (.A(n_1680),
    .B(n_2483),
    .Y(n_3171));
 NAND2xp5_ASAP7_75t_R g217636 (.A(n_2153),
    .B(n_2442),
    .Y(n_3170));
 NAND2xp5_ASAP7_75t_R g217637 (.A(n_2436),
    .B(n_2488),
    .Y(n_3169));
 NOR2xp33_ASAP7_75t_R g217638 (.A(n_2199),
    .B(n_2484),
    .Y(n_3168));
 NOR2xp33_ASAP7_75t_R g217639 (.A(n_2123),
    .B(n_2438),
    .Y(n_3167));
 NAND2xp5_ASAP7_75t_R g217640 (.A(n_2473),
    .B(n_1659),
    .Y(n_3165));
 AND2x2_ASAP7_75t_R g217641 (.A(n_2481),
    .B(n_1351),
    .Y(n_3164));
 NOR2xp33_ASAP7_75t_R g217642 (.A(n_2438),
    .B(n_2129),
    .Y(n_3163));
 NOR2xp33_ASAP7_75t_L g217643 (.A(n_1599),
    .B(n_2478),
    .Y(n_3161));
 NAND2xp5_ASAP7_75t_R g217644 (.A(n_2485),
    .B(n_1597),
    .Y(n_3160));
 NOR2xp33_ASAP7_75t_SL g217645 (.A(n_1644),
    .B(n_2486),
    .Y(n_3159));
 NOR2xp33_ASAP7_75t_L g217646 (.A(n_1503),
    .B(n_2314),
    .Y(n_3158));
 NAND2xp33_ASAP7_75t_R g217647 (.A(n_1852),
    .B(n_2084),
    .Y(n_3157));
 NOR2xp33_ASAP7_75t_R g217648 (.A(n_2106),
    .B(n_2453),
    .Y(n_3156));
 NOR2xp33_ASAP7_75t_L g217649 (.A(sa12[4]),
    .B(n_2319),
    .Y(n_3155));
 NAND2xp5_ASAP7_75t_L g217650 (.A(n_1503),
    .B(n_2134),
    .Y(n_3154));
 NAND2xp5_ASAP7_75t_R g217651 (.A(n_2456),
    .B(n_2186),
    .Y(n_3152));
 NAND2xp5_ASAP7_75t_R g217652 (.A(n_1675),
    .B(n_2450),
    .Y(n_3150));
 NOR2xp33_ASAP7_75t_R g217653 (.A(n_2453),
    .B(n_2217),
    .Y(n_3149));
 NAND2xp33_ASAP7_75t_R g217654 (.A(n_2439),
    .B(n_2464),
    .Y(n_3147));
 NAND2xp5_ASAP7_75t_R g217655 (.A(n_2496),
    .B(n_2067),
    .Y(n_3146));
 NAND2xp5_ASAP7_75t_R g217656 (.A(n_2116),
    .B(n_2448),
    .Y(n_3144));
 NOR2xp33_ASAP7_75t_L g217657 (.A(n_1678),
    .B(n_2311),
    .Y(n_3143));
 NOR2xp33_ASAP7_75t_L g217658 (.A(n_2588),
    .B(n_1378),
    .Y(n_3142));
 NOR2xp33_ASAP7_75t_R g217659 (.A(n_1935),
    .B(n_2437),
    .Y(n_3141));
 NAND2xp5_ASAP7_75t_R g217660 (.A(n_1673),
    .B(n_2477),
    .Y(n_3139));
 NOR2xp33_ASAP7_75t_R g217661 (.A(n_2463),
    .B(n_2482),
    .Y(n_3137));
 NAND2xp5_ASAP7_75t_R g217662 (.A(n_2578),
    .B(n_1606),
    .Y(n_3136));
 NAND2xp33_ASAP7_75t_R g217663 (.A(n_2583),
    .B(n_1448),
    .Y(n_3135));
 NOR2xp33_ASAP7_75t_R g217664 (.A(n_2576),
    .B(n_1583),
    .Y(n_3134));
 AND2x2_ASAP7_75t_R g217665 (.A(n_2568),
    .B(n_2040),
    .Y(n_3132));
 NOR2xp33_ASAP7_75t_R g217666 (.A(n_2562),
    .B(n_2045),
    .Y(n_3130));
 NOR2xp33_ASAP7_75t_R g217667 (.A(n_2489),
    .B(n_2590),
    .Y(n_2735));
 NOR2xp33_ASAP7_75t_L g217668 (.A(n_2472),
    .B(n_2591),
    .Y(n_2734));
 NAND2xp33_ASAP7_75t_R g217669 (.A(n_2593),
    .B(n_2092),
    .Y(n_3129));
 NOR2xp33_ASAP7_75t_L g217670 (.A(n_2530),
    .B(n_1560),
    .Y(n_3128));
 NAND2xp5_ASAP7_75t_R g217671 (.A(n_1687),
    .B(n_2604),
    .Y(n_2733));
 NAND2xp5_ASAP7_75t_L g217672 (.A(n_2282),
    .B(n_2462),
    .Y(n_3127));
 NAND2xp33_ASAP7_75t_R g217673 (.A(n_2471),
    .B(n_2473),
    .Y(n_3125));
 NAND2xp5_ASAP7_75t_R g217674 (.A(n_2500),
    .B(n_2613),
    .Y(n_3124));
 NAND2xp33_ASAP7_75t_R g217675 (.A(n_2062),
    .B(n_2540),
    .Y(n_3122));
 NOR2xp33_ASAP7_75t_R g217676 (.A(n_2506),
    .B(n_2041),
    .Y(n_3121));
 NOR2xp33_ASAP7_75t_R g217677 (.A(n_2515),
    .B(n_2470),
    .Y(n_3119));
 NAND2xp33_ASAP7_75t_R g217678 (.A(n_2132),
    .B(n_2481),
    .Y(n_3118));
 NOR2xp33_ASAP7_75t_R g217679 (.A(n_2131),
    .B(n_2457),
    .Y(n_3117));
 NAND2xp33_ASAP7_75t_R g217680 (.A(n_2065),
    .B(n_2456),
    .Y(n_3116));
 NAND2xp5_ASAP7_75t_R g217681 (.A(n_1673),
    .B(n_2324),
    .Y(n_3115));
 NAND2xp33_ASAP7_75t_R g217682 (.A(n_2502),
    .B(n_2054),
    .Y(n_3113));
 NAND2xp33_ASAP7_75t_R g217683 (.A(n_2062),
    .B(n_2539),
    .Y(n_3112));
 NAND2xp5_ASAP7_75t_L g217684 (.A(n_2521),
    .B(n_2435),
    .Y(n_3111));
 NAND2xp33_ASAP7_75t_R g217685 (.A(n_2443),
    .B(n_2389),
    .Y(n_3110));
 NAND2xp5_ASAP7_75t_R g217686 (.A(n_2448),
    .B(n_1349),
    .Y(n_3108));
 NOR2xp33_ASAP7_75t_L g217687 (.A(n_2138),
    .B(n_2470),
    .Y(n_3106));
 NOR2xp33_ASAP7_75t_R g217688 (.A(n_2451),
    .B(n_2175),
    .Y(n_3104));
 NAND2xp5_ASAP7_75t_R g217689 (.A(n_2440),
    .B(n_2140),
    .Y(n_3103));
 NAND2xp5_ASAP7_75t_R g217690 (.A(n_2436),
    .B(n_2211),
    .Y(n_3101));
 NOR2xp33_ASAP7_75t_L g217691 (.A(n_2492),
    .B(n_2310),
    .Y(n_3099));
 NOR2xp33_ASAP7_75t_L g217692 (.A(n_2438),
    .B(n_2434),
    .Y(n_3098));
 NOR2xp33_ASAP7_75t_R g217693 (.A(n_2143),
    .B(n_2476),
    .Y(n_3097));
 NOR2xp33_ASAP7_75t_L g217694 (.A(n_2495),
    .B(n_2302),
    .Y(n_3095));
 NOR2xp33_ASAP7_75t_R g217695 (.A(n_1601),
    .B(n_2441),
    .Y(n_3094));
 NAND2xp5_ASAP7_75t_L g217696 (.A(n_1345),
    .B(n_2331),
    .Y(n_3093));
 NAND2xp5_ASAP7_75t_L g217697 (.A(n_1613),
    .B(n_2508),
    .Y(n_3091));
 NOR2xp33_ASAP7_75t_R g217698 (.A(n_2158),
    .B(n_2449),
    .Y(n_2732));
 NOR2xp33_ASAP7_75t_R g217699 (.A(n_2470),
    .B(n_2194),
    .Y(n_3090));
 NAND2xp5_ASAP7_75t_R g217700 (.A(n_2509),
    .B(n_2076),
    .Y(n_3089));
 NOR2xp33_ASAP7_75t_R g217701 (.A(n_1679),
    .B(n_2304),
    .Y(n_3088));
 NOR2xp33_ASAP7_75t_L g217702 (.A(n_2066),
    .B(n_2511),
    .Y(n_3087));
 NAND2xp5_ASAP7_75t_R g217703 (.A(n_2512),
    .B(n_2385),
    .Y(n_3085));
 AND2x2_ASAP7_75t_L g217704 (.A(n_2583),
    .B(n_2442),
    .Y(n_3084));
 AND2x2_ASAP7_75t_L g217705 (.A(n_1385),
    .B(n_2154),
    .Y(n_3083));
 NOR2xp33_ASAP7_75t_L g217706 (.A(n_2507),
    .B(n_2411),
    .Y(n_3080));
 NAND2xp5_ASAP7_75t_R g217707 (.A(n_2127),
    .B(n_2466),
    .Y(n_3079));
 NAND2xp5_ASAP7_75t_R g217708 (.A(n_2585),
    .B(n_2055),
    .Y(n_3078));
 AND2x2_ASAP7_75t_L g217709 (.A(n_2094),
    .B(n_8690),
    .Y(n_3077));
 NAND2xp5_ASAP7_75t_L g217710 (.A(n_2537),
    .B(n_2619),
    .Y(n_3076));
 NOR2xp33_ASAP7_75t_L g217711 (.A(n_2555),
    .B(n_2043),
    .Y(n_3074));
 NAND2xp5_ASAP7_75t_R g217712 (.A(n_2094),
    .B(n_2413),
    .Y(n_3072));
 NOR2xp33_ASAP7_75t_R g217713 (.A(n_2214),
    .B(n_2043),
    .Y(n_3070));
 NAND2xp5_ASAP7_75t_R g217714 (.A(n_2060),
    .B(n_2553),
    .Y(n_3069));
 NAND2xp33_ASAP7_75t_R g217715 (.A(sa12[4]),
    .B(n_2133),
    .Y(n_3067));
 OR2x2_ASAP7_75t_SL g217716 (.A(n_2510),
    .B(n_1651),
    .Y(n_3066));
 NOR2x1_ASAP7_75t_L g217717 (.A(n_2252),
    .B(n_1678),
    .Y(n_3064));
 NOR2xp33_ASAP7_75t_R g217718 (.A(n_2576),
    .B(n_2482),
    .Y(n_3063));
 NOR2xp33_ASAP7_75t_SL g217719 (.A(n_1359),
    .B(n_2122),
    .Y(n_3062));
 NAND2xp33_ASAP7_75t_R g217720 (.A(n_2571),
    .B(n_2062),
    .Y(n_3061));
 NAND2xp5_ASAP7_75t_R g217721 (.A(n_2503),
    .B(n_2420),
    .Y(n_3060));
 NAND2xp5_ASAP7_75t_R g217722 (.A(n_2496),
    .B(n_2435),
    .Y(n_3059));
 AND2x2_ASAP7_75t_SL g217723 (.A(n_2585),
    .B(n_2467),
    .Y(n_3058));
 NOR2xp33_ASAP7_75t_L g217724 (.A(n_2474),
    .B(n_2562),
    .Y(n_3057));
 NAND2xp5_ASAP7_75t_SL g217725 (.A(n_1699),
    .B(n_2512),
    .Y(n_3056));
 NOR2x1_ASAP7_75t_L g217726 (.A(n_2567),
    .B(n_2486),
    .Y(n_3055));
 NOR2xp67_ASAP7_75t_SL g217727 (.A(n_1674),
    .B(n_2231),
    .Y(n_1725));
 NAND2xp5_ASAP7_75t_R g217728 (.A(n_2442),
    .B(n_2223),
    .Y(n_3054));
 NOR2xp33_ASAP7_75t_L g217729 (.A(n_2555),
    .B(n_2478),
    .Y(n_3053));
 NAND2xp5_ASAP7_75t_L g217730 (.A(n_2553),
    .B(n_2450),
    .Y(n_3051));
 NAND2xp5_ASAP7_75t_SL g217731 (.A(n_2448),
    .B(n_2529),
    .Y(n_3049));
 AND2x2_ASAP7_75t_L g217732 (.A(n_2197),
    .B(n_2076),
    .Y(n_3047));
 NOR2xp33_ASAP7_75t_L g217733 (.A(n_2299),
    .B(n_1674),
    .Y(n_3046));
 NAND2xp5_ASAP7_75t_R g217734 (.A(n_2119),
    .B(n_1542),
    .Y(n_3045));
 NOR2xp33_ASAP7_75t_L g217735 (.A(n_2465),
    .B(n_2293),
    .Y(n_3044));
 NOR2x1_ASAP7_75t_R g217736 (.A(n_2606),
    .B(n_1690),
    .Y(n_3041));
 NOR2xp67_ASAP7_75t_L g217737 (.A(n_2465),
    .B(n_2235),
    .Y(n_3039));
 AND2x2_ASAP7_75t_SL g217738 (.A(n_2486),
    .B(n_2383),
    .Y(n_3038));
 NOR2xp33_ASAP7_75t_R g217739 (.A(n_2522),
    .B(n_2068),
    .Y(n_3037));
 NAND2xp5_ASAP7_75t_L g217740 (.A(n_1673),
    .B(n_2169),
    .Y(n_3036));
 AND2x2_ASAP7_75t_L g217741 (.A(n_2455),
    .B(n_2268),
    .Y(n_3035));
 NAND2xp5_ASAP7_75t_SL g217742 (.A(n_2618),
    .B(n_2496),
    .Y(n_3034));
 NOR2xp33_ASAP7_75t_L g217743 (.A(n_2486),
    .B(n_2173),
    .Y(n_3033));
 NAND2xp5_ASAP7_75t_L g217744 (.A(n_2531),
    .B(n_2040),
    .Y(n_3032));
 AND2x2_ASAP7_75t_R g217745 (.A(n_2058),
    .B(n_1691),
    .Y(n_3031));
 NAND2xp5_ASAP7_75t_R g217746 (.A(n_1851),
    .B(n_2199),
    .Y(n_3030));
 NAND2xp5_ASAP7_75t_R g217747 (.A(n_2483),
    .B(n_2127),
    .Y(n_3029));
 NAND2xp5_ASAP7_75t_R g217748 (.A(n_1387),
    .B(n_2108),
    .Y(n_3027));
 AND2x2_ASAP7_75t_R g217749 (.A(n_2482),
    .B(n_1351),
    .Y(n_3026));
 NAND2xp5_ASAP7_75t_L g217750 (.A(n_2330),
    .B(n_2471),
    .Y(n_3025));
 NAND2xp5_ASAP7_75t_R g217751 (.A(n_2440),
    .B(n_2427),
    .Y(n_3024));
 NOR2xp33_ASAP7_75t_L g217752 (.A(n_2634),
    .B(n_2520),
    .Y(n_3023));
 NAND2xp5_ASAP7_75t_R g217753 (.A(n_2571),
    .B(n_2401),
    .Y(n_3022));
 NOR2x1_ASAP7_75t_R g217754 (.A(n_2539),
    .B(n_2484),
    .Y(n_3020));
 AND2x2_ASAP7_75t_L g217755 (.A(n_1557),
    .B(n_2457),
    .Y(n_3019));
 AND2x2_ASAP7_75t_R g217756 (.A(n_2534),
    .B(n_2054),
    .Y(n_3017));
 NOR2xp33_ASAP7_75t_L g217757 (.A(n_1688),
    .B(n_2209),
    .Y(n_3016));
 NAND2xp5_ASAP7_75t_L g217758 (.A(n_1687),
    .B(n_2290),
    .Y(n_3015));
 OR2x2_ASAP7_75t_L g217759 (.A(n_2472),
    .B(n_2227),
    .Y(n_3014));
 NAND2xp5_ASAP7_75t_L g217760 (.A(n_2525),
    .B(n_1552),
    .Y(n_3012));
 NAND2xp5_ASAP7_75t_R g217761 (.A(n_2484),
    .B(n_2416),
    .Y(n_3011));
 NAND2xp5_ASAP7_75t_R g217762 (.A(n_2523),
    .B(n_1542),
    .Y(n_3009));
 NAND2xp5_ASAP7_75t_R g217763 (.A(n_2503),
    .B(n_2060),
    .Y(n_3008));
 NAND2xp5_ASAP7_75t_L g217764 (.A(n_1561),
    .B(n_2537),
    .Y(n_3006));
 AND2x2_ASAP7_75t_R g217765 (.A(n_2441),
    .B(n_2397),
    .Y(n_3005));
 NAND2xp5_ASAP7_75t_R g217766 (.A(n_2536),
    .B(n_1705),
    .Y(n_3003));
 AND2x2_ASAP7_75t_R g217767 (.A(n_2476),
    .B(n_1350),
    .Y(n_3002));
 NOR2xp33_ASAP7_75t_R g217768 (.A(n_1386),
    .B(n_2328),
    .Y(n_3001));
 NAND2xp5_ASAP7_75t_L g217769 (.A(n_2196),
    .B(n_2462),
    .Y(n_2999));
 NAND2xp5_ASAP7_75t_R g217770 (.A(n_2534),
    .B(n_1704),
    .Y(n_2997));
 NOR2xp33_ASAP7_75t_R g217771 (.A(n_1361),
    .B(n_1592),
    .Y(n_2995));
 NAND2xp5_ASAP7_75t_SL g217772 (.A(n_2452),
    .B(n_2518),
    .Y(n_1724));
 NAND2xp5_ASAP7_75t_R g217773 (.A(n_2449),
    .B(n_1566),
    .Y(n_2994));
 NOR2xp33_ASAP7_75t_R g217774 (.A(n_2474),
    .B(n_2187),
    .Y(n_2993));
 NAND2xp5_ASAP7_75t_R g217775 (.A(n_1691),
    .B(n_2432),
    .Y(n_2992));
 NOR2xp33_ASAP7_75t_L g217776 (.A(n_2478),
    .B(n_2168),
    .Y(n_2991));
 NOR2xp33_ASAP7_75t_L g217777 (.A(n_2499),
    .B(n_2348),
    .Y(n_2989));
 OR2x2_ASAP7_75t_L g217778 (.A(n_2499),
    .B(n_2182),
    .Y(n_2988));
 NAND2xp5_ASAP7_75t_R g217779 (.A(n_2467),
    .B(n_2241),
    .Y(n_2987));
 AND2x2_ASAP7_75t_L g217780 (.A(n_2534),
    .B(n_2427),
    .Y(n_2985));
 NOR2xp33_ASAP7_75t_R g217781 (.A(n_1591),
    .B(n_1583),
    .Y(n_2984));
 NAND2xp5_ASAP7_75t_L g217782 (.A(n_1683),
    .B(n_2247),
    .Y(n_2982));
 NAND2xp5_ASAP7_75t_R g217783 (.A(n_2531),
    .B(n_1636),
    .Y(n_2980));
 NAND2xp5_ASAP7_75t_R g217784 (.A(n_1609),
    .B(n_2481),
    .Y(n_2979));
 NAND2xp5_ASAP7_75t_L g217785 (.A(n_1605),
    .B(n_2067),
    .Y(n_2977));
 AND2x2_ASAP7_75t_L g217786 (.A(n_1689),
    .B(n_2048),
    .Y(n_2976));
 NOR2xp67_ASAP7_75t_L g217787 (.A(n_2450),
    .B(n_2393),
    .Y(n_1723));
 NOR2xp33_ASAP7_75t_SL g217788 (.A(n_1665),
    .B(n_2526),
    .Y(n_2975));
 NOR2x1_ASAP7_75t_SL g217789 (.A(n_2487),
    .B(n_2213),
    .Y(n_2973));
 NOR2xp33_ASAP7_75t_L g217790 (.A(n_2487),
    .B(n_2308),
    .Y(n_2971));
 NOR2xp33_ASAP7_75t_R g217791 (.A(n_2495),
    .B(n_2249),
    .Y(n_2969));
 NAND2xp5_ASAP7_75t_L g217792 (.A(n_1349),
    .B(n_2537),
    .Y(n_2968));
 NAND2xp5_ASAP7_75t_L g217793 (.A(n_2490),
    .B(n_2254),
    .Y(n_2965));
 NAND2xp5_ASAP7_75t_L g217794 (.A(n_2316),
    .B(n_2490),
    .Y(n_2963));
 NAND2xp5_ASAP7_75t_L g217795 (.A(n_2438),
    .B(n_2400),
    .Y(n_2962));
 NAND2xp33_ASAP7_75t_R g217796 (.A(n_2436),
    .B(n_2092),
    .Y(n_2961));
 NOR2xp67_ASAP7_75t_L g217797 (.A(n_2588),
    .B(n_2457),
    .Y(n_2960));
 NOR2x1_ASAP7_75t_SL g217798 (.A(n_2447),
    .B(n_2256),
    .Y(n_2959));
 NAND2xp5_ASAP7_75t_L g217799 (.A(n_2478),
    .B(n_1445),
    .Y(n_2957));
 NAND2xp5_ASAP7_75t_R g217800 (.A(n_2297),
    .B(n_1682),
    .Y(n_2956));
 NOR2x1_ASAP7_75t_L g217801 (.A(n_2480),
    .B(n_2243),
    .Y(n_2955));
 NAND2xp5_ASAP7_75t_L g217802 (.A(n_1693),
    .B(n_2571),
    .Y(n_2954));
 NAND2xp5_ASAP7_75t_R g217803 (.A(n_2536),
    .B(n_2425),
    .Y(n_2953));
 NAND2xp5_ASAP7_75t_L g217804 (.A(n_2305),
    .B(n_2444),
    .Y(n_2951));
 NAND2xp5_ASAP7_75t_L g217805 (.A(n_2444),
    .B(n_2229),
    .Y(n_2949));
 NOR2xp33_ASAP7_75t_R g217806 (.A(n_2520),
    .B(n_1656),
    .Y(n_2947));
 NAND2xp5_ASAP7_75t_L g217807 (.A(n_2275),
    .B(n_2466),
    .Y(n_2946));
 NOR2xp33_ASAP7_75t_L g217808 (.A(n_1948),
    .B(n_2186),
    .Y(n_2945));
 AND2x2_ASAP7_75t_SL g217809 (.A(n_1699),
    .B(n_2477),
    .Y(n_2943));
 NOR2xp33_ASAP7_75t_SL g217810 (.A(n_1425),
    .B(n_2326),
    .Y(n_2941));
 AND2x2_ASAP7_75t_SL g217811 (.A(n_2436),
    .B(n_1664),
    .Y(n_2940));
 NOR2xp67_ASAP7_75t_SL g217812 (.A(sa31[4]),
    .B(n_2292),
    .Y(n_1722));
 NAND2xp5_ASAP7_75t_SL g217813 (.A(n_1653),
    .B(n_2468),
    .Y(n_1721));
 AND2x2_ASAP7_75t_R g217814 (.A(n_2475),
    .B(n_2425),
    .Y(n_2938));
 AND2x2_ASAP7_75t_L g217815 (.A(n_2474),
    .B(n_1659),
    .Y(n_2937));
 NOR2x1_ASAP7_75t_L g217816 (.A(n_1703),
    .B(n_2441),
    .Y(n_2936));
 AND2x2_ASAP7_75t_SL g217817 (.A(n_1944),
    .B(n_2314),
    .Y(n_2935));
 AND2x2_ASAP7_75t_SL g217818 (.A(n_1949),
    .B(n_1620),
    .Y(n_2934));
 NOR2xp33_ASAP7_75t_SL g217819 (.A(n_2507),
    .B(n_2056),
    .Y(n_2933));
 NAND2xp5_ASAP7_75t_L g217820 (.A(n_2572),
    .B(n_2416),
    .Y(n_2931));
 NAND2xp5_ASAP7_75t_R g217821 (.A(n_2439),
    .B(n_2618),
    .Y(n_2930));
 NAND2xp5_ASAP7_75t_SL g217822 (.A(n_8189),
    .B(n_2279),
    .Y(n_2929));
 OR2x2_ASAP7_75t_L g217823 (.A(n_2620),
    .B(n_2449),
    .Y(n_2927));
 NAND2xp5_ASAP7_75t_L g217824 (.A(n_2483),
    .B(n_1693),
    .Y(n_2924));
 NAND2xp5_ASAP7_75t_L g217825 (.A(n_1705),
    .B(n_2475),
    .Y(n_2922));
 OR2x2_ASAP7_75t_L g217826 (.A(n_2606),
    .B(n_2443),
    .Y(n_2921));
 AND2x2_ASAP7_75t_L g217827 (.A(n_8200),
    .B(n_1613),
    .Y(n_2919));
 AND2x2_ASAP7_75t_L g217828 (.A(n_2633),
    .B(n_2473),
    .Y(n_2918));
 NOR2xp33_ASAP7_75t_L g217829 (.A(n_2045),
    .B(n_2520),
    .Y(n_2917));
 NAND2x1_ASAP7_75t_SL g217830 (.A(n_1940),
    .B(n_2135),
    .Y(n_2916));
 NAND2x1_ASAP7_75t_SL g217831 (.A(n_1957),
    .B(n_2136),
    .Y(n_2914));
 NAND2xp5_ASAP7_75t_SL g217832 (.A(n_1384),
    .B(n_2328),
    .Y(n_2912));
 NAND2xp5_ASAP7_75t_R g217833 (.A(n_1386),
    .B(n_2328),
    .Y(n_2910));
 AND2x2_ASAP7_75t_SL g217834 (.A(n_1952),
    .B(n_2108),
    .Y(n_2908));
 NAND2xp5_ASAP7_75t_R g217835 (.A(n_2097),
    .B(n_8200),
    .Y(n_2905));
 NAND2xp5_ASAP7_75t_SL g217836 (.A(sa31[4]),
    .B(n_2291),
    .Y(n_2903));
 OR2x2_ASAP7_75t_SL g217837 (.A(n_1387),
    .B(n_2108),
    .Y(n_2902));
 NAND2x1_ASAP7_75t_SL g217838 (.A(n_1502),
    .B(n_2638),
    .Y(n_2900));
 NAND2xp5_ASAP7_75t_SL g217839 (.A(n_2200),
    .B(n_8189),
    .Y(n_2899));
 NOR2x1_ASAP7_75t_SL g217840 (.A(n_1425),
    .B(n_2185),
    .Y(n_2897));
 NOR2x1_ASAP7_75t_SL g217841 (.A(sa12[4]),
    .B(n_2133),
    .Y(n_2894));
 OR2x2_ASAP7_75t_SL g217842 (.A(n_1385),
    .B(n_2154),
    .Y(n_2893));
 NAND2xp5_ASAP7_75t_L g217843 (.A(n_1425),
    .B(n_2325),
    .Y(n_2890));
 AND2x2_ASAP7_75t_SL g217844 (.A(n_1852),
    .B(n_2144),
    .Y(n_2889));
 OR2x2_ASAP7_75t_SL g217845 (.A(n_2465),
    .B(n_2497),
    .Y(n_2887));
 AND2x2_ASAP7_75t_L g217846 (.A(n_1947),
    .B(n_2314),
    .Y(n_2885));
 AND2x2_ASAP7_75t_SL g217847 (.A(n_1375),
    .B(n_1620),
    .Y(n_2884));
 NAND2xp5_ASAP7_75t_R g217848 (.A(n_1387),
    .B(n_2287),
    .Y(n_2882));
 NOR2x1_ASAP7_75t_SL g217849 (.A(sa30[4]),
    .B(n_2150),
    .Y(n_1720));
 AND2x2_ASAP7_75t_L g217850 (.A(n_1853),
    .B(n_1613),
    .Y(n_2879));
 NAND2xp5_ASAP7_75t_L g217851 (.A(n_1851),
    .B(n_2279),
    .Y(n_2878));
 NAND2xp5_ASAP7_75t_R g217852 (.A(n_2286),
    .B(sa20[4]),
    .Y(n_1718));
 NAND2xp5_ASAP7_75t_SL g217853 (.A(n_1504),
    .B(n_1615),
    .Y(n_2875));
 NAND2x1_ASAP7_75t_SL g217854 (.A(n_1949),
    .B(n_2623),
    .Y(n_2873));
 AND2x2_ASAP7_75t_SL g217855 (.A(n_1950),
    .B(n_2500),
    .Y(n_2871));
 NAND2xp5_ASAP7_75t_SL g217856 (.A(n_1384),
    .B(n_2154),
    .Y(n_2869));
 NAND2x1_ASAP7_75t_L g217857 (.A(n_1948),
    .B(n_2185),
    .Y(n_2867));
 NOR2xp33_ASAP7_75t_SL g217858 (.A(n_1851),
    .B(n_1695),
    .Y(n_2864));
 OR2x2_ASAP7_75t_SL g217859 (.A(sa20[4]),
    .B(n_2106),
    .Y(n_2863));
 NOR2xp67_ASAP7_75t_SL g217860 (.A(n_1853),
    .B(n_1592),
    .Y(n_2861));
 AND2x2_ASAP7_75t_SL g217861 (.A(n_1949),
    .B(n_2455),
    .Y(n_2860));
 AND2x2_ASAP7_75t_SL g217862 (.A(n_1852),
    .B(n_1682),
    .Y(n_2858));
 AND2x4_ASAP7_75t_SL g217863 (.A(sa31[4]),
    .B(n_2480),
    .Y(n_2856));
 NAND2x1p5_ASAP7_75t_L g217864 (.A(n_8894),
    .B(n_2494),
    .Y(n_1715));
 NAND2x1p5_ASAP7_75t_SL g217865 (.A(n_1375),
    .B(n_1699),
    .Y(n_2854));
 AND2x2_ASAP7_75t_SL g217866 (.A(n_1384),
    .B(n_2606),
    .Y(n_2852));
 AND2x2_ASAP7_75t_L g217867 (.A(n_8189),
    .B(n_2466),
    .Y(n_2850));
 NOR2x1_ASAP7_75t_L g217868 (.A(sa03[4]),
    .B(n_2445),
    .Y(n_2848));
 AND2x4_ASAP7_75t_SL g217869 (.A(n_8896),
    .B(n_2619),
    .Y(n_2846));
 NOR2x1_ASAP7_75t_L g217870 (.A(n_1387),
    .B(n_2472),
    .Y(n_2844));
 AND2x4_ASAP7_75t_SL g217871 (.A(n_1387),
    .B(n_2633),
    .Y(n_2842));
 NAND2x1_ASAP7_75t_L g217872 (.A(n_1695),
    .B(n_1851),
    .Y(n_2840));
 AND2x2_ASAP7_75t_SL g217873 (.A(n_8200),
    .B(n_2490),
    .Y(n_2838));
 AND2x2_ASAP7_75t_SL g217874 (.A(n_1945),
    .B(n_2637),
    .Y(n_2834));
 NAND2x1_ASAP7_75t_SL g217875 (.A(n_1945),
    .B(n_2460),
    .Y(n_2833));
 OR2x2_ASAP7_75t_SL g217876 (.A(n_1385),
    .B(n_2447),
    .Y(n_2831));
 AND2x2_ASAP7_75t_SL g217877 (.A(n_1959),
    .B(n_2459),
    .Y(n_2829));
 OR2x2_ASAP7_75t_SL g217878 (.A(n_1941),
    .B(n_2460),
    .Y(n_2827));
 AND2x4_ASAP7_75t_SL g217879 (.A(n_1386),
    .B(n_2607),
    .Y(n_2825));
 NAND2x1_ASAP7_75t_SL g217880 (.A(n_1386),
    .B(n_2447),
    .Y(n_2823));
 AND2x2_ASAP7_75t_SL g217881 (.A(sa30[4]),
    .B(n_1672),
    .Y(n_2821));
 OR2x2_ASAP7_75t_SL g217882 (.A(n_8189),
    .B(n_2466),
    .Y(n_2819));
 AND2x4_ASAP7_75t_SL g217883 (.A(n_2461),
    .B(n_2637),
    .Y(n_2817));
 OR2x2_ASAP7_75t_SL g217884 (.A(n_2634),
    .B(n_2472),
    .Y(n_2815));
 NAND2x1p5_ASAP7_75t_SL g217885 (.A(n_1385),
    .B(n_2153),
    .Y(n_1713));
 AND2x2_ASAP7_75t_SL g217886 (.A(n_1345),
    .B(n_2607),
    .Y(n_2811));
 OR2x2_ASAP7_75t_SL g217887 (.A(n_1852),
    .B(n_2145),
    .Y(n_2807));
 OR2x2_ASAP7_75t_SL g217888 (.A(n_1952),
    .B(n_2108),
    .Y(n_2805));
 OR2x6_ASAP7_75t_SL g217889 (.A(n_2617),
    .B(n_2465),
    .Y(n_2803));
 NAND2xp5_ASAP7_75t_SL g217890 (.A(sa03[4]),
    .B(n_2186),
    .Y(n_2798));
 AND2x4_ASAP7_75t_SL g217891 (.A(n_1427),
    .B(n_2445),
    .Y(n_2797));
 NAND2xp5_ASAP7_75t_SL g217892 (.A(n_2263),
    .B(n_2097),
    .Y(n_2794));
 AND2x2_ASAP7_75t_SL g217893 (.A(n_2466),
    .B(n_1695),
    .Y(n_2793));
 AND2x2_ASAP7_75t_SL g217894 (.A(n_2455),
    .B(n_2622),
    .Y(n_2791));
 NAND2xp5_ASAP7_75t_SL g217895 (.A(n_1851),
    .B(n_2200),
    .Y(n_2788));
 AND2x4_ASAP7_75t_SL g217896 (.A(n_1947),
    .B(n_2135),
    .Y(n_2786));
 OR2x6_ASAP7_75t_SL g217897 (.A(n_2495),
    .B(n_2620),
    .Y(n_2784));
 AND2x2_ASAP7_75t_SL g217898 (.A(n_2491),
    .B(n_2635),
    .Y(n_2782));
 AND2x4_ASAP7_75t_SL g217899 (.A(n_1853),
    .B(n_1592),
    .Y(n_2780));
 AND2x2_ASAP7_75t_SL g217900 (.A(n_1375),
    .B(n_1598),
    .Y(n_2778));
 INVxp33_ASAP7_75t_R g217901 (.A(n_2730),
    .Y(n_2731));
 INVxp33_ASAP7_75t_R g217902 (.A(n_2727),
    .Y(n_2728));
 INVxp33_ASAP7_75t_R g217903 (.A(n_2725),
    .Y(n_2726));
 INVxp33_ASAP7_75t_R g217904 (.A(n_2714),
    .Y(n_2715));
 INVxp33_ASAP7_75t_R g217905 (.A(n_2710),
    .Y(n_2711));
 INVxp33_ASAP7_75t_R g217906 (.A(n_2708),
    .Y(n_2709));
 INVxp33_ASAP7_75t_R g217907 (.A(n_2705),
    .Y(n_2706));
 INVxp33_ASAP7_75t_R g217908 (.A(n_2703),
    .Y(n_2702));
 INVxp33_ASAP7_75t_R g217909 (.A(n_2699),
    .Y(n_2700));
 INVxp33_ASAP7_75t_R g217910 (.A(n_2697),
    .Y(n_2698));
 INVxp67_ASAP7_75t_R g217911 (.A(n_2692),
    .Y(n_2691));
 INVxp33_ASAP7_75t_R g217912 (.A(n_2689),
    .Y(n_2688));
 INVxp33_ASAP7_75t_R g217913 (.A(n_2686),
    .Y(n_2685));
 INVxp67_ASAP7_75t_R g217914 (.A(n_2683),
    .Y(n_2684));
 INVxp33_ASAP7_75t_R g217915 (.A(n_2682),
    .Y(n_2681));
 INVxp33_ASAP7_75t_R g217916 (.A(n_2679),
    .Y(n_2680));
 INVxp33_ASAP7_75t_R g217917 (.A(n_2678),
    .Y(n_2677));
 INVxp67_ASAP7_75t_L g217918 (.A(n_2675),
    .Y(n_2674));
 INVxp33_ASAP7_75t_R g217919 (.A(n_2672),
    .Y(n_2671));
 INVxp67_ASAP7_75t_R g217921 (.A(n_2668),
    .Y(n_2667));
 INVxp33_ASAP7_75t_R g217922 (.A(n_2666),
    .Y(n_2665));
 INVx1_ASAP7_75t_R g217923 (.A(n_2664),
    .Y(n_2663));
 INVxp67_ASAP7_75t_R g217924 (.A(n_2662),
    .Y(n_2661));
 INVxp67_ASAP7_75t_R g217926 (.A(n_1709),
    .Y(n_2660));
 HB1xp67_ASAP7_75t_SL g217927 (.A(n_2658),
    .Y(n_1709));
 INVxp67_ASAP7_75t_R g217928 (.A(n_2658),
    .Y(n_2659));
 INVx1_ASAP7_75t_L g217929 (.A(n_2657),
    .Y(n_2656));
 INVx1_ASAP7_75t_L g217932 (.A(n_1708),
    .Y(n_1707));
 INVx2_ASAP7_75t_SL g217935 (.A(n_2655),
    .Y(n_1708));
 INVxp33_ASAP7_75t_R g217936 (.A(ld_r),
    .Y(n_2654));
 INVxp67_ASAP7_75t_L g217937 (.A(n_2653),
    .Y(n_2652));
 INVxp67_ASAP7_75t_L g217938 (.A(n_2651),
    .Y(n_2650));
 INVxp67_ASAP7_75t_R g217939 (.A(n_2648),
    .Y(n_2647));
 INVxp33_ASAP7_75t_L g217940 (.A(n_2645),
    .Y(n_2644));
 INVx1_ASAP7_75t_L g217941 (.A(n_2643),
    .Y(n_2642));
 INVx1_ASAP7_75t_SL g217944 (.A(n_2640),
    .Y(n_1706));
 INVx1_ASAP7_75t_SL g217945 (.A(n_2639),
    .Y(n_2640));
 INVx1_ASAP7_75t_SL g217947 (.A(n_1338),
    .Y(n_2639));
 INVx1_ASAP7_75t_L g217948 (.A(n_2637),
    .Y(n_2638));
 INVxp33_ASAP7_75t_R g217950 (.A(n_1705),
    .Y(n_2636));
 BUFx2_ASAP7_75t_SL g217951 (.A(n_2637),
    .Y(n_1705));
 INVxp67_ASAP7_75t_SL g217957 (.A(n_1704),
    .Y(n_1703));
 BUFx2_ASAP7_75t_SL g217958 (.A(n_2635),
    .Y(n_1704));
 INVxp67_ASAP7_75t_R g217960 (.A(n_1701),
    .Y(n_1702));
 INVx2_ASAP7_75t_SL g217962 (.A(n_2634),
    .Y(n_2633));
 INVxp67_ASAP7_75t_L g217963 (.A(n_2632),
    .Y(n_2631));
 INVx1_ASAP7_75t_R g217966 (.A(n_1700),
    .Y(n_2630));
 INVxp67_ASAP7_75t_R g217968 (.A(n_2629),
    .Y(n_2628));
 INVx1_ASAP7_75t_R g217969 (.A(n_2627),
    .Y(n_2626));
 INVxp67_ASAP7_75t_R g217970 (.A(n_2625),
    .Y(n_2624));
 INVxp67_ASAP7_75t_SL g217971 (.A(n_2622),
    .Y(n_2623));
 INVxp67_ASAP7_75t_R g217972 (.A(n_1699),
    .Y(n_2621));
 BUFx3_ASAP7_75t_SL g217974 (.A(n_2622),
    .Y(n_1699));
 INVx2_ASAP7_75t_SL g217975 (.A(n_2620),
    .Y(n_2619));
 INVx2_ASAP7_75t_SL g217976 (.A(n_2618),
    .Y(n_2617));
 INVxp33_ASAP7_75t_R g217981 (.A(n_1698),
    .Y(n_1697));
 HB1xp67_ASAP7_75t_L g217982 (.A(n_2616),
    .Y(n_1698));
 INVxp67_ASAP7_75t_L g217983 (.A(n_2615),
    .Y(n_2614));
 INVx1_ASAP7_75t_R g217984 (.A(n_2613),
    .Y(n_2612));
 INVxp67_ASAP7_75t_R g217985 (.A(n_2611),
    .Y(n_2610));
 INVx1_ASAP7_75t_R g217986 (.A(n_2609),
    .Y(n_2608));
 INVx2_ASAP7_75t_SL g217987 (.A(n_2607),
    .Y(n_2606));
 INVxp67_ASAP7_75t_R g217988 (.A(n_2605),
    .Y(n_2604));
 INVxp67_ASAP7_75t_R g217989 (.A(n_2603),
    .Y(n_2602));
 INVxp67_ASAP7_75t_R g217990 (.A(n_2601),
    .Y(n_2600));
 INVxp33_ASAP7_75t_R g217991 (.A(n_1696),
    .Y(n_2599));
 INVx1_ASAP7_75t_L g218000 (.A(n_1694),
    .Y(n_1693));
 INVx1_ASAP7_75t_L g218002 (.A(n_1695),
    .Y(n_1694));
 INVxp33_ASAP7_75t_R g218004 (.A(n_2598),
    .Y(n_2597));
 INVx1_ASAP7_75t_SL g218005 (.A(n_2596),
    .Y(n_2595));
 INVxp67_ASAP7_75t_R g218006 (.A(n_2594),
    .Y(n_2593));
 INVx1_ASAP7_75t_L g218007 (.A(n_2592),
    .Y(n_2591));
 INVx1_ASAP7_75t_R g218008 (.A(n_2590),
    .Y(n_2589));
 INVx1_ASAP7_75t_L g218009 (.A(n_2588),
    .Y(n_2587));
 INVx1_ASAP7_75t_L g218010 (.A(n_2586),
    .Y(n_2585));
 INVx1_ASAP7_75t_R g218011 (.A(n_2584),
    .Y(n_2583));
 INVxp33_ASAP7_75t_R g218012 (.A(n_2582),
    .Y(n_2581));
 INVxp67_ASAP7_75t_L g218013 (.A(n_2580),
    .Y(n_2579));
 INVx2_ASAP7_75t_L g218014 (.A(n_2578),
    .Y(n_2577));
 INVx1_ASAP7_75t_SL g218015 (.A(n_2576),
    .Y(n_2575));
 INVxp33_ASAP7_75t_R g218016 (.A(n_2574),
    .Y(n_2573));
 INVx1_ASAP7_75t_SL g218017 (.A(n_2572),
    .Y(n_2571));
 INVxp67_ASAP7_75t_R g218018 (.A(n_2570),
    .Y(n_2569));
 INVx2_ASAP7_75t_SL g218019 (.A(n_2568),
    .Y(n_2567));
 INVx1_ASAP7_75t_SL g218020 (.A(n_2566),
    .Y(n_2565));
 INVx1_ASAP7_75t_L g218021 (.A(n_2564),
    .Y(n_2563));
 INVxp67_ASAP7_75t_L g218022 (.A(n_2562),
    .Y(n_2561));
 INVx1_ASAP7_75t_R g218023 (.A(n_2560),
    .Y(n_2559));
 INVx1_ASAP7_75t_L g218024 (.A(n_2558),
    .Y(n_2557));
 INVx1_ASAP7_75t_SL g218025 (.A(n_2556),
    .Y(n_2555));
 INVx2_ASAP7_75t_SL g218026 (.A(n_2554),
    .Y(n_2553));
 INVx1_ASAP7_75t_L g218027 (.A(n_2552),
    .Y(n_2551));
 INVx1_ASAP7_75t_L g218028 (.A(n_2550),
    .Y(n_2549));
 INVxp67_ASAP7_75t_R g218029 (.A(n_2548),
    .Y(n_2547));
 INVx1_ASAP7_75t_R g218030 (.A(n_2546),
    .Y(n_2545));
 INVx1_ASAP7_75t_R g218031 (.A(n_2544),
    .Y(n_2543));
 INVxp67_ASAP7_75t_R g218032 (.A(n_2542),
    .Y(n_2541));
 INVx2_ASAP7_75t_L g218033 (.A(n_2540),
    .Y(n_2539));
 INVx2_ASAP7_75t_SL g218034 (.A(n_2538),
    .Y(n_2537));
 INVx3_ASAP7_75t_SL g218035 (.A(n_2536),
    .Y(n_2535));
 INVx1_ASAP7_75t_SL g218036 (.A(n_2534),
    .Y(n_2533));
 INVx1_ASAP7_75t_SL g218037 (.A(n_2532),
    .Y(n_2531));
 INVx2_ASAP7_75t_SL g218038 (.A(n_2530),
    .Y(n_2529));
 INVx1_ASAP7_75t_R g218039 (.A(n_2528),
    .Y(n_2527));
 INVx1_ASAP7_75t_L g218040 (.A(n_2526),
    .Y(n_2525));
 INVx1_ASAP7_75t_SL g218041 (.A(n_2524),
    .Y(n_2523));
 INVx1_ASAP7_75t_SL g218042 (.A(n_2522),
    .Y(n_2521));
 INVx1_ASAP7_75t_L g218043 (.A(n_2520),
    .Y(n_2519));
 INVx2_ASAP7_75t_SL g218044 (.A(n_2518),
    .Y(n_2517));
 INVx1_ASAP7_75t_SL g218046 (.A(n_1691),
    .Y(n_1690));
 INVx1_ASAP7_75t_SL g218052 (.A(n_2515),
    .Y(n_2514));
 INVx2_ASAP7_75t_L g218053 (.A(n_2513),
    .Y(n_2512));
 INVx2_ASAP7_75t_L g218058 (.A(n_2511),
    .Y(n_1689));
 INVx2_ASAP7_75t_SL g218061 (.A(n_2510),
    .Y(n_2509));
 INVx2_ASAP7_75t_SL g218062 (.A(n_2508),
    .Y(n_2507));
 INVx1_ASAP7_75t_SL g218063 (.A(n_2506),
    .Y(n_2505));
 INVx2_ASAP7_75t_SL g218064 (.A(n_2504),
    .Y(n_2503));
 INVx4_ASAP7_75t_SL g218065 (.A(n_2502),
    .Y(n_2501));
 INVx2_ASAP7_75t_L g218066 (.A(n_2500),
    .Y(n_2499));
 INVx1_ASAP7_75t_L g218071 (.A(n_1688),
    .Y(n_1687));
 INVx1_ASAP7_75t_SL g218074 (.A(n_1686),
    .Y(n_1688));
 INVx2_ASAP7_75t_SL g218076 (.A(n_2497),
    .Y(n_2496));
 INVx2_ASAP7_75t_SL g218077 (.A(n_2495),
    .Y(n_2494));
 INVxp67_ASAP7_75t_L g218084 (.A(n_1683),
    .Y(n_2492));
 BUFx3_ASAP7_75t_SL g218085 (.A(n_2491),
    .Y(n_1683));
 INVx2_ASAP7_75t_SL g218090 (.A(n_2490),
    .Y(n_2489));
 INVx1_ASAP7_75t_SL g218091 (.A(n_2488),
    .Y(n_2487));
 INVx1_ASAP7_75t_SL g218092 (.A(n_2486),
    .Y(n_2485));
 INVx2_ASAP7_75t_SL g218093 (.A(n_2484),
    .Y(n_2483));
 INVx2_ASAP7_75t_L g218094 (.A(n_2482),
    .Y(n_2481));
 INVxp67_ASAP7_75t_L g218097 (.A(n_1682),
    .Y(n_1681));
 BUFx2_ASAP7_75t_SL g218102 (.A(n_2479),
    .Y(n_1682));
 INVx1_ASAP7_75t_L g218103 (.A(n_2479),
    .Y(n_2480));
 INVx3_ASAP7_75t_SL g218104 (.A(n_2478),
    .Y(n_2477));
 INVx2_ASAP7_75t_SL g218105 (.A(n_2476),
    .Y(n_2475));
 INVx2_ASAP7_75t_L g218106 (.A(n_2474),
    .Y(n_2473));
 INVx2_ASAP7_75t_L g218107 (.A(n_2472),
    .Y(n_2471));
 INVx2_ASAP7_75t_L g218108 (.A(n_2470),
    .Y(n_2469));
 INVx2_ASAP7_75t_SL g218109 (.A(n_2468),
    .Y(n_2467));
 INVx1_ASAP7_75t_L g218114 (.A(n_1679),
    .Y(n_1680));
 INVx1_ASAP7_75t_L g218117 (.A(n_2466),
    .Y(n_1679));
 INVx1_ASAP7_75t_L g218120 (.A(n_2465),
    .Y(n_2464));
 INVx3_ASAP7_75t_SL g218121 (.A(n_2463),
    .Y(n_2462));
 INVx1_ASAP7_75t_SL g218122 (.A(n_2460),
    .Y(n_2461));
 INVx2_ASAP7_75t_L g218129 (.A(n_1677),
    .Y(n_1678));
 INVx2_ASAP7_75t_SL g218130 (.A(n_2460),
    .Y(n_1677));
 INVx2_ASAP7_75t_L g218134 (.A(n_1675),
    .Y(n_1676));
 BUFx3_ASAP7_75t_SL g218136 (.A(n_2459),
    .Y(n_1675));
 INVxp33_ASAP7_75t_R g218142 (.A(n_1674),
    .Y(n_2458));
 INVx3_ASAP7_75t_SL g218144 (.A(n_2459),
    .Y(n_1674));
 INVx4_ASAP7_75t_SL g218145 (.A(n_2457),
    .Y(n_2456));
 INVx2_ASAP7_75t_L g218156 (.A(n_1673),
    .Y(n_1671));
 INVx2_ASAP7_75t_L g218157 (.A(n_1672),
    .Y(n_1673));
 INVx2_ASAP7_75t_SL g218158 (.A(n_2455),
    .Y(n_1672));
 INVx2_ASAP7_75t_SL g218159 (.A(n_2453),
    .Y(n_2452));
 INVx3_ASAP7_75t_SL g218160 (.A(n_2451),
    .Y(n_2450));
 INVx3_ASAP7_75t_SL g218161 (.A(n_2449),
    .Y(n_2448));
 INVxp67_ASAP7_75t_L g218165 (.A(n_2446),
    .Y(n_1670));
 INVxp67_ASAP7_75t_SL g218167 (.A(n_1345),
    .Y(n_2446));
 INVx4_ASAP7_75t_SL g218168 (.A(n_2445),
    .Y(n_2444));
 INVx2_ASAP7_75t_R g218169 (.A(n_2443),
    .Y(n_2442));
 INVx2_ASAP7_75t_SL g218170 (.A(n_2441),
    .Y(n_2440));
 INVx2_ASAP7_75t_SL g218171 (.A(n_2439),
    .Y(n_2438));
 INVx2_ASAP7_75t_R g218172 (.A(n_2437),
    .Y(n_2436));
 INVx2_ASAP7_75t_SL g218173 (.A(n_2435),
    .Y(n_2434));
 INVxp33_ASAP7_75t_R g218174 (.A(n_2432),
    .Y(n_2433));
 INVxp67_ASAP7_75t_R g218183 (.A(n_1669),
    .Y(n_1668));
 INVx2_ASAP7_75t_SL g218184 (.A(n_2431),
    .Y(n_1669));
 INVx1_ASAP7_75t_L g218190 (.A(n_1667),
    .Y(n_1666));
 BUFx2_ASAP7_75t_SL g218193 (.A(n_2431),
    .Y(n_1667));
 BUFx3_ASAP7_75t_SL g218195 (.A(n_1665),
    .Y(n_2430));
 BUFx2_ASAP7_75t_L g218209 (.A(n_1664),
    .Y(n_1663));
 INVx1_ASAP7_75t_SL g218215 (.A(n_2429),
    .Y(n_1660));
 BUFx2_ASAP7_75t_SL g218219 (.A(n_1659),
    .Y(n_2429));
 INVx2_ASAP7_75t_SL g218229 (.A(n_1659),
    .Y(n_1662));
 INVx2_ASAP7_75t_SL g218230 (.A(n_2428),
    .Y(n_2427));
 INVx1_ASAP7_75t_SL g218233 (.A(n_1657),
    .Y(n_1658));
 INVx3_ASAP7_75t_SL g218240 (.A(n_1656),
    .Y(n_1657));
 INVx2_ASAP7_75t_R g218255 (.A(n_1656),
    .Y(n_1655));
 INVx2_ASAP7_75t_SL g218257 (.A(n_2425),
    .Y(n_2424));
 BUFx2_ASAP7_75t_L g218259 (.A(n_2423),
    .Y(n_2422));
 BUFx2_ASAP7_75t_R g218262 (.A(n_2420),
    .Y(n_2421));
 HB1xp67_ASAP7_75t_SL g218265 (.A(n_2418),
    .Y(n_2419));
 BUFx2_ASAP7_75t_R g218267 (.A(n_2418),
    .Y(n_1654));
 INVx1_ASAP7_75t_L g218270 (.A(n_2417),
    .Y(n_1652));
 INVx1_ASAP7_75t_R g218272 (.A(n_1653),
    .Y(n_2417));
 INVx2_ASAP7_75t_SL g218275 (.A(n_2416),
    .Y(n_2415));
 BUFx2_ASAP7_75t_SL g218277 (.A(n_2413),
    .Y(n_2414));
 INVxp33_ASAP7_75t_R g218286 (.A(n_1650),
    .Y(n_2412));
 INVxp67_ASAP7_75t_R g218289 (.A(n_1651),
    .Y(n_1650));
 INVx2_ASAP7_75t_R g218290 (.A(n_2411),
    .Y(n_2410));
 INVxp67_ASAP7_75t_R g218315 (.A(n_2404),
    .Y(n_2403));
 BUFx2_ASAP7_75t_R g218316 (.A(n_2401),
    .Y(n_2404));
 INVx2_ASAP7_75t_R g218324 (.A(n_2401),
    .Y(n_1647));
 INVxp67_ASAP7_75t_R g218330 (.A(n_1646),
    .Y(n_2402));
 INVxp67_ASAP7_75t_SL g218332 (.A(n_2401),
    .Y(n_1646));
 INVx4_ASAP7_75t_SL g218338 (.A(n_2400),
    .Y(n_2399));
 INVx2_ASAP7_75t_SL g218348 (.A(n_1642),
    .Y(n_1643));
 INVx2_ASAP7_75t_SL g218354 (.A(n_1645),
    .Y(n_1642));
 INVx2_ASAP7_75t_L g218357 (.A(n_1644),
    .Y(n_2398));
 INVx3_ASAP7_75t_SL g218360 (.A(n_1645),
    .Y(n_1644));
 INVx3_ASAP7_75t_SL g218370 (.A(n_2397),
    .Y(n_2396));
 INVx4_ASAP7_75t_SL g218371 (.A(n_2395),
    .Y(n_2394));
 INVx4_ASAP7_75t_SL g218372 (.A(n_2393),
    .Y(n_2392));
 INVx1_ASAP7_75t_SL g218376 (.A(n_1641),
    .Y(n_1640));
 INVx2_ASAP7_75t_L g218393 (.A(n_1445),
    .Y(n_1639));
 BUFx2_ASAP7_75t_L g218395 (.A(n_2389),
    .Y(n_1638));
 HB1xp67_ASAP7_75t_L g218399 (.A(n_2389),
    .Y(n_2390));
 HB1xp67_ASAP7_75t_L g218408 (.A(n_1637),
    .Y(n_2388));
 INVxp67_ASAP7_75t_SL g218411 (.A(n_1636),
    .Y(n_1635));
 INVx1_ASAP7_75t_L g218424 (.A(n_1632),
    .Y(n_2386));
 INVx2_ASAP7_75t_SL g218426 (.A(n_2387),
    .Y(n_1632));
 INVx2_ASAP7_75t_L g218428 (.A(n_1633),
    .Y(n_1634));
 INVx1_ASAP7_75t_R g218444 (.A(n_1350),
    .Y(n_1629));
 INVx2_ASAP7_75t_L g218456 (.A(n_1628),
    .Y(n_1627));
 INVx4_ASAP7_75t_SL g218457 (.A(n_1350),
    .Y(n_1628));
 INVxp67_ASAP7_75t_SL g218459 (.A(n_2385),
    .Y(n_1626));
 INVx1_ASAP7_75t_SL g218469 (.A(n_1622),
    .Y(n_1623));
 INVx1_ASAP7_75t_SL g218475 (.A(n_1625),
    .Y(n_1624));
 NAND2xp33_ASAP7_75t_R g218478 (.A(n_1950),
    .B(n_1867),
    .Y(n_2384));
 NAND2xp33_ASAP7_75t_R g218479 (.A(n_1507),
    .B(n_8894),
    .Y(n_2730));
 NAND2xp33_ASAP7_75t_R g218480 (.A(n_1967),
    .B(n_1948),
    .Y(n_2729));
 NOR2xp33_ASAP7_75t_R g218481 (.A(sa10[4]),
    .B(n_1972),
    .Y(n_2727));
 NOR2xp33_ASAP7_75t_R g218482 (.A(sa22[4]),
    .B(sa22[3]),
    .Y(n_2725));
 NOR2xp33_ASAP7_75t_R g218483 (.A(sa23[4]),
    .B(sa23[3]),
    .Y(n_2724));
 NAND2xp33_ASAP7_75t_R g218484 (.A(n_8182),
    .B(n_8209),
    .Y(n_2723));
 NOR2xp33_ASAP7_75t_R g218485 (.A(sa32[5]),
    .B(n_1980),
    .Y(n_2722));
 NOR2xp33_ASAP7_75t_R g218486 (.A(sa00[0]),
    .B(sa00[5]),
    .Y(n_2721));
 NOR2xp33_ASAP7_75t_R g218487 (.A(sa32[2]),
    .B(sa32[5]),
    .Y(n_2720));
 NOR2xp33_ASAP7_75t_R g218488 (.A(sa33[2]),
    .B(sa33[5]),
    .Y(n_2719));
 NOR2xp33_ASAP7_75t_R g218489 (.A(sa21[2]),
    .B(n_8183),
    .Y(n_2718));
 NAND2xp33_ASAP7_75t_R g218490 (.A(n_8183),
    .B(n_1968),
    .Y(n_2717));
 NOR2xp33_ASAP7_75t_R g218491 (.A(n_1865),
    .B(sa11[2]),
    .Y(n_2716));
 NOR2xp33_ASAP7_75t_R g218492 (.A(sa01[3]),
    .B(n_1385),
    .Y(n_2714));
 NAND2xp33_ASAP7_75t_R g218493 (.A(n_2009),
    .B(n_1538),
    .Y(n_2713));
 NOR2xp33_ASAP7_75t_R g218494 (.A(n_1532),
    .B(n_2022),
    .Y(n_2712));
 NAND2xp33_ASAP7_75t_R g218495 (.A(n_1888),
    .B(n_1917),
    .Y(n_2710));
 NAND2xp33_ASAP7_75t_R g218496 (.A(n_8208),
    .B(n_1913),
    .Y(n_2708));
 NOR2xp33_ASAP7_75t_R g218497 (.A(sa01[2]),
    .B(sa01[5]),
    .Y(n_2707));
 NOR2xp33_ASAP7_75t_R g218498 (.A(sa33[5]),
    .B(sa33[0]),
    .Y(n_2705));
 NOR2xp33_ASAP7_75t_R g218499 (.A(sa23[0]),
    .B(sa23[5]),
    .Y(n_2704));
 NAND2xp33_ASAP7_75t_R g218500 (.A(n_1494),
    .B(n_8207),
    .Y(n_2703));
 NAND2xp5_ASAP7_75t_R g218501 (.A(n_1884),
    .B(n_1877),
    .Y(n_2701));
 NAND2xp33_ASAP7_75t_R g218502 (.A(sa31[5]),
    .B(n_1926),
    .Y(n_2699));
 NOR2xp33_ASAP7_75t_R g218503 (.A(n_1528),
    .B(sa10[5]),
    .Y(n_2697));
 NOR2xp33_ASAP7_75t_R g218504 (.A(sa30[0]),
    .B(sa30[5]),
    .Y(n_2696));
 NAND2xp5_ASAP7_75t_R g218505 (.A(n_8217),
    .B(n_1879),
    .Y(n_2695));
 NOR2xp33_ASAP7_75t_L g218506 (.A(n_1923),
    .B(sa20[5]),
    .Y(n_2694));
 NOR2xp33_ASAP7_75t_R g218507 (.A(sa22[2]),
    .B(sa22[5]),
    .Y(n_2693));
 NOR2xp33_ASAP7_75t_R g218508 (.A(sa00[2]),
    .B(sa00[5]),
    .Y(n_2692));
 NOR2xp33_ASAP7_75t_L g218509 (.A(sa30[2]),
    .B(sa30[5]),
    .Y(n_2690));
 NOR2xp33_ASAP7_75t_R g218510 (.A(sa31[2]),
    .B(sa31[5]),
    .Y(n_2689));
 NOR2xp33_ASAP7_75t_L g218511 (.A(sa12[2]),
    .B(n_1912),
    .Y(n_2687));
 NAND2xp5_ASAP7_75t_L g218512 (.A(n_8179),
    .B(n_1888),
    .Y(n_2686));
 NAND2xp33_ASAP7_75t_R g218513 (.A(n_1981),
    .B(n_8203),
    .Y(n_2683));
 NOR2xp33_ASAP7_75t_L g218514 (.A(sa21[2]),
    .B(sa21[5]),
    .Y(n_2682));
 NOR2xp33_ASAP7_75t_R g218515 (.A(sa12[2]),
    .B(sa12[0]),
    .Y(n_2679));
 NOR2xp33_ASAP7_75t_R g218516 (.A(sa00[2]),
    .B(sa00[0]),
    .Y(n_2678));
 AND2x2_ASAP7_75t_R g218517 (.A(n_1533),
    .B(n_1509),
    .Y(n_2676));
 OR2x2_ASAP7_75t_SL g218518 (.A(n_1896),
    .B(n_1478),
    .Y(n_2675));
 NOR2xp33_ASAP7_75t_R g218519 (.A(sa30[0]),
    .B(sa30[2]),
    .Y(n_2673));
 NAND2xp5_ASAP7_75t_R g218520 (.A(n_8217),
    .B(n_2026),
    .Y(n_2672));
 NOR2xp33_ASAP7_75t_R g218521 (.A(sa11[2]),
    .B(sa11[0]),
    .Y(n_2670));
 NOR2xp33_ASAP7_75t_R g218522 (.A(sa21[2]),
    .B(sa21[0]),
    .Y(n_2668));
 NOR2xp33_ASAP7_75t_L g218523 (.A(sa01[0]),
    .B(sa01[2]),
    .Y(n_2666));
 NOR2xp33_ASAP7_75t_R g218524 (.A(sa33[0]),
    .B(sa33[2]),
    .Y(n_2664));
 NOR2xp33_ASAP7_75t_L g218525 (.A(n_1495),
    .B(n_1966),
    .Y(n_2662));
 OR2x2_ASAP7_75t_SL g218526 (.A(sa20[1]),
    .B(sa20[7]),
    .Y(n_2658));
 NAND2xp5_ASAP7_75t_L g218527 (.A(sa20[0]),
    .B(n_1923),
    .Y(n_2657));
 NOR2x1_ASAP7_75t_SL g218528 (.A(sa12[1]),
    .B(sa12[7]),
    .Y(n_2655));
 NOR2xp33_ASAP7_75t_L g218530 (.A(n_2034),
    .B(n_1365),
    .Y(n_2653));
 OR2x2_ASAP7_75t_SL g218531 (.A(sa13[7]),
    .B(sa13[1]),
    .Y(n_2651));
 AND2x2_ASAP7_75t_L g218532 (.A(sa21[0]),
    .B(n_1925),
    .Y(n_2649));
 AND2x2_ASAP7_75t_L g218533 (.A(n_2012),
    .B(n_1538),
    .Y(n_2648));
 AND2x2_ASAP7_75t_R g218534 (.A(n_8213),
    .B(n_1926),
    .Y(n_2646));
 OR2x2_ASAP7_75t_SL g218535 (.A(sa10[7]),
    .B(sa10[1]),
    .Y(n_2645));
 NAND2x1p5_ASAP7_75t_SL g218536 (.A(n_1513),
    .B(n_1916),
    .Y(n_2643));
 OR2x2_ASAP7_75t_SL g218538 (.A(sa21[7]),
    .B(sa21[1]),
    .Y(n_2637));
 NAND2xp5_ASAP7_75t_SL g218539 (.A(n_2029),
    .B(n_1874),
    .Y(n_2635));
 OR2x2_ASAP7_75t_SL g218540 (.A(sa03[7]),
    .B(sa03[1]),
    .Y(n_1701));
 AND2x2_ASAP7_75t_SL g218541 (.A(n_8184),
    .B(n_2017),
    .Y(n_2634));
 AND2x2_ASAP7_75t_SL g218542 (.A(sa21[2]),
    .B(n_1968),
    .Y(n_2632));
 NAND2xp5_ASAP7_75t_L g218543 (.A(sa21[0]),
    .B(sa21[2]),
    .Y(n_1700));
 AND2x2_ASAP7_75t_R g218544 (.A(sa30[0]),
    .B(sa30[2]),
    .Y(n_2629));
 AND2x2_ASAP7_75t_L g218545 (.A(sa31[2]),
    .B(n_8213),
    .Y(n_2627));
 NAND2xp5_ASAP7_75t_R g218546 (.A(n_1926),
    .B(n_1866),
    .Y(n_2625));
 NAND2xp5_ASAP7_75t_SL g218547 (.A(n_8187),
    .B(n_8205),
    .Y(n_2622));
 AND2x2_ASAP7_75t_SL g218548 (.A(n_1990),
    .B(n_1908),
    .Y(n_2620));
 OR2x6_ASAP7_75t_SL g218549 (.A(sa02[1]),
    .B(sa02[7]),
    .Y(n_2618));
 NAND2xp5_ASAP7_75t_L g218550 (.A(sa00[0]),
    .B(sa00[2]),
    .Y(n_2616));
 AND2x2_ASAP7_75t_L g218551 (.A(n_1866),
    .B(sa31[2]),
    .Y(n_2615));
 OR2x2_ASAP7_75t_L g218552 (.A(n_1466),
    .B(sa20[4]),
    .Y(n_2613));
 AND2x2_ASAP7_75t_L g218553 (.A(sa12[0]),
    .B(sa12[2]),
    .Y(n_2611));
 NAND2x1_ASAP7_75t_SL g218554 (.A(sa32[2]),
    .B(n_1980),
    .Y(n_2609));
 OR2x2_ASAP7_75t_SL g218555 (.A(sa01[1]),
    .B(sa01[7]),
    .Y(n_2607));
 AND2x2_ASAP7_75t_L g218556 (.A(n_1856),
    .B(n_1513),
    .Y(n_2605));
 AND2x2_ASAP7_75t_R g218557 (.A(sa01[2]),
    .B(sa01[0]),
    .Y(n_2603));
 AND2x2_ASAP7_75t_SL g218558 (.A(n_1532),
    .B(n_1510),
    .Y(n_2601));
 NAND2xp5_ASAP7_75t_R g218559 (.A(sa22[0]),
    .B(sa22[2]),
    .Y(n_1696));
 NAND2x1p5_ASAP7_75t_L g218560 (.A(n_8204),
    .B(n_8191),
    .Y(n_1695));
 AND2x2_ASAP7_75t_R g218561 (.A(sa23[0]),
    .B(sa23[2]),
    .Y(n_2598));
 AND2x2_ASAP7_75t_L g218562 (.A(sa02[0]),
    .B(n_2034),
    .Y(n_2596));
 AND2x2_ASAP7_75t_L g218563 (.A(n_1960),
    .B(n_1871),
    .Y(n_2594));
 NAND2xp5_ASAP7_75t_SL g218564 (.A(n_1480),
    .B(n_1952),
    .Y(n_2592));
 AND2x2_ASAP7_75t_SL g218565 (.A(n_1891),
    .B(n_8200),
    .Y(n_2590));
 AND2x2_ASAP7_75t_SL g218566 (.A(n_2024),
    .B(n_1948),
    .Y(n_2588));
 AND2x2_ASAP7_75t_SL g218567 (.A(n_8200),
    .B(n_8206),
    .Y(n_2586));
 AND2x2_ASAP7_75t_SL g218568 (.A(n_1914),
    .B(n_1384),
    .Y(n_2584));
 NAND2xp5_ASAP7_75t_SL g218569 (.A(sa33[0]),
    .B(sa33[2]),
    .Y(n_2582));
 AND2x2_ASAP7_75t_L g218570 (.A(n_2020),
    .B(n_1948),
    .Y(n_2580));
 NAND2x1p5_ASAP7_75t_L g218571 (.A(n_1466),
    .B(sa20[4]),
    .Y(n_2578));
 AND2x2_ASAP7_75t_SL g218572 (.A(n_1953),
    .B(n_2019),
    .Y(n_2576));
 OR2x2_ASAP7_75t_SL g218573 (.A(n_1941),
    .B(n_1522),
    .Y(n_2574));
 AND2x2_ASAP7_75t_SL g218574 (.A(n_1905),
    .B(n_1851),
    .Y(n_2572));
 AND2x2_ASAP7_75t_R g218575 (.A(n_8204),
    .B(n_8189),
    .Y(n_2570));
 NAND2x1p5_ASAP7_75t_SL g218576 (.A(n_1852),
    .B(n_2006),
    .Y(n_2568));
 AND2x2_ASAP7_75t_SL g218577 (.A(n_1966),
    .B(n_1495),
    .Y(n_2566));
 OR2x2_ASAP7_75t_SL g218578 (.A(n_1492),
    .B(n_1385),
    .Y(n_2564));
 AND2x2_ASAP7_75t_SL g218579 (.A(n_2016),
    .B(n_1952),
    .Y(n_2562));
 AND2x2_ASAP7_75t_SL g218580 (.A(n_1486),
    .B(n_1852),
    .Y(n_2560));
 AND2x2_ASAP7_75t_L g218581 (.A(n_1982),
    .B(n_8212),
    .Y(n_2558));
 OR2x2_ASAP7_75t_SL g218582 (.A(sa30[4]),
    .B(n_1900),
    .Y(n_2556));
 AND2x2_ASAP7_75t_SL g218583 (.A(n_1959),
    .B(n_2001),
    .Y(n_2554));
 AND2x2_ASAP7_75t_L g218584 (.A(n_1475),
    .B(n_1949),
    .Y(n_2552));
 AND2x2_ASAP7_75t_L g218585 (.A(n_1880),
    .B(n_1957),
    .Y(n_2550));
 AND2x2_ASAP7_75t_L g218586 (.A(n_1471),
    .B(n_1855),
    .Y(n_2548));
 AND2x2_ASAP7_75t_SL g218587 (.A(n_1995),
    .B(n_8908),
    .Y(n_2546));
 AND2x2_ASAP7_75t_L g218588 (.A(n_1987),
    .B(n_1953),
    .Y(n_2544));
 AND2x2_ASAP7_75t_R g218589 (.A(sa11[0]),
    .B(sa11[2]),
    .Y(n_2542));
 OR2x2_ASAP7_75t_SL g218590 (.A(n_1851),
    .B(n_2014),
    .Y(n_2540));
 AND2x2_ASAP7_75t_SL g218591 (.A(n_1994),
    .B(sa32[4]),
    .Y(n_2538));
 OR2x2_ASAP7_75t_SL g218592 (.A(n_1940),
    .B(n_1523),
    .Y(n_2536));
 OR2x2_ASAP7_75t_SL g218593 (.A(n_1855),
    .B(n_1469),
    .Y(n_2534));
 AND2x2_ASAP7_75t_SL g218594 (.A(sa31[4]),
    .B(n_1487),
    .Y(n_2532));
 AND2x4_ASAP7_75t_SL g218595 (.A(n_1909),
    .B(n_8894),
    .Y(n_2530));
 AND2x2_ASAP7_75t_SL g218596 (.A(sa23[4]),
    .B(sa23[1]),
    .Y(n_2528));
 AND2x2_ASAP7_75t_SL g218597 (.A(sa10[4]),
    .B(sa10[1]),
    .Y(n_2526));
 AND2x2_ASAP7_75t_SL g218598 (.A(n_2011),
    .B(n_1939),
    .Y(n_2524));
 AND2x2_ASAP7_75t_SL g218599 (.A(n_8212),
    .B(n_2010),
    .Y(n_2522));
 AND2x2_ASAP7_75t_SL g218600 (.A(sa11[4]),
    .B(n_1479),
    .Y(n_2520));
 OR2x2_ASAP7_75t_SL g218601 (.A(sa20[4]),
    .B(sa20[7]),
    .Y(n_2518));
 NAND2x1p5_ASAP7_75t_SL g218602 (.A(sa01[1]),
    .B(sa01[4]),
    .Y(n_1691));
 AND2x4_ASAP7_75t_SL g218603 (.A(n_1856),
    .B(n_1916),
    .Y(n_2515));
 AND2x2_ASAP7_75t_L g218604 (.A(n_1886),
    .B(sa30[4]),
    .Y(n_2513));
 AND2x2_ASAP7_75t_SL g218605 (.A(sa03[4]),
    .B(sa03[1]),
    .Y(n_2511));
 AND2x2_ASAP7_75t_SL g218606 (.A(sa12[4]),
    .B(sa12[1]),
    .Y(n_2510));
 OR2x2_ASAP7_75t_SL g218607 (.A(n_8200),
    .B(n_8198),
    .Y(n_2508));
 AND2x4_ASAP7_75t_SL g218608 (.A(n_1921),
    .B(n_1960),
    .Y(n_2506));
 AND2x4_ASAP7_75t_SL g218609 (.A(n_1506),
    .B(n_1472),
    .Y(n_2504));
 OR2x2_ASAP7_75t_SL g218610 (.A(n_2028),
    .B(sa22[4]),
    .Y(n_2502));
 OR2x6_ASAP7_75t_SL g218611 (.A(n_2013),
    .B(n_1862),
    .Y(n_2500));
 NAND2xp5_ASAP7_75t_SL g218612 (.A(sa23[7]),
    .B(sa23[1]),
    .Y(n_1686));
 AND2x2_ASAP7_75t_SL g218613 (.A(n_1954),
    .B(sa02[1]),
    .Y(n_2497));
 AND2x4_ASAP7_75t_SL g218614 (.A(sa32[1]),
    .B(sa32[7]),
    .Y(n_2495));
 NAND2xp5_ASAP7_75t_L g218615 (.A(sa22[7]),
    .B(sa22[1]),
    .Y(n_2491));
 OR2x2_ASAP7_75t_SL g218616 (.A(n_8206),
    .B(n_8198),
    .Y(n_2490));
 NAND2x2_ASAP7_75t_SL g218617 (.A(sa10[7]),
    .B(sa10[1]),
    .Y(n_2488));
 AND2x2_ASAP7_75t_SL g218618 (.A(sa31[4]),
    .B(n_2008),
    .Y(n_2486));
 AND2x4_ASAP7_75t_SL g218619 (.A(n_1851),
    .B(n_2014),
    .Y(n_2484));
 AND2x4_ASAP7_75t_SL g218620 (.A(sa12[4]),
    .B(sa12[7]),
    .Y(n_2482));
 NAND2xp5_ASAP7_75t_SL g218621 (.A(sa31[7]),
    .B(sa31[1]),
    .Y(n_2479));
 AND2x2_ASAP7_75t_SL g218622 (.A(sa30[4]),
    .B(n_1900),
    .Y(n_2478));
 AND2x2_ASAP7_75t_SL g218623 (.A(sa21[7]),
    .B(sa21[4]),
    .Y(n_2476));
 AND2x4_ASAP7_75t_SL g218624 (.A(sa11[4]),
    .B(n_2018),
    .Y(n_2474));
 AND2x4_ASAP7_75t_SL g218625 (.A(n_1529),
    .B(n_1893),
    .Y(n_2472));
 AND2x4_ASAP7_75t_SL g218626 (.A(sa23[4]),
    .B(sa23[7]),
    .Y(n_2470));
 AND2x4_ASAP7_75t_SL g218627 (.A(n_1853),
    .B(n_1896),
    .Y(n_2468));
 NAND2x2_ASAP7_75t_SL g218628 (.A(n_1905),
    .B(n_2014),
    .Y(n_2466));
 AND2x4_ASAP7_75t_SL g218629 (.A(sa02[7]),
    .B(sa02[1]),
    .Y(n_2465));
 AND2x4_ASAP7_75t_SL g218630 (.A(sa12[1]),
    .B(sa12[7]),
    .Y(n_2463));
 AND2x2_ASAP7_75t_SL g218631 (.A(sa21[7]),
    .B(sa21[1]),
    .Y(n_2460));
 NAND2x1p5_ASAP7_75t_SL g218632 (.A(sa13[7]),
    .B(n_1472),
    .Y(n_2459));
 AND2x4_ASAP7_75t_SL g218633 (.A(sa03[4]),
    .B(n_1534),
    .Y(n_2457));
 NAND2x1_ASAP7_75t_SL g218634 (.A(sa30[1]),
    .B(n_1903),
    .Y(n_2455));
 AND2x4_ASAP7_75t_SL g218635 (.A(sa20[4]),
    .B(sa20[7]),
    .Y(n_2453));
 AND2x4_ASAP7_75t_SL g218636 (.A(sa13[7]),
    .B(n_1955),
    .Y(n_2451));
 AND2x4_ASAP7_75t_SL g218637 (.A(n_1910),
    .B(n_8899),
    .Y(n_2449));
 AND2x2_ASAP7_75t_SL g218638 (.A(sa01[1]),
    .B(sa01[7]),
    .Y(n_2447));
 NAND2xp5_ASAP7_75t_SL g218639 (.A(sa01[7]),
    .B(sa01[1]),
    .Y(n_1345));
 AND2x4_ASAP7_75t_SL g218640 (.A(sa03[1]),
    .B(sa03[7]),
    .Y(n_2445));
 AND2x2_ASAP7_75t_SL g218641 (.A(sa01[7]),
    .B(sa01[4]),
    .Y(n_2443));
 AND2x4_ASAP7_75t_SL g218642 (.A(n_2028),
    .B(sa22[4]),
    .Y(n_2441));
 OR2x6_ASAP7_75t_SL g218643 (.A(n_8212),
    .B(n_2010),
    .Y(n_2439));
 AND2x4_ASAP7_75t_SL g218644 (.A(sa10[7]),
    .B(sa10[4]),
    .Y(n_2437));
 AND2x2_ASAP7_75t_SL g218645 (.A(n_1843),
    .B(n_8210),
    .Y(n_2435));
 NOR2xp33_ASAP7_75t_L g218646 (.A(sa01[6]),
    .B(sa01[3]),
    .Y(n_2432));
 AND2x4_ASAP7_75t_SL g218647 (.A(n_1462),
    .B(n_1859),
    .Y(n_2431));
 OR2x2_ASAP7_75t_SL g218648 (.A(n_1935),
    .B(n_1972),
    .Y(n_1665));
 AND2x4_ASAP7_75t_SL g218649 (.A(n_1371),
    .B(n_8178),
    .Y(n_1664));
 AND2x2_ASAP7_75t_SL g218650 (.A(sa11[3]),
    .B(sa11[6]),
    .Y(n_1659));
 OR2x6_ASAP7_75t_SL g218651 (.A(sa22[6]),
    .B(sa22[3]),
    .Y(n_2428));
 OR2x4_ASAP7_75t_SL g218652 (.A(sa11[3]),
    .B(sa11[6]),
    .Y(n_1656));
 AND2x4_ASAP7_75t_SL g218653 (.A(n_8186),
    .B(n_1975),
    .Y(n_2425));
 OR2x2_ASAP7_75t_SL g218654 (.A(sa13[3]),
    .B(n_1934),
    .Y(n_2423));
 AND2x2_ASAP7_75t_L g218655 (.A(n_8195),
    .B(n_8211),
    .Y(n_2420));
 NAND2xp5_ASAP7_75t_L g218656 (.A(sa00[3]),
    .B(sa00[6]),
    .Y(n_2418));
 AND2x2_ASAP7_75t_SL g218657 (.A(sa00[3]),
    .B(sa00[6]),
    .Y(n_1653));
 AND2x2_ASAP7_75t_SL g218658 (.A(sa33[3]),
    .B(sa33[6]),
    .Y(n_2416));
 AND2x2_ASAP7_75t_SL g218659 (.A(n_1970),
    .B(n_1840),
    .Y(n_2413));
 NAND2x1_ASAP7_75t_SL g218660 (.A(n_1970),
    .B(n_1840),
    .Y(n_1651));
 OR2x2_ASAP7_75t_SL g218661 (.A(sa00[6]),
    .B(sa00[3]),
    .Y(n_2411));
 AND2x2_ASAP7_75t_SL g218662 (.A(n_1511),
    .B(sa12[6]),
    .Y(n_1351));
 AND2x4_ASAP7_75t_SL g218663 (.A(n_1979),
    .B(n_1839),
    .Y(n_2401));
 AND2x4_ASAP7_75t_SL g218664 (.A(sa02[6]),
    .B(n_1860),
    .Y(n_2400));
 AND2x2_ASAP7_75t_SL g218665 (.A(n_1984),
    .B(sa31[6]),
    .Y(n_1645));
 NOR2xp33_ASAP7_75t_R g218666 (.A(n_8181),
    .B(n_1933),
    .Y(n_2383));
 AND2x4_ASAP7_75t_SL g218667 (.A(sa22[3]),
    .B(sa22[6]),
    .Y(n_2397));
 OR2x6_ASAP7_75t_SL g218668 (.A(n_8178),
    .B(n_8180),
    .Y(n_2395));
 OR2x6_ASAP7_75t_SL g218669 (.A(n_8195),
    .B(n_8211),
    .Y(n_2393));
 AND2x2_ASAP7_75t_L g218670_220974 (.A(sa30[3]),
    .B(sa30[6]),
    .Y(n_1445));
 AND2x4_ASAP7_75t_SL g218672 (.A(sa01[3]),
    .B(sa01[6]),
    .Y(n_2389));
 OR2x2_ASAP7_75t_SL g218673 (.A(n_1859),
    .B(n_1462),
    .Y(n_1637));
 AND2x2_ASAP7_75t_SL g218674 (.A(n_8181),
    .B(n_1933),
    .Y(n_1636));
 AND2x4_ASAP7_75t_SL g218675 (.A(n_1933),
    .B(n_8181),
    .Y(n_2387));
 AND2x4_ASAP7_75t_SL g218676 (.A(sa21[3]),
    .B(sa21[6]),
    .Y(n_1350));
 AND2x2_ASAP7_75t_SL g218677 (.A(n_8177),
    .B(n_1938),
    .Y(n_2385));
 AND2x2_ASAP7_75t_SL g218678_0 (.A(n_1938),
    .B(n_8177),
    .Y(n_1622));
 INVxp33_ASAP7_75t_R g218679 (.A(n_2373),
    .Y(n_2374));
 INVxp33_ASAP7_75t_R g218680 (.A(n_2371),
    .Y(n_2372));
 INVxp33_ASAP7_75t_R g218681 (.A(n_2367),
    .Y(n_2368));
 INVxp33_ASAP7_75t_R g218682 (.A(n_2366),
    .Y(n_2365));
 INVxp33_ASAP7_75t_R g218683 (.A(n_2361),
    .Y(n_2362));
 INVxp33_ASAP7_75t_R g218684 (.A(n_2356),
    .Y(n_2357));
 INVxp33_ASAP7_75t_R g218685 (.A(n_2352),
    .Y(n_2351));
 INVxp67_ASAP7_75t_R g218686 (.A(n_2350),
    .Y(n_2349));
 INVxp33_ASAP7_75t_R g218689 (.A(n_1621),
    .Y(n_2345));
 INVxp33_ASAP7_75t_R g218690 (.A(n_2344),
    .Y(n_2343));
 INVxp33_ASAP7_75t_R g218691 (.A(n_2341),
    .Y(n_2340));
 INVxp33_ASAP7_75t_R g218692 (.A(n_2338),
    .Y(n_2339));
 INVxp67_ASAP7_75t_R g218693 (.A(n_2336),
    .Y(n_2337));
 INVxp33_ASAP7_75t_R g218694 (.A(n_2334),
    .Y(n_2335));
 INVxp33_ASAP7_75t_R g218695 (.A(n_1620),
    .Y(n_2333));
 INVxp67_ASAP7_75t_R g218697 (.A(n_2332),
    .Y(n_2331));
 INVxp67_ASAP7_75t_R g218698 (.A(n_2330),
    .Y(n_2329));
 INVxp33_ASAP7_75t_R g218699 (.A(n_2328),
    .Y(n_2327));
 INVx1_ASAP7_75t_L g218700 (.A(n_2326),
    .Y(n_2325));
 INVxp67_ASAP7_75t_R g218701 (.A(n_2324),
    .Y(n_2323));
 INVxp33_ASAP7_75t_R g218702 (.A(n_1619),
    .Y(n_2322));
 INVxp33_ASAP7_75t_R g218705 (.A(n_2320),
    .Y(n_2321));
 HB1xp67_ASAP7_75t_R g218706 (.A(n_2319),
    .Y(n_2320));
 INVxp67_ASAP7_75t_L g218707 (.A(n_2318),
    .Y(n_2317));
 INVxp33_ASAP7_75t_R g218708 (.A(n_2316),
    .Y(n_2315));
 INVxp33_ASAP7_75t_R g218709 (.A(n_2314),
    .Y(n_2313));
 INVxp67_ASAP7_75t_R g218710 (.A(n_2311),
    .Y(n_2312));
 INVxp33_ASAP7_75t_R g218711 (.A(n_2310),
    .Y(n_2309));
 INVxp67_ASAP7_75t_SL g218712 (.A(n_2308),
    .Y(n_2307));
 INVx1_ASAP7_75t_R g218713 (.A(n_2306),
    .Y(n_2305));
 INVxp67_ASAP7_75t_R g218714 (.A(n_2304),
    .Y(n_2303));
 INVxp33_ASAP7_75t_R g218715 (.A(n_2302),
    .Y(n_2301));
 INVxp33_ASAP7_75t_R g218716 (.A(n_1618),
    .Y(n_2300));
 INVxp33_ASAP7_75t_R g218719 (.A(n_1617),
    .Y(n_2298));
 INVxp67_ASAP7_75t_R g218720 (.A(n_2297),
    .Y(n_2296));
 INVxp67_ASAP7_75t_R g218721 (.A(n_2295),
    .Y(n_2294));
 INVx2_ASAP7_75t_SL g218722 (.A(n_2292),
    .Y(n_2291));
 INVxp67_ASAP7_75t_R g218723 (.A(n_2290),
    .Y(n_2289));
 INVxp33_ASAP7_75t_R g218724 (.A(n_1616),
    .Y(n_2288));
 HB1xp67_ASAP7_75t_L g218726 (.A(n_2287),
    .Y(n_1616));
 INVxp33_ASAP7_75t_R g218727 (.A(n_2286),
    .Y(n_2285));
 INVxp67_ASAP7_75t_R g218728 (.A(n_2284),
    .Y(n_2283));
 INVxp67_ASAP7_75t_R g218729 (.A(n_2282),
    .Y(n_2281));
 INVxp33_ASAP7_75t_R g218730 (.A(n_1615),
    .Y(n_2280));
 INVxp33_ASAP7_75t_R g218732 (.A(n_2279),
    .Y(n_2278));
 INVxp33_ASAP7_75t_R g218733 (.A(n_2277),
    .Y(n_2276));
 INVxp67_ASAP7_75t_R g218734 (.A(n_2275),
    .Y(n_2274));
 INVxp67_ASAP7_75t_R g218735 (.A(n_2273),
    .Y(n_2272));
 HB1xp67_ASAP7_75t_SL g218736 (.A(n_2270),
    .Y(n_2271));
 INVx1_ASAP7_75t_L g218737 (.A(n_2269),
    .Y(n_2270));
 INVx1_ASAP7_75t_L g218738 (.A(n_2268),
    .Y(n_2269));
 INVxp67_ASAP7_75t_R g218739 (.A(n_2267),
    .Y(n_2266));
 INVxp67_ASAP7_75t_R g218740 (.A(n_2265),
    .Y(n_2264));
 INVxp67_ASAP7_75t_L g218743 (.A(n_1613),
    .Y(n_1614));
 BUFx2_ASAP7_75t_SL g218744 (.A(n_2263),
    .Y(n_1613));
 INVxp67_ASAP7_75t_R g218745 (.A(n_2262),
    .Y(n_2261));
 INVxp33_ASAP7_75t_R g218746 (.A(n_2260),
    .Y(n_2259));
 INVxp33_ASAP7_75t_R g218747 (.A(n_2258),
    .Y(n_2257));
 INVx1_ASAP7_75t_SL g218748 (.A(n_2256),
    .Y(n_2255));
 INVxp67_ASAP7_75t_R g218753 (.A(n_1611),
    .Y(n_1612));
 INVx1_ASAP7_75t_L g218754 (.A(n_2254),
    .Y(n_1611));
 INVx2_ASAP7_75t_SL g218755 (.A(n_2253),
    .Y(n_2252));
 INVx1_ASAP7_75t_L g218756 (.A(n_2251),
    .Y(n_2250));
 INVxp33_ASAP7_75t_R g218757 (.A(n_2249),
    .Y(n_2248));
 INVx2_ASAP7_75t_SL g218760 (.A(n_2247),
    .Y(n_1610));
 INVxp33_ASAP7_75t_R g218763 (.A(n_1609),
    .Y(n_2246));
 INVxp67_ASAP7_75t_R g218765 (.A(n_2245),
    .Y(n_2244));
 INVx2_ASAP7_75t_L g218766 (.A(n_2243),
    .Y(n_2242));
 INVxp67_ASAP7_75t_L g218767 (.A(n_2241),
    .Y(n_2240));
 INVxp33_ASAP7_75t_R g218768 (.A(n_2239),
    .Y(n_2238));
 INVxp33_ASAP7_75t_R g218770 (.A(n_1608),
    .Y(n_2237));
 HB1xp67_ASAP7_75t_L g218772 (.A(n_2236),
    .Y(n_1608));
 INVxp33_ASAP7_75t_R g218773 (.A(n_2235),
    .Y(n_2234));
 INVxp33_ASAP7_75t_R g218774 (.A(n_2233),
    .Y(n_2232));
 INVx1_ASAP7_75t_L g218775 (.A(n_2231),
    .Y(n_2230));
 INVx1_ASAP7_75t_L g218776 (.A(n_2229),
    .Y(n_2228));
 INVx1_ASAP7_75t_SL g218777 (.A(n_2227),
    .Y(n_2226));
 INVxp67_ASAP7_75t_R g218778 (.A(n_2225),
    .Y(n_2224));
 INVx2_ASAP7_75t_SL g218779 (.A(n_2223),
    .Y(n_2222));
 INVx1_ASAP7_75t_SL g218780 (.A(n_2221),
    .Y(n_2220));
 INVx1_ASAP7_75t_L g218784 (.A(n_1606),
    .Y(n_1607));
 INVx2_ASAP7_75t_L g218785 (.A(n_2219),
    .Y(n_1606));
 INVx2_ASAP7_75t_SL g218786 (.A(n_2218),
    .Y(n_2219));
 INVxp67_ASAP7_75t_R g218787 (.A(n_2217),
    .Y(n_2216));
 INVx1_ASAP7_75t_SL g218788 (.A(n_2215),
    .Y(n_2214));
 INVxp33_ASAP7_75t_R g218794 (.A(n_1605),
    .Y(n_1604));
 INVx2_ASAP7_75t_SL g218795 (.A(n_2213),
    .Y(n_2212));
 INVxp67_ASAP7_75t_SL g218796 (.A(n_2211),
    .Y(n_2210));
 INVx1_ASAP7_75t_L g218797 (.A(n_2209),
    .Y(n_2208));
 INVx1_ASAP7_75t_L g218799 (.A(n_2205),
    .Y(n_2206));
 INVxp33_ASAP7_75t_R g218800 (.A(n_2204),
    .Y(n_2203));
 INVx1_ASAP7_75t_R g218801 (.A(n_2202),
    .Y(n_2201));
 INVxp67_ASAP7_75t_R g218802 (.A(n_2200),
    .Y(n_2199));
 INVxp67_ASAP7_75t_L g218804 (.A(n_2198),
    .Y(n_1603));
 INVx1_ASAP7_75t_L g218805 (.A(n_2197),
    .Y(n_2198));
 INVx1_ASAP7_75t_L g218806 (.A(n_2196),
    .Y(n_2195));
 INVxp33_ASAP7_75t_R g218807 (.A(n_2194),
    .Y(n_2193));
 INVxp67_ASAP7_75t_R g218808 (.A(n_2191),
    .Y(n_2190));
 INVxp33_ASAP7_75t_R g218809 (.A(n_2189),
    .Y(n_2188));
 INVx2_ASAP7_75t_SL g218810 (.A(n_2186),
    .Y(n_2185));
 INVxp67_ASAP7_75t_R g218811 (.A(n_2184),
    .Y(n_2183));
 INVxp33_ASAP7_75t_R g218812 (.A(n_2182),
    .Y(n_2181));
 INVx1_ASAP7_75t_R g218814 (.A(n_2180),
    .Y(n_2179));
 INVx1_ASAP7_75t_R g218816 (.A(n_2178),
    .Y(n_2177));
 HB1xp67_ASAP7_75t_SL g218817 (.A(n_2176),
    .Y(n_2178));
 INVxp67_ASAP7_75t_R g218818 (.A(n_2175),
    .Y(n_2174));
 INVxp67_ASAP7_75t_R g218819 (.A(n_2173),
    .Y(n_2172));
 INVx1_ASAP7_75t_L g218820 (.A(n_2171),
    .Y(n_2170));
 INVx1_ASAP7_75t_L g218821 (.A(n_2169),
    .Y(n_2168));
 INVx1_ASAP7_75t_L g218824 (.A(n_1602),
    .Y(n_2167));
 INVx1_ASAP7_75t_L g218825 (.A(n_2166),
    .Y(n_1602));
 INVx1_ASAP7_75t_SL g218826 (.A(n_2165),
    .Y(n_2166));
 INVx1_ASAP7_75t_R g218827 (.A(n_2164),
    .Y(n_2163));
 INVxp67_ASAP7_75t_L g218832 (.A(n_1601),
    .Y(n_1600));
 INVx1_ASAP7_75t_SL g218833 (.A(n_2162),
    .Y(n_1601));
 INVx2_ASAP7_75t_L g218834 (.A(n_2161),
    .Y(n_2162));
 INVx1_ASAP7_75t_L g218835 (.A(n_2160),
    .Y(n_2159));
 INVxp33_ASAP7_75t_R g218836 (.A(n_2158),
    .Y(n_2157));
 INVx1_ASAP7_75t_SL g218837 (.A(n_2156),
    .Y(n_2155));
 INVx2_ASAP7_75t_SL g218838 (.A(n_2154),
    .Y(n_2153));
 INVxp67_ASAP7_75t_R g218839 (.A(n_2152),
    .Y(n_2151));
 INVx1_ASAP7_75t_SL g218840 (.A(n_1598),
    .Y(n_2150));
 INVxp33_ASAP7_75t_R g218842 (.A(n_1599),
    .Y(n_2149));
 INVx1_ASAP7_75t_SL g218845 (.A(n_1598),
    .Y(n_1599));
 INVxp67_ASAP7_75t_L g218847 (.A(n_2147),
    .Y(n_2148));
 INVxp67_ASAP7_75t_R g218848 (.A(n_1597),
    .Y(n_2146));
 BUFx2_ASAP7_75t_SL g218849 (.A(n_2147),
    .Y(n_1597));
 HB1xp67_ASAP7_75t_SL g218850 (.A(n_2144),
    .Y(n_2147));
 INVx1_ASAP7_75t_SL g218851 (.A(n_2144),
    .Y(n_2145));
 INVx1_ASAP7_75t_R g218852 (.A(n_2143),
    .Y(n_2142));
 INVxp67_ASAP7_75t_R g218853 (.A(n_2141),
    .Y(n_2140));
 INVx1_ASAP7_75t_SL g218854 (.A(n_2139),
    .Y(n_2138));
 INVx3_ASAP7_75t_SL g218855 (.A(n_2137),
    .Y(n_2136));
 INVx1_ASAP7_75t_L g218856 (.A(n_2135),
    .Y(n_2134));
 INVx3_ASAP7_75t_SL g218857 (.A(n_2133),
    .Y(n_2132));
 INVxp67_ASAP7_75t_R g218858 (.A(n_2131),
    .Y(n_2130));
 INVx1_ASAP7_75t_L g218859 (.A(n_2129),
    .Y(n_2128));
 INVxp67_ASAP7_75t_R g218860 (.A(n_2127),
    .Y(n_2126));
 INVx1_ASAP7_75t_L g218861 (.A(n_2125),
    .Y(n_2124));
 INVx4_ASAP7_75t_SL g218862 (.A(n_2123),
    .Y(n_2122));
 INVxp67_ASAP7_75t_L g218863 (.A(n_2119),
    .Y(n_2121));
 INVx1_ASAP7_75t_L g218864 (.A(n_1596),
    .Y(n_2120));
 HB1xp67_ASAP7_75t_SL g218867 (.A(n_2119),
    .Y(n_1596));
 INVx1_ASAP7_75t_SL g218868 (.A(n_2112),
    .Y(n_2118));
 INVxp67_ASAP7_75t_L g218869 (.A(n_2116),
    .Y(n_2117));
 HB1xp67_ASAP7_75t_SL g218871 (.A(n_2114),
    .Y(n_2116));
 INVxp67_ASAP7_75t_L g218872 (.A(n_2114),
    .Y(n_2115));
 INVxp67_ASAP7_75t_SL g218873 (.A(n_2113),
    .Y(n_2114));
 INVx1_ASAP7_75t_SL g218874 (.A(n_2112),
    .Y(n_2113));
 INVx2_ASAP7_75t_SL g218875 (.A(n_2111),
    .Y(n_2110));
 INVxp33_ASAP7_75t_R g218880 (.A(n_1595),
    .Y(n_1594));
 INVx1_ASAP7_75t_L g218882 (.A(n_2108),
    .Y(n_2107));
 INVxp67_ASAP7_75t_R g218883 (.A(n_2106),
    .Y(n_2105));
 INVx3_ASAP7_75t_SL g218884 (.A(n_2104),
    .Y(n_2103));
 INVxp67_ASAP7_75t_R g218885 (.A(n_2102),
    .Y(n_2101));
 INVxp67_ASAP7_75t_R g218886 (.A(n_2100),
    .Y(n_2099));
 INVxp33_ASAP7_75t_R g218887 (.A(n_1593),
    .Y(n_2098));
 INVx1_ASAP7_75t_L g218891 (.A(n_1592),
    .Y(n_1593));
 BUFx3_ASAP7_75t_SL g218893 (.A(n_2097),
    .Y(n_1592));
 INVx1_ASAP7_75t_R g218894 (.A(n_2096),
    .Y(n_2095));
 INVx1_ASAP7_75t_L g218895 (.A(n_1591),
    .Y(n_2094));
 INVx3_ASAP7_75t_SL g218900 (.A(n_1337),
    .Y(n_2092));
 INVx2_ASAP7_75t_SL g218901 (.A(n_2091),
    .Y(n_2090));
 INVx4_ASAP7_75t_SL g218902 (.A(n_2089),
    .Y(n_2088));
 INVxp67_ASAP7_75t_R g218909 (.A(n_1588),
    .Y(n_2087));
 INVx1_ASAP7_75t_SL g218919 (.A(n_1590),
    .Y(n_1587));
 INVx3_ASAP7_75t_L g218920 (.A(n_1589),
    .Y(n_1590));
 INVx2_ASAP7_75t_SL g218925 (.A(n_1589),
    .Y(n_1588));
 INVx4_ASAP7_75t_SL g218926 (.A(n_2084),
    .Y(n_2083));
 INVx4_ASAP7_75t_SL g218927 (.A(n_2082),
    .Y(n_2081));
 INVx2_ASAP7_75t_SL g218942 (.A(n_2080),
    .Y(n_1586));
 INVx1_ASAP7_75t_L g218949 (.A(n_1585),
    .Y(n_1584));
 INVx1_ASAP7_75t_L g218951 (.A(n_2080),
    .Y(n_1585));
 INVx4_ASAP7_75t_SL g218952 (.A(n_2079),
    .Y(n_2078));
 BUFx2_ASAP7_75t_SL g218955 (.A(n_2076),
    .Y(n_2077));
 BUFx2_ASAP7_75t_SL g218959 (.A(n_1583),
    .Y(n_1582));
 INVx1_ASAP7_75t_SL g218972 (.A(n_1580),
    .Y(n_1581));
 INVx2_ASAP7_75t_SL g218974 (.A(n_1577),
    .Y(n_1580));
 INVx1_ASAP7_75t_R g218981 (.A(n_1577),
    .Y(n_1578));
 INVx3_ASAP7_75t_L g218985 (.A(n_2075),
    .Y(n_2074));
 INVx3_ASAP7_75t_SL g218986 (.A(n_2073),
    .Y(n_2072));
 INVx2_ASAP7_75t_SL g218990 (.A(n_1575),
    .Y(n_1576));
 INVx2_ASAP7_75t_SL g218994 (.A(n_1344),
    .Y(n_2069));
 BUFx3_ASAP7_75t_SL g218997 (.A(n_1575),
    .Y(n_1344));
 INVxp67_ASAP7_75t_R g218999 (.A(n_1576),
    .Y(n_2070));
 INVx4_ASAP7_75t_SL g219012 (.A(n_2068),
    .Y(n_2067));
 INVx3_ASAP7_75t_SL g219013 (.A(n_2066),
    .Y(n_2065));
 INVxp67_ASAP7_75t_L g219016 (.A(n_1572),
    .Y(n_1573));
 INVx2_ASAP7_75t_R g219027 (.A(n_1570),
    .Y(n_1571));
 INVx2_ASAP7_75t_SL g219028 (.A(n_1342),
    .Y(n_1570));
 INVx2_ASAP7_75t_SL g219033 (.A(n_1342),
    .Y(n_1572));
 INVx4_ASAP7_75t_SL g219036 (.A(n_2064),
    .Y(n_2063));
 INVx3_ASAP7_75t_SL g219037 (.A(n_2062),
    .Y(n_2061));
 INVx3_ASAP7_75t_SL g219054 (.A(n_1568),
    .Y(n_1349));
 INVx3_ASAP7_75t_SL g219055 (.A(n_1569),
    .Y(n_1568));
 INVx2_ASAP7_75t_L g219059 (.A(n_1567),
    .Y(n_1348));
 INVx3_ASAP7_75t_SL g219061 (.A(n_1569),
    .Y(n_1567));
 INVx2_ASAP7_75t_SL g219068 (.A(n_2060),
    .Y(n_2059));
 INVx2_ASAP7_75t_L g219069 (.A(n_2058),
    .Y(n_2057));
 INVx3_ASAP7_75t_L g219070 (.A(n_2056),
    .Y(n_2055));
 INVx4_ASAP7_75t_SL g219071 (.A(n_2054),
    .Y(n_2053));
 INVx2_ASAP7_75t_SL g219077 (.A(n_2052),
    .Y(n_2051));
 INVx2_ASAP7_75t_SL g219078 (.A(n_1566),
    .Y(n_2052));
 INVx1_ASAP7_75t_R g219090 (.A(n_1565),
    .Y(n_2050));
 INVx2_ASAP7_75t_L g219094 (.A(n_1566),
    .Y(n_1565));
 INVx3_ASAP7_75t_SL g219102 (.A(n_1560),
    .Y(n_1559));
 INVxp67_ASAP7_75t_SL g219109 (.A(n_1561),
    .Y(n_1562));
 INVx4_ASAP7_75t_SL g219117 (.A(n_1560),
    .Y(n_1561));
 INVx3_ASAP7_75t_SL g219119 (.A(n_2048),
    .Y(n_2047));
 INVx2_ASAP7_75t_SL g219123 (.A(n_1558),
    .Y(n_2046));
 INVx2_ASAP7_75t_SL g219131 (.A(n_1557),
    .Y(n_1558));
 INVxp33_ASAP7_75t_R g219136 (.A(n_1556),
    .Y(n_1555));
 INVx1_ASAP7_75t_L g219137 (.A(n_1557),
    .Y(n_1556));
 INVx2_ASAP7_75t_SL g219144 (.A(n_1554),
    .Y(n_1553));
 BUFx3_ASAP7_75t_SL g219146 (.A(n_1557),
    .Y(n_1554));
 INVx2_ASAP7_75t_SL g219147 (.A(n_2045),
    .Y(n_2044));
 INVx3_ASAP7_75t_SL g219148 (.A(n_2043),
    .Y(n_2042));
 INVx4_ASAP7_75t_SL g219154 (.A(n_1552),
    .Y(n_2041));
 INVx1_ASAP7_75t_L g219163 (.A(n_1551),
    .Y(n_1550));
 INVx2_ASAP7_75t_SL g219165 (.A(n_1552),
    .Y(n_1551));
 INVx2_ASAP7_75t_SL g219172 (.A(n_2041),
    .Y(n_1549));
 INVx2_ASAP7_75t_L g219184 (.A(n_1548),
    .Y(n_1547));
 INVx2_ASAP7_75t_L g219187 (.A(n_2040),
    .Y(n_1548));
 INVxp67_ASAP7_75t_L g219192 (.A(n_1546),
    .Y(n_2039));
 INVx2_ASAP7_75t_L g219197 (.A(n_2040),
    .Y(n_1546));
 INVx2_ASAP7_75t_L g219201 (.A(n_1544),
    .Y(n_1545));
 INVx2_ASAP7_75t_SL g219205 (.A(n_1542),
    .Y(n_1544));
 INVx1_ASAP7_75t_L g219209 (.A(n_1542),
    .Y(n_1541));
 INVx1_ASAP7_75t_SL g219213 (.A(n_1542),
    .Y(n_1543));
 NAND2xp33_ASAP7_75t_R g219219 (.A(sa23[5]),
    .B(n_1538),
    .Y(n_2038));
 NAND2xp33_ASAP7_75t_R g219220 (.A(n_2014),
    .B(n_1979),
    .Y(n_2382));
 NAND2xp33_ASAP7_75t_R g219221 (.A(sa30[5]),
    .B(n_1924),
    .Y(n_2381));
 NAND2xp33_ASAP7_75t_R g219222 (.A(sa02[7]),
    .B(n_8210),
    .Y(n_2380));
 NAND2xp33_ASAP7_75t_R g219223 (.A(sa20[7]),
    .B(n_1867),
    .Y(n_2379));
 NAND2xp5_ASAP7_75t_R g219224 (.A(n_8177),
    .B(n_1484),
    .Y(n_2378));
 NAND2xp33_ASAP7_75t_R g219225 (.A(n_1975),
    .B(sa21[7]),
    .Y(n_2377));
 NAND2xp33_ASAP7_75t_R g219226 (.A(n_1915),
    .B(sa01[5]),
    .Y(n_2376));
 NOR2xp33_ASAP7_75t_R g219227 (.A(sa22[2]),
    .B(n_1879),
    .Y(n_2375));
 NOR2xp33_ASAP7_75t_R g219228 (.A(n_2001),
    .B(n_1519),
    .Y(n_2373));
 NAND2xp33_ASAP7_75t_R g219229 (.A(sa10[4]),
    .B(n_8178),
    .Y(n_2371));
 NAND2xp5_ASAP7_75t_R g219230 (.A(n_1971),
    .B(sa12[4]),
    .Y(n_2370));
 NOR2xp33_ASAP7_75t_SL g219231 (.A(n_2034),
    .B(n_1913),
    .Y(n_2369));
 NAND2xp33_ASAP7_75t_R g219232 (.A(n_1387),
    .B(n_1986),
    .Y(n_2367));
 NAND2xp33_ASAP7_75t_R g219233 (.A(n_1967),
    .B(n_1425),
    .Y(n_2366));
 NAND2xp33_ASAP7_75t_R g219234 (.A(n_1954),
    .B(n_8210),
    .Y(n_2364));
 NAND2xp5_ASAP7_75t_R g219235 (.A(n_1878),
    .B(n_1494),
    .Y(n_2363));
 NAND2xp33_ASAP7_75t_R g219236 (.A(n_2022),
    .B(n_1533),
    .Y(n_2361));
 NAND2xp5_ASAP7_75t_R g219237 (.A(n_1491),
    .B(n_1507),
    .Y(n_2360));
 NAND2xp5_ASAP7_75t_R g219238 (.A(n_1912),
    .B(n_8199),
    .Y(n_2359));
 NOR2xp33_ASAP7_75t_R g219239 (.A(sa01[3]),
    .B(n_1384),
    .Y(n_2358));
 NOR2xp33_ASAP7_75t_R g219240 (.A(n_1361),
    .B(sa00[3]),
    .Y(n_2356));
 NAND2xp33_ASAP7_75t_R g219241 (.A(n_1506),
    .B(n_1518),
    .Y(n_2355));
 NAND2xp33_ASAP7_75t_R g219242 (.A(n_1851),
    .B(n_1979),
    .Y(n_2354));
 AND2x2_ASAP7_75t_R g219243 (.A(sa22[4]),
    .B(n_1985),
    .Y(n_2353));
 NAND2xp33_ASAP7_75t_R g219244 (.A(n_8181),
    .B(sa31[4]),
    .Y(n_2352));
 NAND2xp5_ASAP7_75t_R g219245 (.A(n_8177),
    .B(n_1375),
    .Y(n_2350));
 AND2x2_ASAP7_75t_R g219246 (.A(n_1862),
    .B(sa20[4]),
    .Y(n_2348));
 AND2x2_ASAP7_75t_R g219247 (.A(n_1975),
    .B(n_1947),
    .Y(n_2347));
 NAND2xp5_ASAP7_75t_R g219248 (.A(sa10[7]),
    .B(n_8178),
    .Y(n_2346));
 NAND2xp5_ASAP7_75t_L g219249 (.A(n_1507),
    .B(sa32[4]),
    .Y(n_1621));
 NOR2xp33_ASAP7_75t_R g219250 (.A(n_1950),
    .B(sa20[3]),
    .Y(n_2344));
 NOR2xp33_ASAP7_75t_R g219251 (.A(n_1914),
    .B(sa01[3]),
    .Y(n_2342));
 NOR2xp33_ASAP7_75t_R g219252 (.A(n_1856),
    .B(sa23[3]),
    .Y(n_2341));
 NAND2xp33_ASAP7_75t_R g219253 (.A(n_1534),
    .B(n_1967),
    .Y(n_2338));
 NOR2xp33_ASAP7_75t_L g219254 (.A(n_1535),
    .B(sa22[3]),
    .Y(n_2336));
 NAND2xp5_ASAP7_75t_R g219255 (.A(sa23[7]),
    .B(n_1983),
    .Y(n_2334));
 NAND2xp5_ASAP7_75t_SL g219256 (.A(n_1886),
    .B(n_1902),
    .Y(n_1620));
 AND2x2_ASAP7_75t_L g219257 (.A(n_1493),
    .B(n_1386),
    .Y(n_2332));
 NAND2xp5_ASAP7_75t_L g219258 (.A(n_1387),
    .B(n_1480),
    .Y(n_2330));
 OR2x2_ASAP7_75t_SL g219259 (.A(n_1918),
    .B(sa01[7]),
    .Y(n_2328));
 AND2x2_ASAP7_75t_SL g219260 (.A(sa03[1]),
    .B(n_2024),
    .Y(n_2326));
 NAND2xp5_ASAP7_75t_L g219261 (.A(n_1474),
    .B(n_1375),
    .Y(n_2324));
 NAND2xp5_ASAP7_75t_SL g219262 (.A(sa02[1]),
    .B(n_2010),
    .Y(n_1619));
 NAND2xp5_ASAP7_75t_SL g219263 (.A(sa12[1]),
    .B(n_2019),
    .Y(n_2319));
 OR2x2_ASAP7_75t_SL g219264 (.A(n_1995),
    .B(n_1910),
    .Y(n_2318));
 NAND2xp5_ASAP7_75t_L g219265 (.A(n_1853),
    .B(n_1477),
    .Y(n_2316));
 OR2x2_ASAP7_75t_L g219266 (.A(n_1523),
    .B(sa21[7]),
    .Y(n_2314));
 NOR2xp33_ASAP7_75t_L g219267 (.A(sa21[1]),
    .B(n_1939),
    .Y(n_2311));
 AND2x2_ASAP7_75t_R g219268 (.A(sa22[4]),
    .B(n_1471),
    .Y(n_2310));
 NOR2xp33_ASAP7_75t_SL g219269 (.A(n_1960),
    .B(sa10[1]),
    .Y(n_2308));
 AND2x2_ASAP7_75t_SL g219270 (.A(n_2020),
    .B(n_1425),
    .Y(n_2306));
 AND2x2_ASAP7_75t_L g219271 (.A(n_8204),
    .B(n_1851),
    .Y(n_2304));
 AND2x2_ASAP7_75t_SL g219272 (.A(n_8899),
    .B(n_1995),
    .Y(n_2302));
 NAND2xp5_ASAP7_75t_SL g219273 (.A(sa10[1]),
    .B(n_1921),
    .Y(n_1618));
 AND2x2_ASAP7_75t_SL g219274 (.A(n_1880),
    .B(n_1958),
    .Y(n_2299));
 NOR2x1_ASAP7_75t_SL g219275 (.A(n_1513),
    .B(sa23[7]),
    .Y(n_1617));
 NAND2xp5_ASAP7_75t_R g219276 (.A(n_1486),
    .B(sa31[4]),
    .Y(n_2297));
 OR2x2_ASAP7_75t_SL g219277 (.A(n_1469),
    .B(n_2028),
    .Y(n_2295));
 AND2x2_ASAP7_75t_SL g219278 (.A(n_1982),
    .B(n_1954),
    .Y(n_2293));
 AND2x2_ASAP7_75t_SL g219279 (.A(n_1487),
    .B(n_2007),
    .Y(n_2292));
 NAND2xp5_ASAP7_75t_L g219280 (.A(sa23[4]),
    .B(n_1513),
    .Y(n_2290));
 NAND2xp5_ASAP7_75t_SL g219281 (.A(n_1481),
    .B(n_2016),
    .Y(n_2287));
 OR2x2_ASAP7_75t_SL g219282 (.A(n_1862),
    .B(sa20[7]),
    .Y(n_2286));
 AND2x2_ASAP7_75t_L g219283 (.A(sa20[0]),
    .B(n_8179),
    .Y(n_2284));
 NAND2xp5_ASAP7_75t_R g219284 (.A(n_1987),
    .B(sa12[4]),
    .Y(n_2282));
 NAND2xp5_ASAP7_75t_SL g219285 (.A(n_1472),
    .B(n_2001),
    .Y(n_1615));
 OR2x2_ASAP7_75t_SL g219286 (.A(n_8204),
    .B(n_2014),
    .Y(n_2279));
 AND2x2_ASAP7_75t_SL g219287 (.A(sa03[2]),
    .B(n_8215),
    .Y(n_2277));
 OR2x2_ASAP7_75t_SL g219288 (.A(n_8189),
    .B(n_2014),
    .Y(n_2275));
 AND2x2_ASAP7_75t_R g219289 (.A(sa30[0]),
    .B(n_1924),
    .Y(n_2273));
 NAND2xp5_ASAP7_75t_SL g219290 (.A(sa30[4]),
    .B(n_1901),
    .Y(n_2268));
 AND2x2_ASAP7_75t_L g219291 (.A(n_1980),
    .B(n_1981),
    .Y(n_2267));
 NAND2xp5_ASAP7_75t_R g219292 (.A(sa33[0]),
    .B(n_1540),
    .Y(n_2265));
 NAND2xp5_ASAP7_75t_SL g219293 (.A(sa00[1]),
    .B(n_8206),
    .Y(n_2263));
 AND2x2_ASAP7_75t_R g219294 (.A(sa23[0]),
    .B(n_2031),
    .Y(n_2262));
 NAND2xp5_ASAP7_75t_L g219295 (.A(sa22[0]),
    .B(n_2026),
    .Y(n_2260));
 AND2x2_ASAP7_75t_L g219296 (.A(sa00[0]),
    .B(n_1531),
    .Y(n_2258));
 AND2x2_ASAP7_75t_SL g219297 (.A(n_1914),
    .B(sa01[4]),
    .Y(n_2256));
 NAND2xp5_ASAP7_75t_SL g219298 (.A(n_1853),
    .B(n_1482),
    .Y(n_2254));
 OR2x2_ASAP7_75t_SL g219299 (.A(n_1940),
    .B(sa21[7]),
    .Y(n_2253));
 AND2x2_ASAP7_75t_L g219300 (.A(sa32[2]),
    .B(n_8203),
    .Y(n_2251));
 AND2x2_ASAP7_75t_SL g219301 (.A(sa32[4]),
    .B(n_1490),
    .Y(n_2249));
 OR2x2_ASAP7_75t_SL g219302 (.A(n_1855),
    .B(sa22[7]),
    .Y(n_2247));
 NAND2xp5_ASAP7_75t_SL g219303 (.A(sa12[1]),
    .B(n_1953),
    .Y(n_1609));
 AND2x2_ASAP7_75t_R g219304 (.A(sa01[0]),
    .B(n_1915),
    .Y(n_2245));
 AND2x2_ASAP7_75t_SL g219305 (.A(sa31[4]),
    .B(n_2007),
    .Y(n_2243));
 OR2x2_ASAP7_75t_SL g219306 (.A(n_1891),
    .B(n_1853),
    .Y(n_2241));
 AND2x2_ASAP7_75t_R g219307 (.A(sa11[0]),
    .B(n_2005),
    .Y(n_2239));
 NOR2xp33_ASAP7_75t_SL g219308 (.A(sa12[0]),
    .B(n_8199),
    .Y(n_2236));
 AND2x2_ASAP7_75t_SL g219309 (.A(n_1954),
    .B(n_2010),
    .Y(n_2235));
 OR2x2_ASAP7_75t_SL g219310 (.A(n_8179),
    .B(sa20[0]),
    .Y(n_2233));
 AND2x2_ASAP7_75t_SL g219311 (.A(n_1506),
    .B(n_2001),
    .Y(n_2231));
 NAND2x1p5_ASAP7_75t_SL g219312 (.A(n_2023),
    .B(sa03[4]),
    .Y(n_2229));
 AND2x2_ASAP7_75t_SL g219313 (.A(sa11[4]),
    .B(n_2016),
    .Y(n_2227));
 OR2x2_ASAP7_75t_SL g219314 (.A(sa02[0]),
    .B(n_8208),
    .Y(n_2225));
 OR2x2_ASAP7_75t_SL g219315 (.A(n_1493),
    .B(n_1385),
    .Y(n_2223));
 NAND2xp5_ASAP7_75t_SL g219316 (.A(n_1966),
    .B(n_1494),
    .Y(n_2221));
 NAND2xp5_ASAP7_75t_SL g219317 (.A(n_1950),
    .B(sa20[7]),
    .Y(n_2218));
 AND2x2_ASAP7_75t_L g219318 (.A(n_1466),
    .B(n_1950),
    .Y(n_2217));
 OR2x2_ASAP7_75t_SL g219319 (.A(n_8205),
    .B(sa30[4]),
    .Y(n_2215));
 NAND2x1_ASAP7_75t_SL g219320 (.A(n_8212),
    .B(sa02[7]),
    .Y(n_1605));
 AND2x2_ASAP7_75t_SL g219321 (.A(sa10[4]),
    .B(n_1921),
    .Y(n_2213));
 NAND2x1p5_ASAP7_75t_SL g219322 (.A(n_1871),
    .B(sa10[7]),
    .Y(n_2211));
 AND2x2_ASAP7_75t_SL g219323 (.A(sa23[4]),
    .B(n_1916),
    .Y(n_2209));
 NAND2xp5_ASAP7_75t_SL g219324 (.A(sa32[7]),
    .B(n_8894),
    .Y(n_2205));
 NAND2x1_ASAP7_75t_SL g219325 (.A(sa22[2]),
    .B(n_8217),
    .Y(n_2204));
 AND2x2_ASAP7_75t_SL g219326 (.A(sa13[2]),
    .B(n_8188),
    .Y(n_2202));
 NAND2x1p5_ASAP7_75t_SL g219327 (.A(n_2014),
    .B(n_8204),
    .Y(n_2200));
 NAND2xp5_ASAP7_75t_SL g219328 (.A(n_1953),
    .B(sa12[7]),
    .Y(n_2197));
 OR2x2_ASAP7_75t_SL g219329 (.A(n_1953),
    .B(sa12[7]),
    .Y(n_2196));
 AND2x2_ASAP7_75t_SL g219330 (.A(sa23[1]),
    .B(n_1856),
    .Y(n_2194));
 OR2x2_ASAP7_75t_R g219331 (.A(n_1482),
    .B(n_1853),
    .Y(n_2192));
 AND2x2_ASAP7_75t_SL g219332 (.A(sa11[2]),
    .B(n_8182),
    .Y(n_2191));
 AND2x2_ASAP7_75t_SL g219333 (.A(sa30[2]),
    .B(n_1870),
    .Y(n_2189));
 AND2x2_ASAP7_75t_L g219334 (.A(n_1479),
    .B(n_1952),
    .Y(n_2187));
 OR2x2_ASAP7_75t_SL g219335 (.A(sa03[1]),
    .B(n_2024),
    .Y(n_2186));
 AND2x2_ASAP7_75t_SL g219336 (.A(sa00[2]),
    .B(n_8196),
    .Y(n_2184));
 AND2x2_ASAP7_75t_L g219337 (.A(sa20[4]),
    .B(n_2013),
    .Y(n_2182));
 AND2x2_ASAP7_75t_L g219338 (.A(n_1365),
    .B(n_8208),
    .Y(n_2180));
 NAND2xp5_ASAP7_75t_L g219339 (.A(sa13[7]),
    .B(n_1959),
    .Y(n_2176));
 AND2x2_ASAP7_75t_L g219340 (.A(n_1472),
    .B(n_1959),
    .Y(n_2175));
 AND2x2_ASAP7_75t_L g219341 (.A(n_1487),
    .B(n_1852),
    .Y(n_2173));
 NAND2xp5_ASAP7_75t_L g219342 (.A(sa01[7]),
    .B(n_1384),
    .Y(n_2171));
 OR2x2_ASAP7_75t_SL g219343 (.A(n_8187),
    .B(sa30[4]),
    .Y(n_2169));
 AND2x2_ASAP7_75t_SL g219344 (.A(n_2028),
    .B(n_1855),
    .Y(n_2165));
 OR2x2_ASAP7_75t_SL g219345 (.A(n_2032),
    .B(sa33[0]),
    .Y(n_2164));
 AND2x2_ASAP7_75t_SL g219346 (.A(n_2028),
    .B(n_1874),
    .Y(n_2161));
 AND2x2_ASAP7_75t_SL g219347 (.A(n_1856),
    .B(sa23[7]),
    .Y(n_2160));
 AND2x2_ASAP7_75t_SL g219348 (.A(n_1994),
    .B(n_8894),
    .Y(n_2158));
 NAND2xp5_ASAP7_75t_SL g219349 (.A(sa23[2]),
    .B(n_2012),
    .Y(n_2156));
 AND2x2_ASAP7_75t_SL g219350 (.A(sa01[7]),
    .B(n_1918),
    .Y(n_2154));
 AND2x2_ASAP7_75t_L g219351 (.A(sa01[2]),
    .B(n_1877),
    .Y(n_2152));
 NAND2x1_ASAP7_75t_SL g219352 (.A(n_8187),
    .B(n_1900),
    .Y(n_1598));
 NAND2xp5_ASAP7_75t_SL g219353 (.A(n_2008),
    .B(n_1486),
    .Y(n_2144));
 AND2x2_ASAP7_75t_L g219354 (.A(n_1522),
    .B(n_1502),
    .Y(n_2143));
 AND2x2_ASAP7_75t_SL g219355 (.A(n_1876),
    .B(n_1855),
    .Y(n_2141));
 NAND2x1p5_ASAP7_75t_SL g219356 (.A(sa23[7]),
    .B(n_1513),
    .Y(n_2139));
 AND2x4_ASAP7_75t_SL g219357 (.A(sa13[7]),
    .B(n_8192),
    .Y(n_2137));
 OR2x2_ASAP7_75t_SL g219358 (.A(sa21[1]),
    .B(n_2011),
    .Y(n_2135));
 AND2x4_ASAP7_75t_SL g219359 (.A(sa12[7]),
    .B(n_1987),
    .Y(n_2133));
 AND2x2_ASAP7_75t_L g219360 (.A(sa03[1]),
    .B(n_1948),
    .Y(n_2131));
 AND2x2_ASAP7_75t_R g219361 (.A(sa02[1]),
    .B(n_8212),
    .Y(n_2129));
 OR2x2_ASAP7_75t_L g219362 (.A(n_8204),
    .B(n_1851),
    .Y(n_2127));
 NAND2xp5_ASAP7_75t_SL g219363 (.A(n_1510),
    .B(n_1533),
    .Y(n_2125));
 AND2x4_ASAP7_75t_SL g219364 (.A(sa02[7]),
    .B(n_1982),
    .Y(n_2123));
 NAND2xp5_ASAP7_75t_SL g219365 (.A(sa21[7]),
    .B(n_1939),
    .Y(n_2119));
 NAND2xp5_ASAP7_75t_SL g219366 (.A(sa32[7]),
    .B(n_1990),
    .Y(n_2112));
 AND2x2_ASAP7_75t_SL g219367 (.A(n_1960),
    .B(sa10[7]),
    .Y(n_2111));
 OR2x2_ASAP7_75t_SL g219368 (.A(n_2023),
    .B(sa03[4]),
    .Y(n_1595));
 AND2x2_ASAP7_75t_SL g219369 (.A(n_8184),
    .B(n_2018),
    .Y(n_2108));
 AND2x2_ASAP7_75t_SL g219370 (.A(sa20[7]),
    .B(n_1862),
    .Y(n_2106));
 AND2x4_ASAP7_75t_SL g219371 (.A(n_2008),
    .B(n_1852),
    .Y(n_2104));
 AND2x2_ASAP7_75t_SL g219372 (.A(n_2014),
    .B(n_8189),
    .Y(n_2102));
 OR2x2_ASAP7_75t_L g219373 (.A(n_1871),
    .B(sa10[4]),
    .Y(n_2100));
 NAND2x1p5_ASAP7_75t_SL g219374 (.A(n_1896),
    .B(n_8198),
    .Y(n_2097));
 AND2x2_ASAP7_75t_SL g219375 (.A(n_1529),
    .B(n_1952),
    .Y(n_2096));
 NAND2xp5_ASAP7_75t_L g219376 (.A(sa12[0]),
    .B(n_8199),
    .Y(n_1591));
 OR2x6_ASAP7_75t_SL g219377 (.A(n_1972),
    .B(n_8180),
    .Y(n_1337));
 OR2x2_ASAP7_75t_SL g219378 (.A(sa32[3]),
    .B(n_8214),
    .Y(n_2091));
 AND2x4_ASAP7_75t_SL g219379 (.A(n_1930),
    .B(n_1967),
    .Y(n_2089));
 AND2x4_ASAP7_75t_SL g219380 (.A(n_1859),
    .B(sa01[6]),
    .Y(n_1589));
 AND2x4_ASAP7_75t_SL g219381 (.A(sa31[6]),
    .B(n_8181),
    .Y(n_2084));
 AND2x4_ASAP7_75t_SL g219382 (.A(n_1985),
    .B(sa22[6]),
    .Y(n_2082));
 OR2x4_ASAP7_75t_SL g219383 (.A(n_8211),
    .B(sa13[3]),
    .Y(n_2080));
 AND2x4_ASAP7_75t_SL g219384 (.A(sa30[6]),
    .B(n_8177),
    .Y(n_2079));
 AND2x2_ASAP7_75t_L g219385 (.A(n_1511),
    .B(n_1840),
    .Y(n_2076));
 OR2x2_ASAP7_75t_SL g219386 (.A(n_1970),
    .B(sa12[6]),
    .Y(n_1583));
 AND2x4_ASAP7_75t_SL g219387 (.A(sa33[6]),
    .B(n_1979),
    .Y(n_1577));
 AND2x4_ASAP7_75t_SL g219388 (.A(sa02[6]),
    .B(n_8210),
    .Y(n_2075));
 OR2x4_ASAP7_75t_SL g219389 (.A(n_8186),
    .B(sa21[3]),
    .Y(n_2073));
 OR2x2_ASAP7_75t_SL g219390 (.A(sa11[3]),
    .B(n_1850),
    .Y(n_1575));
 OR2x6_ASAP7_75t_L g219391 (.A(n_8210),
    .B(sa02[6]),
    .Y(n_2068));
 OR2x6_ASAP7_75t_SL g219392 (.A(n_1930),
    .B(sa03[3]),
    .Y(n_2066));
 AND2x4_ASAP7_75t_L g219394 (.A(sa12[6]),
    .B(n_1969),
    .Y(n_2064));
 AND2x4_ASAP7_75t_SL g219395 (.A(sa33[3]),
    .B(n_1839),
    .Y(n_2062));
 AND2x2_ASAP7_75t_SL g219396 (.A(n_1961),
    .B(n_8214),
    .Y(n_1569));
 AND2x4_ASAP7_75t_SL g219397 (.A(sa13[3]),
    .B(n_8211),
    .Y(n_2060));
 AND2x4_ASAP7_75t_SL g219398 (.A(sa01[3]),
    .B(n_1462),
    .Y(n_2058));
 OR2x6_ASAP7_75t_SL g219399 (.A(n_1467),
    .B(sa00[6]),
    .Y(n_2056));
 AND2x4_ASAP7_75t_SL g219400 (.A(sa22[3]),
    .B(n_1844),
    .Y(n_2054));
 NOR2xp33_ASAP7_75t_R g219401 (.A(n_1961),
    .B(n_8214),
    .Y(n_2037));
 AND2x4_ASAP7_75t_SL g219402 (.A(n_1964),
    .B(sa32[6]),
    .Y(n_1566));
 OR2x4_ASAP7_75t_SL g219403 (.A(sa32[6]),
    .B(n_1961),
    .Y(n_1560));
 AND2x4_ASAP7_75t_SL g219404 (.A(sa03[3]),
    .B(n_1929),
    .Y(n_2048));
 AND2x2_ASAP7_75t_SL g219405 (.A(sa03[3]),
    .B(n_1930),
    .Y(n_1557));
 OR2x2_ASAP7_75t_SL g219406 (.A(n_1986),
    .B(sa11[6]),
    .Y(n_2045));
 OR2x6_ASAP7_75t_SL g219407 (.A(n_8177),
    .B(sa30[6]),
    .Y(n_2043));
 AND2x2_ASAP7_75t_SL g219408 (.A(n_1972),
    .B(n_8180),
    .Y(n_1552));
 AND2x4_ASAP7_75t_SL g219409 (.A(n_1984),
    .B(n_1933),
    .Y(n_2040));
 INVxp33_ASAP7_75t_R g219412 (.A(w0[14]),
    .Y(n_2035));
 INVx2_ASAP7_75t_L g219413 (.A(n_8208),
    .Y(n_2034));
 INVx1_ASAP7_75t_L g219414 (.A(sa30[5]),
    .Y(n_2033));
 INVx2_ASAP7_75t_L g219425 (.A(sa33[2]),
    .Y(n_1540));
 INVx1_ASAP7_75t_SL g219426 (.A(sa33[2]),
    .Y(n_2032));
 INVxp33_ASAP7_75t_R g219427 (.A(sa23[2]),
    .Y(n_2031));
 INVx1_ASAP7_75t_SL g219433 (.A(n_1537),
    .Y(n_1538));
 HB1xp67_ASAP7_75t_SL g219434 (.A(sa23[2]),
    .Y(n_1537));
 INVx2_ASAP7_75t_SL g219435 (.A(n_2029),
    .Y(n_2028));
 INVxp67_ASAP7_75t_R g219439 (.A(n_1535),
    .Y(n_1536));
 HB1xp67_ASAP7_75t_L g219441 (.A(n_2029),
    .Y(n_1535));
 INVx3_ASAP7_75t_SL g219445 (.A(sa22[7]),
    .Y(n_2029));
 INVx1_ASAP7_75t_L g219446 (.A(sa22[2]),
    .Y(n_2026));
 INVx2_ASAP7_75t_SL g219448 (.A(sa03[7]),
    .Y(n_2024));
 INVx2_ASAP7_75t_SL g219455 (.A(n_2023),
    .Y(n_1534));
 INVx2_ASAP7_75t_SL g219457 (.A(sa03[7]),
    .Y(n_2023));
 INVx2_ASAP7_75t_R g219458 (.A(n_8197),
    .Y(n_2022));
 INVx1_ASAP7_75t_L g219467 (.A(n_1532),
    .Y(n_1533));
 BUFx2_ASAP7_75t_SL g219469 (.A(sa03[2]),
    .Y(n_1532));
 INVx1_ASAP7_75t_SL g219478 (.A(sa00[2]),
    .Y(n_1531));
 INVx1_ASAP7_75t_L g219479 (.A(sa03[1]),
    .Y(n_2020));
 INVx2_ASAP7_75t_R g219480 (.A(sa12[7]),
    .Y(n_2019));
 INVx1_ASAP7_75t_SL g219481 (.A(n_2017),
    .Y(n_2018));
 INVxp67_ASAP7_75t_SL g219482 (.A(sa11[7]),
    .Y(n_2017));
 INVxp67_ASAP7_75t_L g219487 (.A(n_2015),
    .Y(n_1530));
 HB1xp67_ASAP7_75t_SL g219488 (.A(n_1529),
    .Y(n_2015));
 INVx1_ASAP7_75t_SL g219490 (.A(n_1529),
    .Y(n_2016));
 BUFx3_ASAP7_75t_SL g219491 (.A(sa11[7]),
    .Y(n_1529));
 INVx4_ASAP7_75t_SL g219492 (.A(n_8191),
    .Y(n_2014));
 INVx1_ASAP7_75t_L g219497 (.A(n_1528),
    .Y(n_1527));
 BUFx2_ASAP7_75t_L g219503 (.A(sa10[0]),
    .Y(n_1528));
 INVx4_ASAP7_75t_SL g219504 (.A(sa20[7]),
    .Y(n_2013));
 INVx1_ASAP7_75t_L g219505 (.A(sa23[0]),
    .Y(n_2012));
 INVx2_ASAP7_75t_SL g219506 (.A(sa21[7]),
    .Y(n_2011));
 INVx4_ASAP7_75t_SL g219507 (.A(sa02[7]),
    .Y(n_2010));
 INVx1_ASAP7_75t_R g219508 (.A(sa23[5]),
    .Y(n_2009));
 INVx2_ASAP7_75t_L g219514 (.A(n_1526),
    .Y(n_1525));
 BUFx2_ASAP7_75t_SL g219515 (.A(n_2007),
    .Y(n_1526));
 INVx2_ASAP7_75t_SL g219516 (.A(n_2008),
    .Y(n_2007));
 INVx1_ASAP7_75t_SL g219518 (.A(n_2008),
    .Y(n_2006));
 BUFx3_ASAP7_75t_SL g219519 (.A(sa31[7]),
    .Y(n_2008));
 INVx1_ASAP7_75t_L g219520 (.A(sa11[2]),
    .Y(n_2005));
 INVxp33_ASAP7_75t_R g219521 (.A(sa10[5]),
    .Y(n_2004));
 INVx1_ASAP7_75t_L g219522 (.A(sa33[5]),
    .Y(n_2003));
 INVx4_ASAP7_75t_SL g219524 (.A(sa13[7]),
    .Y(n_2001));
 INVx2_ASAP7_75t_SL g219527 (.A(n_1995),
    .Y(n_1994));
 INVx1_ASAP7_75t_SL g219530 (.A(n_1524),
    .Y(n_1992));
 BUFx2_ASAP7_75t_SL g219534 (.A(n_1994),
    .Y(n_1524));
 INVx3_ASAP7_75t_SL g219536 (.A(sa32[1]),
    .Y(n_1995));
 INVx2_ASAP7_75t_SL g219537 (.A(sa32[1]),
    .Y(n_1990));
 INVx2_ASAP7_75t_L g219549 (.A(n_1523),
    .Y(n_1522));
 INVx2_ASAP7_75t_SL g219550 (.A(sa21[1]),
    .Y(n_1523));
 INVx4_ASAP7_75t_SL g219551 (.A(sa12[1]),
    .Y(n_1987));
 INVx3_ASAP7_75t_SL g219555 (.A(sa11[3]),
    .Y(n_1986));
 INVx3_ASAP7_75t_SL g219562 (.A(sa22[3]),
    .Y(n_1985));
 INVx4_ASAP7_75t_SL g219563 (.A(n_8181),
    .Y(n_1984));
 INVx2_ASAP7_75t_SL g219564 (.A(sa23[3]),
    .Y(n_1983));
 INVx4_ASAP7_75t_SL g219565 (.A(sa02[1]),
    .Y(n_1982));
 INVx2_ASAP7_75t_R g219566 (.A(sa32[2]),
    .Y(n_1981));
 INVx3_ASAP7_75t_SL g219567 (.A(n_8203),
    .Y(n_1980));
 INVx3_ASAP7_75t_SL g219568 (.A(sa33[3]),
    .Y(n_1979));
 INVx1_ASAP7_75t_SL g219581 (.A(n_1518),
    .Y(n_1519));
 INVx2_ASAP7_75t_SL g219582 (.A(sa13[3]),
    .Y(n_1518));
 INVx4_ASAP7_75t_SL g219585 (.A(sa21[3]),
    .Y(n_1975));
 INVx1_ASAP7_75t_SL g219589 (.A(n_1513),
    .Y(n_1517));
 INVx4_ASAP7_75t_SL g219602 (.A(sa23[1]),
    .Y(n_1513));
 INVx4_ASAP7_75t_SL g219603 (.A(n_8178),
    .Y(n_1972));
 INVx2_ASAP7_75t_SL g219612 (.A(n_1971),
    .Y(n_1512));
 BUFx2_ASAP7_75t_L g219613 (.A(n_1970),
    .Y(n_1971));
 INVx1_ASAP7_75t_SL g219614 (.A(sa12[3]),
    .Y(n_1970));
 INVx1_ASAP7_75t_SL g219616 (.A(n_1969),
    .Y(n_1511));
 INVx2_ASAP7_75t_SL g219617 (.A(sa12[3]),
    .Y(n_1969));
 INVx1_ASAP7_75t_L g219618 (.A(sa21[0]),
    .Y(n_1968));
 INVx2_ASAP7_75t_L g219630 (.A(n_1510),
    .Y(n_1509));
 INVx2_ASAP7_75t_SL g219631 (.A(n_8215),
    .Y(n_1510));
 INVx3_ASAP7_75t_SL g219632 (.A(sa03[3]),
    .Y(n_1967));
 INVx3_ASAP7_75t_SL g219633 (.A(n_8188),
    .Y(n_1966));
 INVxp67_ASAP7_75t_R g219634 (.A(sa12[0]),
    .Y(n_1965));
 INVxp67_ASAP7_75t_SL g219635 (.A(n_1961),
    .Y(n_1964));
 INVx2_ASAP7_75t_R g219643 (.A(n_1507),
    .Y(n_1343));
 BUFx2_ASAP7_75t_SL g219644 (.A(n_1961),
    .Y(n_1507));
 INVx2_ASAP7_75t_SL g219645 (.A(sa32[3]),
    .Y(n_1961));
 INVx4_ASAP7_75t_SL g219647 (.A(sa10[4]),
    .Y(n_1960));
 INVxp67_ASAP7_75t_SL g219657 (.A(n_1505),
    .Y(n_1504));
 INVx2_ASAP7_75t_R g219658 (.A(n_1506),
    .Y(n_1505));
 INVx3_ASAP7_75t_SL g219659 (.A(n_1959),
    .Y(n_1506));
 INVx1_ASAP7_75t_R g219660 (.A(n_1959),
    .Y(n_1958));
 INVxp67_ASAP7_75t_SL g219661 (.A(n_1955),
    .Y(n_1957));
 INVx2_ASAP7_75t_SL g219664 (.A(n_1959),
    .Y(n_1955));
 INVx4_ASAP7_75t_SL g219665 (.A(n_8212),
    .Y(n_1954));
 INVx5_ASAP7_75t_SL g219666 (.A(sa12[4]),
    .Y(n_1953));
 INVx3_ASAP7_75t_L g219667 (.A(sa11[4]),
    .Y(n_1952));
 INVx4_ASAP7_75t_SL g219668 (.A(sa01[4]),
    .Y(n_1384));
 INVx4_ASAP7_75t_SL g219669 (.A(sa20[4]),
    .Y(n_1950));
 INVx2_ASAP7_75t_L g219670 (.A(sa30[4]),
    .Y(n_1949));
 INVx2_ASAP7_75t_SL g219671 (.A(sa03[4]),
    .Y(n_1948));
 INVx1_ASAP7_75t_R g219672 (.A(n_1939),
    .Y(n_1947));
 INVx1_ASAP7_75t_SL g219675 (.A(n_1945),
    .Y(n_1944));
 BUFx2_ASAP7_75t_SL g219677 (.A(sa21[4]),
    .Y(n_1945));
 INVx1_ASAP7_75t_L g219682 (.A(n_1502),
    .Y(n_1503));
 INVx1_ASAP7_75t_SL g219685 (.A(sa21[4]),
    .Y(n_1502));
 INVx2_ASAP7_75t_SL g219687 (.A(n_1940),
    .Y(n_1941));
 BUFx3_ASAP7_75t_SL g219690 (.A(n_1939),
    .Y(n_1940));
 INVx3_ASAP7_75t_SL g219691 (.A(sa21[4]),
    .Y(n_1939));
 INVx3_ASAP7_75t_SL g219692 (.A(sa30[6]),
    .Y(n_1938));
 INVx1_ASAP7_75t_L g219697 (.A(n_1501),
    .Y(n_1336));
 INVx1_ASAP7_75t_R g219707 (.A(n_1501),
    .Y(n_1500));
 BUFx2_ASAP7_75t_L g219709 (.A(n_8186),
    .Y(n_1501));
 INVx5_ASAP7_75t_SL g219711 (.A(n_8180),
    .Y(n_1935));
 INVx2_ASAP7_75t_SL g219712 (.A(n_8211),
    .Y(n_1934));
 INVx4_ASAP7_75t_SL g219713 (.A(sa31[6]),
    .Y(n_1933));
 INVx2_ASAP7_75t_SL g219727 (.A(n_1499),
    .Y(n_1498));
 BUFx2_ASAP7_75t_SL g219730 (.A(n_8214),
    .Y(n_1499));
 INVx2_ASAP7_75t_L g219751 (.A(n_1497),
    .Y(n_1496));
 BUFx3_ASAP7_75t_SL g219752 (.A(n_1930),
    .Y(n_1497));
 INVx3_ASAP7_75t_SL g219753 (.A(n_1929),
    .Y(n_1930));
 INVx2_ASAP7_75t_SL g219755 (.A(sa03[6]),
    .Y(n_1929));
 INVxp33_ASAP7_75t_R g219756 (.A(dcnt[0]),
    .Y(n_1928));
 INVx1_ASAP7_75t_L g219758 (.A(sa31[2]),
    .Y(n_1926));
 INVx1_ASAP7_75t_L g219759 (.A(sa21[2]),
    .Y(n_1925));
 INVx1_ASAP7_75t_R g219760 (.A(sa30[2]),
    .Y(n_1924));
 INVx2_ASAP7_75t_SL g219761 (.A(n_8179),
    .Y(n_1923));
 INVx1_ASAP7_75t_SL g219771 (.A(n_1495),
    .Y(n_1494));
 BUFx3_ASAP7_75t_SL g219772 (.A(sa13[2]),
    .Y(n_1495));
 INVx2_ASAP7_75t_SL g219774 (.A(sa10[7]),
    .Y(n_1921));
 INVx1_ASAP7_75t_SL g219782 (.A(n_1493),
    .Y(n_1492));
 INVx1_ASAP7_75t_SL g219784 (.A(sa01[1]),
    .Y(n_1493));
 INVx2_ASAP7_75t_SL g219785 (.A(sa01[1]),
    .Y(n_1918));
 INVx2_ASAP7_75t_L g219786 (.A(sa20[5]),
    .Y(n_1917));
 INVx3_ASAP7_75t_SL g219787 (.A(sa23[7]),
    .Y(n_1916));
 INVx1_ASAP7_75t_R g219788 (.A(sa01[2]),
    .Y(n_1915));
 INVx1_ASAP7_75t_SL g219789 (.A(sa01[7]),
    .Y(n_1914));
 INVx1_ASAP7_75t_SL g219790 (.A(sa02[5]),
    .Y(n_1913));
 INVx1_ASAP7_75t_L g219791 (.A(n_8190),
    .Y(n_1912));
 BUFx3_ASAP7_75t_SL g219793 (.A(sa32[7]),
    .Y(n_1910));
 INVxp67_ASAP7_75t_SL g219794 (.A(sa32[7]),
    .Y(n_1909));
 INVx2_ASAP7_75t_SL g219795 (.A(sa32[7]),
    .Y(n_1908));
 INVx1_ASAP7_75t_L g219801 (.A(n_1490),
    .Y(n_1491));
 INVxp67_ASAP7_75t_SL g219804 (.A(sa32[7]),
    .Y(n_1490));
 INVx3_ASAP7_75t_SL g219805 (.A(n_8204),
    .Y(n_1905));
 INVxp33_ASAP7_75t_R g219810 (.A(n_1487),
    .Y(n_1904));
 INVx3_ASAP7_75t_SL g219815 (.A(sa31[1]),
    .Y(n_1486));
 INVx2_ASAP7_75t_SL g219819 (.A(n_1486),
    .Y(n_1487));
 INVx2_ASAP7_75t_SL g219822 (.A(n_8205),
    .Y(n_1903));
 HB1xp67_ASAP7_75t_SL g219823 (.A(n_8205),
    .Y(n_1902));
 INVx1_ASAP7_75t_L g219828 (.A(n_1485),
    .Y(n_1484));
 BUFx2_ASAP7_75t_SL g219829 (.A(n_1901),
    .Y(n_1485));
 INVxp67_ASAP7_75t_SL g219830 (.A(n_1900),
    .Y(n_1901));
 INVx2_ASAP7_75t_SL g219831 (.A(n_8205),
    .Y(n_1900));
 INVx5_ASAP7_75t_SL g219832 (.A(n_8206),
    .Y(n_1896));
 INVxp67_ASAP7_75t_R g219838 (.A(n_1482),
    .Y(n_1483));
 INVx2_ASAP7_75t_SL g219840 (.A(n_1896),
    .Y(n_1482));
 INVx1_ASAP7_75t_R g219842 (.A(sa31[5]),
    .Y(n_1895));
 INVxp33_ASAP7_75t_R g219843 (.A(n_1481),
    .Y(n_1894));
 INVxp67_ASAP7_75t_L g219845 (.A(n_8184),
    .Y(n_1481));
 INVx2_ASAP7_75t_SL g219851 (.A(n_1479),
    .Y(n_1480));
 INVx2_ASAP7_75t_L g219853 (.A(n_8184),
    .Y(n_1479));
 INVx1_ASAP7_75t_L g219854 (.A(n_8184),
    .Y(n_1893));
 INVxp67_ASAP7_75t_R g219856 (.A(n_1891),
    .Y(n_1890));
 BUFx2_ASAP7_75t_L g219857 (.A(n_8198),
    .Y(n_1891));
 INVx1_ASAP7_75t_SL g219863 (.A(n_1478),
    .Y(n_1477));
 INVx2_ASAP7_75t_SL g219864 (.A(n_8198),
    .Y(n_1478));
 INVx1_ASAP7_75t_R g219865 (.A(sa20[0]),
    .Y(n_1888));
 INVx1_ASAP7_75t_SL g219870 (.A(n_1475),
    .Y(n_1476));
 BUFx2_ASAP7_75t_SL g219874 (.A(n_8187),
    .Y(n_1475));
 INVx1_ASAP7_75t_SL g219875 (.A(n_8187),
    .Y(n_1886));
 INVx1_ASAP7_75t_R g219877 (.A(n_1886),
    .Y(n_1474));
 INVx1_ASAP7_75t_R g219880 (.A(sa01[5]),
    .Y(n_1884));
 INVx2_ASAP7_75t_SL g219888 (.A(n_1880),
    .Y(n_1473));
 BUFx3_ASAP7_75t_SL g219891 (.A(n_8192),
    .Y(n_1880));
 INVx2_ASAP7_75t_SL g219893 (.A(n_8192),
    .Y(n_1472));
 INVx1_ASAP7_75t_L g219894 (.A(sa22[5]),
    .Y(n_1879));
 INVx1_ASAP7_75t_L g219895 (.A(n_8207),
    .Y(n_1878));
 INVx1_ASAP7_75t_SL g219896 (.A(sa01[0]),
    .Y(n_1877));
 INVx1_ASAP7_75t_SL g219902 (.A(n_1471),
    .Y(n_1470));
 INVx2_ASAP7_75t_SL g219903 (.A(sa22[1]),
    .Y(n_1471));
 INVxp67_ASAP7_75t_L g219905 (.A(n_1469),
    .Y(n_1876));
 INVxp67_ASAP7_75t_SL g219906 (.A(sa22[1]),
    .Y(n_1469));
 INVx2_ASAP7_75t_SL g219908 (.A(sa22[1]),
    .Y(n_1874));
 INVx2_ASAP7_75t_L g219909 (.A(sa32[5]),
    .Y(n_1873));
 INVx3_ASAP7_75t_SL g219911 (.A(sa10[1]),
    .Y(n_1871));
 INVx1_ASAP7_75t_SL g219912 (.A(sa30[0]),
    .Y(n_1870));
 INVx1_ASAP7_75t_R g219913 (.A(sa33[0]),
    .Y(n_1869));
 INVx3_ASAP7_75t_SL g219922 (.A(sa00[3]),
    .Y(n_1467));
 INVx4_ASAP7_75t_SL g219924 (.A(sa20[3]),
    .Y(n_1867));
 INVx3_ASAP7_75t_SL g219925 (.A(n_8213),
    .Y(n_1866));
 INVx1_ASAP7_75t_L g219926 (.A(n_8209),
    .Y(n_1865));
 INVx2_ASAP7_75t_SL g219936 (.A(n_1862),
    .Y(n_1466));
 INVx3_ASAP7_75t_SL g219947 (.A(n_8210),
    .Y(n_1860));
 INVx3_ASAP7_75t_SL g219948 (.A(sa01[3]),
    .Y(n_1859));
 INVx1_ASAP7_75t_R g219950 (.A(sa02[0]),
    .Y(n_1857));
 INVx6_ASAP7_75t_SL g219951 (.A(sa23[4]),
    .Y(n_1856));
 INVx5_ASAP7_75t_SL g219952 (.A(sa22[4]),
    .Y(n_1855));
 INVx5_ASAP7_75t_SL g219954 (.A(n_8200),
    .Y(n_1853));
 INVx5_ASAP7_75t_SL g219955 (.A(sa31[4]),
    .Y(n_1852));
 INVx4_ASAP7_75t_SL g219956 (.A(n_8189),
    .Y(n_1851));
 INVx4_ASAP7_75t_SL g219957 (.A(sa11[6]),
    .Y(n_1850));
 INVx1_ASAP7_75t_R g219963 (.A(n_1464),
    .Y(n_1465));
 INVx1_ASAP7_75t_R g219979 (.A(n_1464),
    .Y(n_1463));
 INVx2_ASAP7_75t_L g219982 (.A(sa01[6]),
    .Y(n_1464));
 INVx2_ASAP7_75t_SL g219984 (.A(sa01[6]),
    .Y(n_1462));
 INVx1_ASAP7_75t_L g219985 (.A(sa00[6]),
    .Y(n_1846));
 INVx1_ASAP7_75t_R g219987 (.A(n_1461),
    .Y(n_1845));
 INVxp67_ASAP7_75t_SL g219997 (.A(n_1461),
    .Y(n_1460));
 BUFx2_ASAP7_75t_L g220004 (.A(sa00[6]),
    .Y(n_1461));
 INVx3_ASAP7_75t_SL g220005 (.A(sa22[6]),
    .Y(n_1844));
 INVxp67_ASAP7_75t_R g220006 (.A(sa02[6]),
    .Y(n_1843));
 INVx1_ASAP7_75t_L g220017 (.A(n_1458),
    .Y(n_1459));
 INVx1_ASAP7_75t_L g220025 (.A(n_1458),
    .Y(n_1457));
 BUFx2_ASAP7_75t_L g220031 (.A(sa02[6]),
    .Y(n_1458));
 INVx2_ASAP7_75t_L g220052 (.A(n_1456),
    .Y(n_1454));
 INVx1_ASAP7_75t_SL g220053 (.A(n_1455),
    .Y(n_1456));
 BUFx3_ASAP7_75t_SL g220054 (.A(sa12[6]),
    .Y(n_1455));
 INVx1_ASAP7_75t_SL g220056 (.A(sa12[6]),
    .Y(n_1840));
 INVx3_ASAP7_75t_SL g220058 (.A(sa33[6]),
    .Y(n_1839));
 AND2x2_ASAP7_75t_L g220848 (.A(sa30[3]),
    .B(sa30[6]),
    .Y(n_1641));
 AND2x2_ASAP7_75t_SL g220868 (.A(n_1938),
    .B(n_8177),
    .Y(n_1625));
 AND2x4_ASAP7_75t_SL g220975 (.A(sa21[3]),
    .B(n_8186),
    .Y(n_1542));
 XOR2xp5_ASAP7_75t_R g220976 (.A(n_3976),
    .B(n_8177),
    .Y(n_1341));
 OR2x2_ASAP7_75t_SL g220977 (.A(n_2919),
    .B(n_3298),
    .Y(n_1340));
 AOI21xp33_ASAP7_75t_R g220978 (.A1(n_1663),
    .A2(n_4345),
    .B(n_7660),
    .Y(n_1339));
 OR2x2_ASAP7_75t_SL g220979 (.A(sa31[7]),
    .B(sa31[1]),
    .Y(n_1338));
 XNOR2xp5_ASAP7_75t_SL g220981 (.A(n_936),
    .B(n_1141),
    .Y(n_26));
 OAI21xp33_ASAP7_75t_SL g221261 (.A1(sa11[2]),
    .A2(n_7124),
    .B(n_7182),
    .Y(n_8992));
 OAI21xp5_ASAP7_75t_SL g221262 (.A1(n_7163),
    .A2(n_6782),
    .B(sa22[5]),
    .Y(n_8993));
 O2A1O1Ixp33_ASAP7_75t_SL g221263 (.A1(n_5872),
    .A2(n_5750),
    .B(n_3360),
    .C(n_6787),
    .Y(n_8994));
 XNOR2xp5_ASAP7_75t_SL g221264 (.A(w3[27]),
    .B(n_8234),
    .Y(n_8995));
 XOR2xp5_ASAP7_75t_R g221265 (.A(w1[0]),
    .B(n_8261),
    .Y(n_8996));
 XOR2xp5_ASAP7_75t_L g221266 (.A(w1[7]),
    .B(n_8280),
    .Y(n_8997));
 XNOR2xp5_ASAP7_75t_L g221267 (.A(n_8234),
    .B(n_8656),
    .Y(n_8998));
 XOR2xp5_ASAP7_75t_SL g221268 (.A(w2[17]),
    .B(n_8343),
    .Y(n_8999));
 XOR2xp5_ASAP7_75t_SL g221269 (.A(n_8299),
    .B(n_8311),
    .Y(n_9000));
 XOR2x2_ASAP7_75t_SL g221270 (.A(n_207),
    .B(n_8253),
    .Y(n_9001));
 OR2x2_ASAP7_75t_SL g222998 (.A(n_8625),
    .B(u0_n_31924),
    .Y(n_11516));
 A2O1A1Ixp33_ASAP7_75t_L g222999 (.A1(n_1547),
    .A2(n_5414),
    .B(n_5778),
    .C(n_3509),
    .Y(n_11517));
 FAx1_ASAP7_75t_SL g223000 (.SN(n_11518),
    .A(n_724),
    .B(n_729),
    .CI(n_725),
    .CON(UNCONNECTED));
 HAxp5_ASAP7_75t_R g223002 (.A(u0_r0_rcnt[1]),
    .B(u0_r0_rcnt[0]),
    .CON(n_11521),
    .SN(n_11520));
 OAI21xp33_ASAP7_75t_SL g223780 (.A1(sa20[3]),
    .A2(n_2182),
    .B(n_7842),
    .Y(n_12816));
 INVx5_ASAP7_75t_SL g95636 (.A(sa33[1]),
    .Y(n_8204));
 INVx2_ASAP7_75t_SL g95637 (.A(sa00[0]),
    .Y(n_8196));
 INVx5_ASAP7_75t_SL g95638 (.A(sa00[4]),
    .Y(n_8200));
 INVx4_ASAP7_75t_SL g95639 (.A(sa02[3]),
    .Y(n_8210));
 INVx5_ASAP7_75t_SL g95640 (.A(sa10[3]),
    .Y(n_8178));
 INVx2_ASAP7_75t_L g95641 (.A(sa11[5]),
    .Y(n_8209));
 INVx4_ASAP7_75t_SL g95643 (.A(sa13[0]),
    .Y(n_8188));
 INVx2_ASAP7_75t_SL g95644 (.A(sa20[2]),
    .Y(n_8179));
 INVx5_ASAP7_75t_SL g95645 (.A(sa20[1]),
    .Y(n_1862));
 INVx2_ASAP7_75t_SL g95646 (.A(sa21[5]),
    .Y(n_8183));
 INVx3_ASAP7_75t_SL g95647 (.A(sa22[0]),
    .Y(n_8217));
 INVx5_ASAP7_75t_SL g95648 (.A(sa31[3]),
    .Y(n_8181));
 INVx5_ASAP7_75t_SL g95649 (.A(sa30[3]),
    .Y(n_8177));
 INVx3_ASAP7_75t_SL g95650 (.A(sa13[1]),
    .Y(n_8192));
 INVx4_ASAP7_75t_SL g95651 (.A(sa13[6]),
    .Y(n_8211));
 INVx2_ASAP7_75t_SL g95652 (.A(sa13[5]),
    .Y(n_8207));
 INVx3_ASAP7_75t_L g95653 (.A(sa11[0]),
    .Y(n_8182));
 INVx5_ASAP7_75t_SL g95654 (.A(sa10[6]),
    .Y(n_8180));
 INVx2_ASAP7_75t_L g95655 (.A(sa03[5]),
    .Y(n_8197));
 INVx5_ASAP7_75t_SL g95656 (.A(sa02[4]),
    .Y(n_8212));
 INVx4_ASAP7_75t_SL g95657 (.A(sa00[7]),
    .Y(n_8206));
 INVx3_ASAP7_75t_SL g95658 (.A(sa31[0]),
    .Y(n_8213));
 INVx4_ASAP7_75t_SL g95659 (.A(sa30[1]),
    .Y(n_8187));
 INVx2_ASAP7_75t_SL g95660 (.A(sa21[6]),
    .Y(n_8186));
 INVx2_ASAP7_75t_SL g95661 (.A(sa13[3]),
    .Y(n_8195));
 INVx1_ASAP7_75t_SL g95662 (.A(sa03[0]),
    .Y(n_8215));
 INVx3_ASAP7_75t_SL g95663 (.A(sa02[2]),
    .Y(n_8208));
 INVx5_ASAP7_75t_SL g95664 (.A(sa13[4]),
    .Y(n_1959));
 INVx4_ASAP7_75t_SL g95665 (.A(sa11[1]),
    .Y(n_8184));
 INVx4_ASAP7_75t_SL g95666 (.A(sa00[1]),
    .Y(n_8198));
 INVx2_ASAP7_75t_SL g95668 (.A(sa32[0]),
    .Y(n_8203));
 INVx4_ASAP7_75t_SL g95669 (.A(sa30[7]),
    .Y(n_8205));
 INVx2_ASAP7_75t_R g95670 (.A(sa12[5]),
    .Y(n_8190));
 INVx2_ASAP7_75t_L g95671 (.A(sa32[6]),
    .Y(n_8214));
 INVx2_ASAP7_75t_SL g95672 (.A(sa12[2]),
    .Y(n_8199));
 INVx4_ASAP7_75t_SL g95673 (.A(sa33[4]),
    .Y(n_8189));
 INVx3_ASAP7_75t_R g95674 (.A(sa00[5]),
    .Y(n_8202));
 INVx4_ASAP7_75t_SL g95675 (.A(sa33[7]),
    .Y(n_8191));
 DFFHQNx1_ASAP7_75t_R ld_r_reg (.CLK(clk),
    .D(u0_n_32835),
    .QN(ld_r));
 SDFHx4_ASAP7_75t_SL \sa00_reg[0]  (.CLK(clk),
    .D(n_470),
    .QN(sa00[0]),
    .SE(n_107),
    .SI(n_1178));
 SDFHx4_ASAP7_75t_SL \sa00_reg[1]  (.CLK(clk),
    .D(n_462),
    .QN(sa00[1]),
    .SE(n_109),
    .SI(n_1199));
 DFFHQx4_ASAP7_75t_SL \sa00_reg[2]  (.CLK(clk),
    .D(n_1335),
    .Q(sa00[2]));
 SDFHx4_ASAP7_75t_SL \sa00_reg[3]  (.CLK(clk),
    .D(n_442),
    .QN(sa00[3]),
    .SE(n_104),
    .SI(n_1206));
 SDFHx4_ASAP7_75t_SL \sa00_reg[4]  (.CLK(clk),
    .D(n_487),
    .QN(sa00[4]),
    .SE(n_105),
    .SI(n_1207));
 DFFHQx4_ASAP7_75t_SL \sa00_reg[5]  (.CLK(clk),
    .D(n_1279),
    .Q(sa00[5]));
 SDFHx4_ASAP7_75t_SL \sa00_reg[6]  (.CLK(clk),
    .D(n_512),
    .QN(sa00[6]),
    .SE(n_108),
    .SI(n_1251));
 SDFHx4_ASAP7_75t_SL \sa00_reg[7]  (.CLK(clk),
    .D(n_520),
    .QN(sa00[7]),
    .SE(n_106),
    .SI(n_1249));
 SDFHx4_ASAP7_75t_SL \sa01_reg[0]  (.CLK(clk),
    .D(n_526),
    .QN(sa01[0]),
    .SE(n_105),
    .SI(n_1173));
 SDFHx4_ASAP7_75t_SL \sa01_reg[1]  (.CLK(clk),
    .D(n_534),
    .QN(sa01[1]),
    .SE(n_104),
    .SI(n_1284));
 SDFHx4_ASAP7_75t_SL \sa01_reg[2]  (.CLK(clk),
    .D(n_544),
    .QN(sa01[2]),
    .SE(n_104),
    .SI(n_1208));
 SDFHx4_ASAP7_75t_SL \sa01_reg[3]  (.CLK(clk),
    .D(n_550),
    .QN(sa01[3]),
    .SE(n_104),
    .SI(n_1303));
 SDFHx4_ASAP7_75t_SL \sa01_reg[4]  (.CLK(clk),
    .D(n_449),
    .QN(sa01[4]),
    .SE(n_112),
    .SI(n_1283));
 SDFHx4_ASAP7_75t_SL \sa01_reg[5]  (.CLK(clk),
    .D(n_493),
    .QN(sa01[5]),
    .SE(n_103),
    .SI(n_1210));
 SDFHx4_ASAP7_75t_SL \sa01_reg[6]  (.CLK(clk),
    .D(n_498),
    .QN(sa01[6]),
    .SE(n_104),
    .SI(n_1211));
 SDFHx4_ASAP7_75t_SL \sa01_reg[7]  (.CLK(clk),
    .D(n_500),
    .QN(sa01[7]),
    .SE(n_103),
    .SI(n_1196));
 SDFHx4_ASAP7_75t_L \sa02_reg[0]  (.CLK(clk),
    .D(n_467),
    .QN(sa02[0]),
    .SE(n_103),
    .SI(n_1182));
 SDFHx4_ASAP7_75t_SL \sa02_reg[1]  (.CLK(clk),
    .D(n_455),
    .QN(sa02[1]),
    .SE(n_102),
    .SI(n_1282));
 DFFHQx4_ASAP7_75t_SL \sa02_reg[2]  (.CLK(clk),
    .D(n_1332),
    .Q(sa02[2]));
 SDFHx4_ASAP7_75t_SL \sa02_reg[3]  (.CLK(clk),
    .D(n_468),
    .QN(sa02[3]),
    .SE(n_107),
    .SI(n_1194));
 SDFHx4_ASAP7_75t_SL \sa02_reg[4]  (.CLK(clk),
    .D(n_478),
    .QN(sa02[4]),
    .SE(n_109),
    .SI(n_1278));
 SDFHx2_ASAP7_75t_SL \sa02_reg[5]  (.CLK(clk),
    .D(n_473),
    .QN(sa02[5]),
    .SE(n_110),
    .SI(n_1195));
 SDFHx4_ASAP7_75t_SL \sa02_reg[6]  (.CLK(clk),
    .D(n_469),
    .QN(sa02[6]),
    .SE(n_107),
    .SI(n_1190));
 SDFHx4_ASAP7_75t_SL \sa02_reg[7]  (.CLK(clk),
    .D(n_464),
    .QN(sa02[7]),
    .SE(n_106),
    .SI(n_1267));
 DFFHQx4_ASAP7_75t_SL \sa03_reg[0]  (.CLK(clk),
    .D(n_1331),
    .Q(sa03[0]));
 SDFHx4_ASAP7_75t_SL \sa03_reg[1]  (.CLK(clk),
    .D(n_454),
    .QN(sa03[1]),
    .SE(n_102),
    .SI(n_1200));
 SDFHx1_ASAP7_75t_SL \sa03_reg[2]  (.CLK(clk),
    .QN(sa03[2]),
    .D(n_448),
    .SE(n_103),
    .SI(n_1201));
 SDFHx4_ASAP7_75t_SL \sa03_reg[3]  (.CLK(clk),
    .D(n_444),
    .QN(sa03[3]),
    .SE(n_108),
    .SI(n_1323));
 SDFHx4_ASAP7_75t_SL \sa03_reg[4]  (.CLK(clk),
    .D(n_440),
    .QN(sa03[4]),
    .SE(n_105),
    .SI(n_1286));
 SDFHx1_ASAP7_75t_L \sa03_reg[5]  (.CLK(clk),
    .QN(sa03[5]),
    .D(n_484),
    .SE(n_110),
    .SI(n_16));
 SDFHx1_ASAP7_75t_SL \sa03_reg[6]  (.CLK(clk),
    .QN(sa03[6]),
    .D(n_489),
    .SE(n_109),
    .SI(n_1260));
 SDFHx4_ASAP7_75t_SL \sa03_reg[7]  (.CLK(clk),
    .D(n_495),
    .QN(sa03[7]),
    .SE(n_110),
    .SI(n_1319));
 SDFHx1_ASAP7_75t_SL \sa10_reg[0]  (.CLK(clk),
    .QN(sa10[0]),
    .D(n_504),
    .SE(n_106),
    .SI(n_1257));
 SDFHx4_ASAP7_75t_SL \sa10_reg[1]  (.CLK(clk),
    .D(n_510),
    .QN(sa10[1]),
    .SE(n_104),
    .SI(n_1288));
 SDFHx4_ASAP7_75t_SL \sa10_reg[2]  (.CLK(clk),
    .D(n_2774),
    .QN(sa10[2]),
    .SE(n_2654),
    .SI(n_7613));
 SDFHx4_ASAP7_75t_SL \sa10_reg[3]  (.CLK(clk),
    .D(n_511),
    .QN(sa10[3]),
    .SE(n_102),
    .SI(n_1316));
 SDFHx4_ASAP7_75t_SL \sa10_reg[4]  (.CLK(clk),
    .D(n_516),
    .QN(sa10[4]),
    .SE(n_104),
    .SI(n_1314));
 DFFHQx4_ASAP7_75t_L \sa10_reg[5]  (.CLK(clk),
    .D(n_1329),
    .Q(sa10[5]));
 SDFHx4_ASAP7_75t_SL \sa10_reg[6]  (.CLK(clk),
    .D(n_524),
    .QN(sa10[6]),
    .SE(n_102),
    .SI(n_1248));
 SDFHx4_ASAP7_75t_SL \sa10_reg[7]  (.CLK(clk),
    .D(n_528),
    .QN(sa10[7]),
    .SE(n_106),
    .SI(n_1246));
 SDFHx4_ASAP7_75t_SL \sa11_reg[0]  (.CLK(clk),
    .D(n_1187),
    .QN(sa11[0]),
    .SE(n_40),
    .SI(n_532));
 SDFHx4_ASAP7_75t_SL \sa11_reg[1]  (.CLK(clk),
    .D(n_536),
    .QN(sa11[1]),
    .SE(n_103),
    .SI(n_1309));
 SDFHx4_ASAP7_75t_SL \sa11_reg[2]  (.CLK(clk),
    .D(n_488),
    .QN(sa11[2]),
    .SE(n_106),
    .SI(n_1186));
 SDFHx4_ASAP7_75t_SL \sa11_reg[3]  (.CLK(clk),
    .D(n_542),
    .QN(sa11[3]),
    .SE(n_110),
    .SI(n_1304));
 SDFHx4_ASAP7_75t_SL \sa11_reg[4]  (.CLK(clk),
    .D(n_545),
    .QN(sa11[4]),
    .SE(n_103),
    .SI(n_1276));
 SDFHx1_ASAP7_75t_L \sa11_reg[5]  (.CLK(clk),
    .QN(sa11[5]),
    .D(n_552),
    .SE(n_108),
    .SI(n_1209));
 SDFHx4_ASAP7_75t_SL \sa11_reg[6]  (.CLK(clk),
    .D(n_1205),
    .QN(sa11[6]),
    .SE(n_40),
    .SI(n_558));
 SDFHx4_ASAP7_75t_SL \sa11_reg[7]  (.CLK(clk),
    .D(n_560),
    .QN(sa11[7]),
    .SE(n_109),
    .SI(n_1203));
 SDFHx4_ASAP7_75t_SL \sa12_reg[0]  (.CLK(clk),
    .D(n_1183),
    .QN(sa12[0]),
    .SE(n_41),
    .SI(n_563));
 SDFHx4_ASAP7_75t_SL \sa12_reg[1]  (.CLK(clk),
    .D(n_518),
    .QN(sa12[1]),
    .SE(n_107),
    .SI(n_1281));
 SDFHx4_ASAP7_75t_SL \sa12_reg[2]  (.CLK(clk),
    .D(n_499),
    .QN(sa12[2]),
    .SE(n_109),
    .SI(n_1185));
 SDFHx1_ASAP7_75t_SL \sa12_reg[3]  (.CLK(clk),
    .QN(sa12[3]),
    .D(n_494),
    .SE(n_105),
    .SI(n_1299));
 SDFHx4_ASAP7_75t_SL \sa12_reg[4]  (.CLK(clk),
    .D(n_496),
    .QN(sa12[4]),
    .SE(n_107),
    .SI(n_1280));
 SDFHx1_ASAP7_75t_SL \sa12_reg[5]  (.CLK(clk),
    .QN(sa12[5]),
    .D(n_513),
    .SE(n_105),
    .SI(n_1197));
 SDFHx4_ASAP7_75t_L \sa12_reg[6]  (.CLK(clk),
    .D(n_459),
    .QN(sa12[6]),
    .SE(n_112),
    .SI(n_1177));
 SDFHx4_ASAP7_75t_SL \sa12_reg[7]  (.CLK(clk),
    .D(n_501),
    .QN(sa12[7]),
    .SE(n_105),
    .SI(n_1179));
 SDFHx4_ASAP7_75t_L \sa13_reg[0]  (.CLK(clk),
    .D(n_1188),
    .QN(sa13[0]),
    .SE(n_41),
    .SI(n_457));
 SDFHx4_ASAP7_75t_SL \sa13_reg[1]  (.CLK(clk),
    .D(n_507),
    .QN(sa13[1]),
    .SE(n_106),
    .SI(n_1298));
 SDFHx1_ASAP7_75t_SL \sa13_reg[2]  (.CLK(clk),
    .QN(sa13[2]),
    .D(n_1184),
    .SE(n_40),
    .SI(n_551));
 SDFHx4_ASAP7_75t_SL \sa13_reg[3]  (.CLK(clk),
    .D(n_553),
    .QN(sa13[3]),
    .SE(n_102),
    .SI(n_1297));
 SDFHx4_ASAP7_75t_SL \sa13_reg[4]  (.CLK(clk),
    .D(n_555),
    .QN(sa13[4]),
    .SE(n_109),
    .SI(n_1296));
 SDFHx1_ASAP7_75t_L \sa13_reg[5]  (.CLK(clk),
    .QN(sa13[5]),
    .D(n_557),
    .SE(n_102),
    .SI(n_11518));
 SDFHx4_ASAP7_75t_SL \sa13_reg[6]  (.CLK(clk),
    .D(n_561),
    .QN(sa13[6]),
    .SE(n_107),
    .SI(n_1212));
 SDFHx4_ASAP7_75t_SL \sa13_reg[7]  (.CLK(clk),
    .D(n_480),
    .QN(sa13[7]),
    .SE(n_109),
    .SI(n_1189));
 SDFHx4_ASAP7_75t_SL \sa20_reg[0]  (.CLK(clk),
    .D(n_479),
    .QN(sa20[0]),
    .SE(n_109),
    .SI(n_1270));
 SDFHx4_ASAP7_75t_SL \sa20_reg[1]  (.CLK(clk),
    .D(n_477),
    .QN(sa20[1]),
    .SE(n_102),
    .SI(n_1294));
 SDFHx1_ASAP7_75t_SL \sa20_reg[2]  (.CLK(clk),
    .QN(sa20[2]),
    .D(n_476),
    .SE(n_111),
    .SI(n_1328));
 SDFHx4_ASAP7_75t_SL \sa20_reg[3]  (.CLK(clk),
    .D(n_474),
    .QN(sa20[3]),
    .SE(n_102),
    .SI(n_1327));
 SDFHx4_ASAP7_75t_SL \sa20_reg[4]  (.CLK(clk),
    .D(n_472),
    .QN(sa20[4]),
    .SE(n_103),
    .SI(n_1293));
 SDFHx1_ASAP7_75t_SL \sa20_reg[5]  (.CLK(clk),
    .QN(sa20[5]),
    .D(n_471),
    .SE(n_111),
    .SI(n_1269));
 SDFHx1_ASAP7_75t_SL \sa20_reg[6]  (.CLK(clk),
    .QN(sa20[6]),
    .D(n_2775),
    .SE(n_2654),
    .SI(n_7614));
 SDFHx4_ASAP7_75t_SL \sa20_reg[7]  (.CLK(clk),
    .D(n_564),
    .QN(sa20[7]),
    .SE(n_104),
    .SI(n_1213));
 SDFHx4_ASAP7_75t_SL \sa21_reg[0]  (.CLK(clk),
    .D(n_1268),
    .QN(sa21[0]),
    .SE(n_41),
    .SI(n_466));
 SDFHx4_ASAP7_75t_SL \sa21_reg[1]  (.CLK(clk),
    .D(n_463),
    .QN(sa21[1]),
    .SE(n_109),
    .SI(n_1198));
 SDFHx4_ASAP7_75t_SL \sa21_reg[2]  (.CLK(clk),
    .D(n_461),
    .QN(sa21[2]),
    .SE(n_103),
    .SI(n_1326));
 SDFHx4_ASAP7_75t_SL \sa21_reg[3]  (.CLK(clk),
    .D(n_460),
    .QN(sa21[3]),
    .SE(n_102),
    .SI(n_19));
 SDFHx4_ASAP7_75t_SL \sa21_reg[4]  (.CLK(clk),
    .D(n_456),
    .QN(sa21[4]),
    .SE(n_103),
    .SI(n_1324));
 SDFHx2_ASAP7_75t_SL \sa21_reg[5]  (.CLK(clk),
    .D(n_453),
    .QN(sa21[5]),
    .SE(n_105),
    .SI(n_1266));
 SDFHx4_ASAP7_75t_SL \sa21_reg[6]  (.CLK(clk),
    .D(n_452),
    .QN(sa21[6]),
    .SE(n_106),
    .SI(n_1265));
 SDFHx4_ASAP7_75t_SL \sa21_reg[7]  (.CLK(clk),
    .D(n_450),
    .QN(sa21[7]),
    .SE(n_108),
    .SI(n_1264));
 SDFHx4_ASAP7_75t_SL \sa22_reg[0]  (.CLK(clk),
    .D(n_447),
    .QN(sa22[0]),
    .SE(n_103),
    .SI(n_1263));
 SDFHx4_ASAP7_75t_SL \sa22_reg[1]  (.CLK(clk),
    .D(n_446),
    .QN(sa22[1]),
    .SE(n_109),
    .SI(n_1292));
 SDFHx4_ASAP7_75t_SL \sa22_reg[2]  (.CLK(clk),
    .D(n_445),
    .QN(sa22[2]),
    .SE(n_102),
    .SI(n_1322));
 SDFHx4_ASAP7_75t_SL \sa22_reg[3]  (.CLK(clk),
    .D(n_443),
    .QN(sa22[3]),
    .SE(n_106),
    .SI(n_1321));
 SDFHx4_ASAP7_75t_SL \sa22_reg[4]  (.CLK(clk),
    .D(n_441),
    .QN(sa22[4]),
    .SE(n_107),
    .SI(n_1291));
 SDFHx2_ASAP7_75t_SL \sa22_reg[5]  (.CLK(clk),
    .D(n_481),
    .QN(sa22[5]),
    .SE(n_105),
    .SI(n_1262));
 SDFHx4_ASAP7_75t_SL \sa22_reg[6]  (.CLK(clk),
    .D(n_482),
    .QN(sa22[6]),
    .SE(n_104),
    .SI(n_1261));
 SDFHx4_ASAP7_75t_SL \sa22_reg[7]  (.CLK(clk),
    .D(n_483),
    .QN(sa22[7]),
    .SE(n_111),
    .SI(n_1320));
 SDFHx4_ASAP7_75t_L \sa23_reg[0]  (.CLK(clk),
    .D(n_485),
    .QN(sa23[0]),
    .SE(n_105),
    .SI(n_1176));
 SDFHx4_ASAP7_75t_SL \sa23_reg[1]  (.CLK(clk),
    .D(n_486),
    .QN(sa23[1]),
    .SE(n_109),
    .SI(n_1290));
 SDFHx1_ASAP7_75t_L \sa23_reg[2]  (.CLK(clk),
    .QN(sa23[2]),
    .D(n_490),
    .SE(n_110),
    .SI(n_1259));
 SDFHx4_ASAP7_75t_SL \sa23_reg[3]  (.CLK(clk),
    .D(n_491),
    .QN(sa23[3]),
    .SE(n_105),
    .SI(n_1277));
 SDFHx4_ASAP7_75t_SL \sa23_reg[4]  (.CLK(clk),
    .D(n_497),
    .QN(sa23[4]),
    .SE(n_104),
    .SI(n_1289));
 SDFHx2_ASAP7_75t_SL \sa23_reg[5]  (.CLK(clk),
    .D(n_502),
    .QN(sa23[5]),
    .SE(n_107),
    .SI(n_1258));
 SDFHx1_ASAP7_75t_SL \sa23_reg[6]  (.CLK(clk),
    .QN(sa23[6]),
    .D(n_2776),
    .SE(n_2654),
    .SI(n_7945));
 SDFHx4_ASAP7_75t_SL \sa23_reg[7]  (.CLK(clk),
    .D(n_505),
    .QN(sa23[7]),
    .SE(n_103),
    .SI(n_1193));
 SDFHx4_ASAP7_75t_SL \sa30_reg[0]  (.CLK(clk),
    .D(n_506),
    .QN(sa30[0]),
    .SE(n_107),
    .SI(n_1256));
 SDFHx4_ASAP7_75t_SL \sa30_reg[1]  (.CLK(clk),
    .D(n_508),
    .QN(sa30[1]),
    .SE(n_106),
    .SI(n_1318));
 SDFHx4_ASAP7_75t_SL \sa30_reg[2]  (.CLK(clk),
    .D(n_492),
    .QN(sa30[2]),
    .SE(n_106),
    .SI(n_1255));
 SDFHx4_ASAP7_75t_SL \sa30_reg[3]  (.CLK(clk),
    .D(n_475),
    .QN(sa30[3]),
    .SE(n_108),
    .SI(n_1317));
 SDFHx4_ASAP7_75t_SL \sa30_reg[4]  (.CLK(clk),
    .D(n_514),
    .QN(sa30[4]),
    .SE(n_110),
    .SI(n_1315));
 SDFHx1_ASAP7_75t_SL \sa30_reg[5]  (.CLK(clk),
    .QN(sa30[5]),
    .D(n_515),
    .SE(n_110),
    .SI(n_1254));
 SDFHx4_ASAP7_75t_SL \sa30_reg[6]  (.CLK(clk),
    .D(n_517),
    .QN(sa30[6]),
    .SE(n_108),
    .SI(n_1253));
 SDFHx4_ASAP7_75t_SL \sa30_reg[7]  (.CLK(clk),
    .D(n_519),
    .QN(sa30[7]),
    .SE(n_110),
    .SI(n_1252));
 SDFHx1_ASAP7_75t_SL \sa31_reg[0]  (.CLK(clk),
    .QN(sa31[0]),
    .D(n_521),
    .SE(n_107),
    .SI(n_1174));
 SDFHx4_ASAP7_75t_SL \sa31_reg[1]  (.CLK(clk),
    .D(n_522),
    .QN(sa31[1]),
    .SE(n_107),
    .SI(n_1285));
 DFFHQNx1_ASAP7_75t_L \sa31_reg[2]  (.CLK(clk),
    .D(n_1334),
    .QN(sa31[2]));
 SDFHx4_ASAP7_75t_SL \sa31_reg[3]  (.CLK(clk),
    .D(n_525),
    .QN(sa31[3]),
    .SE(n_107),
    .SI(n_1312));
 SDFHx4_ASAP7_75t_SL \sa31_reg[4]  (.CLK(clk),
    .D(n_509),
    .QN(sa31[4]),
    .SE(n_109),
    .SI(n_1311));
 SDFHx1_ASAP7_75t_SL \sa31_reg[5]  (.CLK(clk),
    .QN(sa31[5]),
    .D(n_527),
    .SE(n_104),
    .SI(n_1247));
 SDFHx4_ASAP7_75t_SL \sa31_reg[6]  (.CLK(clk),
    .D(n_1273),
    .QN(sa31[6]),
    .SE(n_41),
    .SI(n_530));
 SDFHx4_ASAP7_75t_SL \sa31_reg[7]  (.CLK(clk),
    .D(n_531),
    .QN(sa31[7]),
    .SE(n_108),
    .SI(n_1180));
 SDFHx1_ASAP7_75t_SL \sa32_reg[0]  (.CLK(clk),
    .QN(sa32[0]),
    .D(n_539),
    .SE(n_102),
    .SI(n_1172));
 SDFHx4_ASAP7_75t_SL \sa32_reg[1]  (.CLK(clk),
    .D(n_535),
    .QN(sa32[1]),
    .SE(n_102),
    .SI(n_1310));
 SDFHx4_ASAP7_75t_SL \sa32_reg[2]  (.CLK(clk),
    .D(n_537),
    .QN(sa32[2]),
    .SE(n_105),
    .SI(n_1308));
 SDFHx1_ASAP7_75t_SL \sa32_reg[3]  (.CLK(clk),
    .QN(sa32[3]),
    .D(n_538),
    .SE(n_104),
    .SI(n_1307));
 SDFHx4_ASAP7_75t_SL \sa32_reg[4]  (.CLK(clk),
    .D(n_540),
    .QN(sa32[4]),
    .SE(n_108),
    .SI(n_1306));
 DFFHQx4_ASAP7_75t_SL \sa32_reg[5]  (.CLK(clk),
    .D(n_1333),
    .Q(sa32[5]));
 SDFHx4_ASAP7_75t_SL \sa32_reg[6]  (.CLK(clk),
    .D(n_543),
    .QN(sa32[6]),
    .SE(n_106),
    .SI(n_1171));
 SDFHx4_ASAP7_75t_SL \sa32_reg[7]  (.CLK(clk),
    .D(n_546),
    .QN(sa32[7]),
    .SE(n_108),
    .SI(n_1181));
 SDFHx4_ASAP7_75t_SL \sa33_reg[0]  (.CLK(clk),
    .D(n_547),
    .QN(sa33[0]),
    .SE(n_105),
    .SI(n_1170));
 SDFHx4_ASAP7_75t_SL \sa33_reg[1]  (.CLK(clk),
    .D(n_548),
    .QN(sa33[1]),
    .SE(n_108),
    .SI(n_1302));
 DFFHQx4_ASAP7_75t_SL \sa33_reg[2]  (.CLK(clk),
    .D(n_1330),
    .Q(sa33[2]));
 SDFHx4_ASAP7_75t_SL \sa33_reg[3]  (.CLK(clk),
    .D(n_554),
    .QN(sa33[3]),
    .SE(n_108),
    .SI(n_1301));
 SDFHx4_ASAP7_75t_SL \sa33_reg[4]  (.CLK(clk),
    .D(n_529),
    .QN(sa33[4]),
    .SE(n_103),
    .SI(n_1300));
 SDFHx2_ASAP7_75t_SL \sa33_reg[5]  (.CLK(clk),
    .D(n_559),
    .QN(sa33[5]),
    .SE(n_108),
    .SI(n_1204));
 SDFHx4_ASAP7_75t_SL \sa33_reg[6]  (.CLK(clk),
    .D(n_1192),
    .QN(sa33[6]),
    .SE(n_40),
    .SI(n_465));
 SDFHx4_ASAP7_75t_SL \sa33_reg[7]  (.CLK(clk),
    .D(n_562),
    .QN(sa33[7]),
    .SE(n_106),
    .SI(n_1202));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[0]  (.CLK(clk),
    .D(n_872),
    .QN(text_in_r[0]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[100]  (.CLK(clk),
    .D(n_783),
    .QN(text_in_r[100]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[101]  (.CLK(clk),
    .D(n_782),
    .QN(text_in_r[101]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[102]  (.CLK(clk),
    .D(n_781),
    .QN(text_in_r[102]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[103]  (.CLK(clk),
    .D(n_780),
    .QN(text_in_r[103]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[104]  (.CLK(clk),
    .D(n_779),
    .QN(text_in_r[104]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[105]  (.CLK(clk),
    .D(n_778),
    .QN(text_in_r[105]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[106]  (.CLK(clk),
    .D(n_777),
    .QN(text_in_r[106]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[107]  (.CLK(clk),
    .D(n_776),
    .QN(text_in_r[107]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[108]  (.CLK(clk),
    .D(n_775),
    .QN(text_in_r[108]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[109]  (.CLK(clk),
    .D(n_774),
    .QN(text_in_r[109]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[10]  (.CLK(clk),
    .D(n_863),
    .QN(text_in_r[10]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[110]  (.CLK(clk),
    .D(n_773),
    .QN(text_in_r[110]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[111]  (.CLK(clk),
    .D(n_772),
    .QN(text_in_r[111]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[112]  (.CLK(clk),
    .D(n_771),
    .QN(text_in_r[112]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[113]  (.CLK(clk),
    .D(n_770),
    .QN(text_in_r[113]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[114]  (.CLK(clk),
    .D(n_769),
    .QN(text_in_r[114]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[115]  (.CLK(clk),
    .D(n_768),
    .QN(text_in_r[115]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[116]  (.CLK(clk),
    .D(n_846),
    .QN(text_in_r[116]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[117]  (.CLK(clk),
    .D(n_767),
    .QN(text_in_r[117]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[118]  (.CLK(clk),
    .D(n_766),
    .QN(text_in_r[118]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[119]  (.CLK(clk),
    .D(n_765),
    .QN(text_in_r[119]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[11]  (.CLK(clk),
    .D(n_862),
    .QN(text_in_r[11]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[120]  (.CLK(clk),
    .D(n_760),
    .QN(text_in_r[120]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[121]  (.CLK(clk),
    .D(n_764),
    .QN(text_in_r[121]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[122]  (.CLK(clk),
    .D(n_873),
    .QN(text_in_r[122]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[123]  (.CLK(clk),
    .D(n_763),
    .QN(text_in_r[123]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[124]  (.CLK(clk),
    .D(n_762),
    .QN(text_in_r[124]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[125]  (.CLK(clk),
    .D(n_761),
    .QN(text_in_r[125]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[126]  (.CLK(clk),
    .D(n_884),
    .QN(text_in_r[126]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[127]  (.CLK(clk),
    .D(n_888),
    .QN(text_in_r[127]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[12]  (.CLK(clk),
    .D(n_861),
    .QN(text_in_r[12]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[13]  (.CLK(clk),
    .D(n_860),
    .QN(text_in_r[13]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[14]  (.CLK(clk),
    .D(n_859),
    .QN(text_in_r[14]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[15]  (.CLK(clk),
    .D(n_858),
    .QN(text_in_r[15]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[16]  (.CLK(clk),
    .D(n_857),
    .QN(text_in_r[16]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[17]  (.CLK(clk),
    .D(n_856),
    .QN(text_in_r[17]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[18]  (.CLK(clk),
    .D(n_855),
    .QN(text_in_r[18]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[19]  (.CLK(clk),
    .D(n_854),
    .QN(text_in_r[19]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[1]  (.CLK(clk),
    .D(n_871),
    .QN(text_in_r[1]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[20]  (.CLK(clk),
    .D(n_853),
    .QN(text_in_r[20]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[21]  (.CLK(clk),
    .D(n_852),
    .QN(text_in_r[21]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[22]  (.CLK(clk),
    .D(n_851),
    .QN(text_in_r[22]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[23]  (.CLK(clk),
    .D(n_850),
    .QN(text_in_r[23]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[24]  (.CLK(clk),
    .D(n_875),
    .QN(text_in_r[24]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[25]  (.CLK(clk),
    .D(n_849),
    .QN(text_in_r[25]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[26]  (.CLK(clk),
    .D(n_848),
    .QN(text_in_r[26]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[27]  (.CLK(clk),
    .D(n_847),
    .QN(text_in_r[27]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[28]  (.CLK(clk),
    .D(n_878),
    .QN(text_in_r[28]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[29]  (.CLK(clk),
    .D(n_882),
    .QN(text_in_r[29]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[2]  (.CLK(clk),
    .D(n_885),
    .QN(text_in_r[2]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[30]  (.CLK(clk),
    .D(n_845),
    .QN(text_in_r[30]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[31]  (.CLK(clk),
    .D(n_844),
    .QN(text_in_r[31]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[32]  (.CLK(clk),
    .D(n_843),
    .QN(text_in_r[32]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[33]  (.CLK(clk),
    .D(n_842),
    .QN(text_in_r[33]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[34]  (.CLK(clk),
    .D(n_841),
    .QN(text_in_r[34]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[35]  (.CLK(clk),
    .D(n_840),
    .QN(text_in_r[35]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[36]  (.CLK(clk),
    .D(n_839),
    .QN(text_in_r[36]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[37]  (.CLK(clk),
    .D(n_838),
    .QN(text_in_r[37]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[38]  (.CLK(clk),
    .D(n_886),
    .QN(text_in_r[38]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[39]  (.CLK(clk),
    .D(n_837),
    .QN(text_in_r[39]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[3]  (.CLK(clk),
    .D(n_870),
    .QN(text_in_r[3]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[40]  (.CLK(clk),
    .D(n_836),
    .QN(text_in_r[40]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[41]  (.CLK(clk),
    .D(n_835),
    .QN(text_in_r[41]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[42]  (.CLK(clk),
    .D(n_865),
    .QN(text_in_r[42]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[43]  (.CLK(clk),
    .D(n_834),
    .QN(text_in_r[43]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[44]  (.CLK(clk),
    .D(n_792),
    .QN(text_in_r[44]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[45]  (.CLK(clk),
    .D(n_833),
    .QN(text_in_r[45]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[46]  (.CLK(clk),
    .D(n_832),
    .QN(text_in_r[46]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[47]  (.CLK(clk),
    .D(n_831),
    .QN(text_in_r[47]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[48]  (.CLK(clk),
    .D(n_830),
    .QN(text_in_r[48]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[49]  (.CLK(clk),
    .D(n_829),
    .QN(text_in_r[49]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[4]  (.CLK(clk),
    .D(n_869),
    .QN(text_in_r[4]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[50]  (.CLK(clk),
    .D(n_828),
    .QN(text_in_r[50]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[51]  (.CLK(clk),
    .D(n_827),
    .QN(text_in_r[51]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[52]  (.CLK(clk),
    .D(n_826),
    .QN(text_in_r[52]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[53]  (.CLK(clk),
    .D(n_825),
    .QN(text_in_r[53]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[54]  (.CLK(clk),
    .D(n_824),
    .QN(text_in_r[54]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[55]  (.CLK(clk),
    .D(n_823),
    .QN(text_in_r[55]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[56]  (.CLK(clk),
    .D(n_822),
    .QN(text_in_r[56]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[57]  (.CLK(clk),
    .D(n_821),
    .QN(text_in_r[57]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[58]  (.CLK(clk),
    .D(n_820),
    .QN(text_in_r[58]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[59]  (.CLK(clk),
    .D(n_819),
    .QN(text_in_r[59]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[5]  (.CLK(clk),
    .D(n_868),
    .QN(text_in_r[5]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[60]  (.CLK(clk),
    .D(n_883),
    .QN(text_in_r[60]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[61]  (.CLK(clk),
    .D(n_818),
    .QN(text_in_r[61]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[62]  (.CLK(clk),
    .D(n_817),
    .QN(text_in_r[62]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[63]  (.CLK(clk),
    .D(n_816),
    .QN(text_in_r[63]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[64]  (.CLK(clk),
    .D(n_815),
    .QN(text_in_r[64]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[65]  (.CLK(clk),
    .D(n_877),
    .QN(text_in_r[65]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[66]  (.CLK(clk),
    .D(n_814),
    .QN(text_in_r[66]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[67]  (.CLK(clk),
    .D(n_813),
    .QN(text_in_r[67]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[68]  (.CLK(clk),
    .D(n_812),
    .QN(text_in_r[68]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[69]  (.CLK(clk),
    .D(n_811),
    .QN(text_in_r[69]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[6]  (.CLK(clk),
    .D(n_874),
    .QN(text_in_r[6]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[70]  (.CLK(clk),
    .D(n_810),
    .QN(text_in_r[70]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[71]  (.CLK(clk),
    .D(n_809),
    .QN(text_in_r[71]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[72]  (.CLK(clk),
    .D(n_808),
    .QN(text_in_r[72]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[73]  (.CLK(clk),
    .D(n_807),
    .QN(text_in_r[73]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[74]  (.CLK(clk),
    .D(n_806),
    .QN(text_in_r[74]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[75]  (.CLK(clk),
    .D(n_805),
    .QN(text_in_r[75]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[76]  (.CLK(clk),
    .D(n_881),
    .QN(text_in_r[76]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[77]  (.CLK(clk),
    .D(n_804),
    .QN(text_in_r[77]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[78]  (.CLK(clk),
    .D(n_803),
    .QN(text_in_r[78]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[79]  (.CLK(clk),
    .D(n_802),
    .QN(text_in_r[79]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[7]  (.CLK(clk),
    .D(n_867),
    .QN(text_in_r[7]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[80]  (.CLK(clk),
    .D(n_879),
    .QN(text_in_r[80]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[81]  (.CLK(clk),
    .D(n_801),
    .QN(text_in_r[81]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[82]  (.CLK(clk),
    .D(n_800),
    .QN(text_in_r[82]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[83]  (.CLK(clk),
    .D(n_799),
    .QN(text_in_r[83]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[84]  (.CLK(clk),
    .D(n_798),
    .QN(text_in_r[84]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[85]  (.CLK(clk),
    .D(n_797),
    .QN(text_in_r[85]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[86]  (.CLK(clk),
    .D(n_796),
    .QN(text_in_r[86]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[87]  (.CLK(clk),
    .D(n_795),
    .QN(text_in_r[87]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[88]  (.CLK(clk),
    .D(n_876),
    .QN(text_in_r[88]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[89]  (.CLK(clk),
    .D(n_794),
    .QN(text_in_r[89]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[8]  (.CLK(clk),
    .D(n_866),
    .QN(text_in_r[8]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[90]  (.CLK(clk),
    .D(n_793),
    .QN(text_in_r[90]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[91]  (.CLK(clk),
    .D(n_791),
    .QN(text_in_r[91]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[92]  (.CLK(clk),
    .D(n_790),
    .QN(text_in_r[92]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[93]  (.CLK(clk),
    .D(n_789),
    .QN(text_in_r[93]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[94]  (.CLK(clk),
    .D(n_788),
    .QN(text_in_r[94]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[95]  (.CLK(clk),
    .D(n_787),
    .QN(text_in_r[95]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[96]  (.CLK(clk),
    .D(n_786),
    .QN(text_in_r[96]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[97]  (.CLK(clk),
    .D(n_785),
    .QN(text_in_r[97]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[98]  (.CLK(clk),
    .D(n_880),
    .QN(text_in_r[98]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[99]  (.CLK(clk),
    .D(n_784),
    .QN(text_in_r[99]));
 DFFHQNx1_ASAP7_75t_R \text_in_r_reg[9]  (.CLK(clk),
    .D(n_864),
    .QN(text_in_r[9]));
 SDFHx1_ASAP7_75t_R \text_out_reg[0]  (.CLK(clk),
    .QN(\text_out[0]_3160 ),
    .D(n_7518),
    .SE(w3[0]),
    .SI(n_7519));
 SDFHx1_ASAP7_75t_R \text_out_reg[100]  (.CLK(clk),
    .QN(\text_out[100]_3140 ),
    .D(n_8923),
    .SE(w0[4]),
    .SI(n_8922));
 SDFHx1_ASAP7_75t_R \text_out_reg[101]  (.CLK(clk),
    .QN(\text_out[101]_3141 ),
    .D(n_8260),
    .SE(w0[5]),
    .SI(n_148));
 SDFHx1_ASAP7_75t_R \text_out_reg[102]  (.CLK(clk),
    .QN(\text_out[102]_3142 ),
    .D(n_8279),
    .SE(w0[6]),
    .SI(n_194));
 SDFHx1_ASAP7_75t_R \text_out_reg[103]  (.CLK(clk),
    .QN(\text_out[103]_3143 ),
    .D(n_8259),
    .SE(w0[7]),
    .SI(n_119));
 SDFHx1_ASAP7_75t_R \text_out_reg[104]  (.CLK(clk),
    .QN(\text_out[104]_3104 ),
    .D(n_7564),
    .SE(w0[8]),
    .SI(n_7565));
 SDFHx1_ASAP7_75t_R \text_out_reg[105]  (.CLK(clk),
    .QN(\text_out[105]_3105 ),
    .D(n_203),
    .SE(w0[9]),
    .SI(n_8325));
 SDFHx1_ASAP7_75t_R \text_out_reg[106]  (.CLK(clk),
    .QN(\text_out[106]_3106 ),
    .D(n_324),
    .SE(w0[10]),
    .SI(n_62));
 SDFHx1_ASAP7_75t_R \text_out_reg[107]  (.CLK(clk),
    .QN(\text_out[107]_3107 ),
    .D(n_7554),
    .SE(w0[11]),
    .SI(n_7555));
 SDFHx1_ASAP7_75t_R \text_out_reg[108]  (.CLK(clk),
    .QN(\text_out[108]_3108 ),
    .D(n_150),
    .SE(w0[12]),
    .SI(n_8323));
 SDFHx1_ASAP7_75t_R \text_out_reg[109]  (.CLK(clk),
    .QN(\text_out[109]_3109 ),
    .D(n_8252),
    .SE(w0[13]),
    .SI(n_361));
 SDFHx1_ASAP7_75t_R \text_out_reg[10]  (.CLK(clk),
    .QN(\text_out[10]_3130 ),
    .D(n_68),
    .SE(w3[10]),
    .SI(n_8333));
 SDFHx1_ASAP7_75t_R \text_out_reg[110]  (.CLK(clk),
    .QN(\text_out[110]_3110 ),
    .D(w0[14]),
    .SE(n_8275),
    .SI(n_2035));
 SDFHx1_ASAP7_75t_R \text_out_reg[111]  (.CLK(clk),
    .QN(\text_out[111]_3111 ),
    .D(n_7537),
    .SE(w0[15]),
    .SI(n_332));
 SDFHx1_ASAP7_75t_R \text_out_reg[112]  (.CLK(clk),
    .QN(\text_out[112]_3072 ),
    .D(n_8287),
    .SE(w0[16]),
    .SI(n_174));
 SDFHx1_ASAP7_75t_R \text_out_reg[113]  (.CLK(clk),
    .QN(\text_out[113]_3073 ),
    .D(n_240),
    .SE(w0[17]),
    .SI(n_8313));
 SDFHx1_ASAP7_75t_R \text_out_reg[114]  (.CLK(clk),
    .QN(\text_out[114]_3074 ),
    .D(n_211),
    .SE(w0[18]),
    .SI(n_8312));
 SDFHx1_ASAP7_75t_R \text_out_reg[115]  (.CLK(clk),
    .QN(\text_out[115]_3075 ),
    .D(n_357),
    .SE(w0[19]),
    .SI(n_356));
 SDFHx1_ASAP7_75t_R \text_out_reg[116]  (.CLK(clk),
    .QN(\text_out[116]_3076 ),
    .D(n_355),
    .SE(w0[20]),
    .SI(n_8311));
 SDFHx1_ASAP7_75t_R \text_out_reg[117]  (.CLK(clk),
    .QN(\text_out[117]_3077 ),
    .D(n_8244),
    .SE(w0[21]),
    .SI(n_238));
 SDFHx1_ASAP7_75t_R \text_out_reg[118]  (.CLK(clk),
    .QN(\text_out[118]_3078 ),
    .D(n_8271),
    .SE(w0[22]),
    .SI(n_364));
 SDFHx1_ASAP7_75t_R \text_out_reg[119]  (.CLK(clk),
    .QN(\text_out[119]_3079 ),
    .D(n_8243),
    .SE(w0[23]),
    .SI(n_122));
 SDFHx1_ASAP7_75t_R \text_out_reg[11]  (.CLK(clk),
    .QN(\text_out[11]_3131 ),
    .D(n_7539),
    .SE(w3[11]),
    .SI(n_7540));
 SDFHx1_ASAP7_75t_R \text_out_reg[120]  (.CLK(clk),
    .QN(\text_out[120]_3040 ),
    .D(n_8283),
    .SE(w0[24]),
    .SI(n_214));
 SDFHx1_ASAP7_75t_R \text_out_reg[121]  (.CLK(clk),
    .QN(\text_out[121]_3041 ),
    .D(n_8879),
    .SE(w0[25]),
    .SI(n_8877));
 SDFHx1_ASAP7_75t_R \text_out_reg[122]  (.CLK(clk),
    .QN(\text_out[122]_3042 ),
    .D(n_235),
    .SE(w0[26]),
    .SI(n_8300));
 SDFHx1_ASAP7_75t_R \text_out_reg[123]  (.CLK(clk),
    .QN(\text_out[123]_3043 ),
    .D(n_7502),
    .SE(w0[27]),
    .SI(n_7503));
 SDFHx1_ASAP7_75t_R \text_out_reg[124]  (.CLK(clk),
    .QN(\text_out[124]_3044 ),
    .D(n_8792),
    .SE(w0[28]),
    .SI(n_8299));
 SDFHx1_ASAP7_75t_R \text_out_reg[125]  (.CLK(clk),
    .QN(\text_out[125]_3045 ),
    .D(n_8236),
    .SE(w0[29]),
    .SI(n_173));
 SDFHx1_ASAP7_75t_R \text_out_reg[126]  (.CLK(clk),
    .QN(\text_out[126]_3046 ),
    .D(n_8267),
    .SE(w0[30]),
    .SI(n_228));
 SDFHx1_ASAP7_75t_R \text_out_reg[127]  (.CLK(clk),
    .QN(\text_out[127]_3047 ),
    .D(n_7546),
    .SE(w0[31]),
    .SI(n_7547));
 SDFHx1_ASAP7_75t_R \text_out_reg[12]  (.CLK(clk),
    .QN(\text_out[12]_3132 ),
    .D(n_184),
    .SE(w3[12]),
    .SI(n_8332));
 SDFHx1_ASAP7_75t_R \text_out_reg[13]  (.CLK(clk),
    .QN(\text_out[13]_3133 ),
    .D(n_8258),
    .SE(w3[13]),
    .SI(n_242));
 SDFHx1_ASAP7_75t_R \text_out_reg[14]  (.CLK(clk),
    .QN(\text_out[14]_3134 ),
    .D(w3[14]),
    .SE(n_8278),
    .SI(n_8801));
 SDFHx1_ASAP7_75t_R \text_out_reg[15]  (.CLK(clk),
    .QN(\text_out[15]_3135 ),
    .D(n_7447),
    .SE(w3[15]),
    .SI(n_7448));
 SDFHx1_ASAP7_75t_R \text_out_reg[16]  (.CLK(clk),
    .QN(\text_out[16]_3096 ),
    .D(n_8290),
    .SE(w3[16]),
    .SI(n_156));
 SDFHx1_ASAP7_75t_R \text_out_reg[17]  (.CLK(clk),
    .QN(\text_out[17]_3097 ),
    .D(n_292),
    .SE(w3[17]),
    .SI(n_8322));
 SDFHx1_ASAP7_75t_R \text_out_reg[18]  (.CLK(clk),
    .QN(\text_out[18]_3098 ),
    .D(n_154),
    .SE(w3[18]),
    .SI(n_8321));
 SDFHx1_ASAP7_75t_R \text_out_reg[19]  (.CLK(clk),
    .QN(\text_out[19]_3099 ),
    .D(n_8226),
    .SE(n_8668),
    .SI(n_208));
 SDFHx1_ASAP7_75t_R \text_out_reg[1]  (.CLK(clk),
    .QN(\text_out[1]_3161 ),
    .D(n_125),
    .SE(n_8748),
    .SI(n_8344));
 SDFHx1_ASAP7_75t_R \text_out_reg[20]  (.CLK(clk),
    .QN(\text_out[20]_3100 ),
    .D(n_350),
    .SE(w3[20]),
    .SI(n_8320));
 SDFHx1_ASAP7_75t_R \text_out_reg[21]  (.CLK(clk),
    .QN(\text_out[21]_3101 ),
    .D(n_8250),
    .SE(w3[21]),
    .SI(n_221));
 SDFHx1_ASAP7_75t_R \text_out_reg[22]  (.CLK(clk),
    .QN(\text_out[22]_3102 ),
    .D(n_8274),
    .SE(w3[22]),
    .SI(n_153));
 SDFHx1_ASAP7_75t_R \text_out_reg[23]  (.CLK(clk),
    .QN(\text_out[23]_3103 ),
    .D(n_8249),
    .SE(n_8831),
    .SI(n_338));
 SDFHx1_ASAP7_75t_R \text_out_reg[24]  (.CLK(clk),
    .QN(\text_out[24]_3064 ),
    .D(n_8286),
    .SE(w3[24]),
    .SI(n_222));
 SDFHx1_ASAP7_75t_R \text_out_reg[25]  (.CLK(clk),
    .QN(\text_out[25]_3065 ),
    .D(n_159),
    .SE(w3[25]),
    .SI(n_8310));
 SDFHx1_ASAP7_75t_R \text_out_reg[26]  (.CLK(clk),
    .QN(\text_out[26]_3066 ),
    .D(n_7556),
    .SE(w3[26]),
    .SI(n_8309));
 SDFHx1_ASAP7_75t_R \text_out_reg[27]  (.CLK(clk),
    .QN(\text_out[27]_3067 ),
    .D(n_8222),
    .SE(w3[27]),
    .SI(n_152));
 SDFHx1_ASAP7_75t_R \text_out_reg[28]  (.CLK(clk),
    .QN(\text_out[28]_3068 ),
    .D(n_196),
    .SE(n_8942),
    .SI(n_8308));
 SDFHx1_ASAP7_75t_R \text_out_reg[29]  (.CLK(clk),
    .QN(\text_out[29]_3069 ),
    .D(n_8242),
    .SE(w3[29]),
    .SI(n_349));
 SDFHx1_ASAP7_75t_R \text_out_reg[2]  (.CLK(clk),
    .QN(\text_out[2]_3162 ),
    .D(n_166),
    .SE(w3[2]),
    .SI(n_8346));
 SDFHx1_ASAP7_75t_R \text_out_reg[30]  (.CLK(clk),
    .QN(\text_out[30]_3070 ),
    .D(n_8270),
    .SE(w3[30]),
    .SI(n_158));
 SDFHx1_ASAP7_75t_R \text_out_reg[31]  (.CLK(clk),
    .QN(\text_out[31]_3071 ),
    .D(n_7491),
    .SE(w3[31]),
    .SI(n_7492));
 SDFHx1_ASAP7_75t_R \text_out_reg[32]  (.CLK(clk),
    .QN(\text_out[32]_3152 ),
    .D(n_7494),
    .SE(w2[0]),
    .SI(n_7495));
 SDFHx1_ASAP7_75t_R \text_out_reg[33]  (.CLK(clk),
    .QN(\text_out[33]_3153 ),
    .D(n_136),
    .SE(w2[1]),
    .SI(n_8343));
 SDFHx1_ASAP7_75t_R \text_out_reg[34]  (.CLK(clk),
    .QN(\text_out[34]_3154 ),
    .D(n_195),
    .SE(w2[2]),
    .SI(n_8342));
 SDFHx1_ASAP7_75t_R \text_out_reg[35]  (.CLK(clk),
    .QN(\text_out[35]_3155 ),
    .D(n_7541),
    .SE(w2[3]),
    .SI(n_7542));
 SDFHx1_ASAP7_75t_R \text_out_reg[36]  (.CLK(clk),
    .QN(\text_out[36]_3156 ),
    .D(n_49),
    .SE(w2[4]),
    .SI(n_129));
 SDFHx1_ASAP7_75t_R \text_out_reg[37]  (.CLK(clk),
    .QN(\text_out[37]_3157 ),
    .D(n_7584),
    .SE(w2[5]),
    .SI(n_7585));
 SDFHx1_ASAP7_75t_R \text_out_reg[38]  (.CLK(clk),
    .QN(\text_out[38]_3158 ),
    .D(n_8281),
    .SE(w2[6]),
    .SI(n_145));
 SDFHx1_ASAP7_75t_R \text_out_reg[39]  (.CLK(clk),
    .QN(\text_out[39]_3159 ),
    .D(n_121),
    .SE(w2[7]),
    .SI(n_42));
 SDFHx1_ASAP7_75t_R \text_out_reg[3]  (.CLK(clk),
    .QN(\text_out[3]_3163 ),
    .D(n_8887),
    .SE(w3[3]),
    .SI(n_8884));
 SDFHx1_ASAP7_75t_R \text_out_reg[40]  (.CLK(clk),
    .QN(\text_out[40]_3120 ),
    .D(n_8293),
    .SE(w2[8]),
    .SI(n_60));
 SDFHx1_ASAP7_75t_R \text_out_reg[41]  (.CLK(clk),
    .QN(\text_out[41]_3121 ),
    .D(n_223),
    .SE(w2[9]),
    .SI(n_8331));
 SDFHx1_ASAP7_75t_R \text_out_reg[42]  (.CLK(clk),
    .QN(\text_out[42]_3122 ),
    .D(n_189),
    .SE(w2[10]),
    .SI(n_8330));
 SDFHx1_ASAP7_75t_R \text_out_reg[43]  (.CLK(clk),
    .QN(\text_out[43]_3123 ),
    .D(n_8229),
    .SE(w2[11]),
    .SI(n_226));
 SDFHx1_ASAP7_75t_R \text_out_reg[44]  (.CLK(clk),
    .QN(\text_out[44]_3124 ),
    .D(n_347),
    .SE(w2[12]),
    .SI(n_8329));
 SDFHx1_ASAP7_75t_R \text_out_reg[45]  (.CLK(clk),
    .QN(\text_out[45]_3125 ),
    .D(n_8256),
    .SE(w2[13]),
    .SI(n_59));
 SDFHx1_ASAP7_75t_R \text_out_reg[46]  (.CLK(clk),
    .QN(\text_out[46]_3126 ),
    .D(n_8277),
    .SE(w2[14]),
    .SI(n_341));
 SDFHx1_ASAP7_75t_R \text_out_reg[47]  (.CLK(clk),
    .QN(\text_out[47]_3127 ),
    .D(n_8255),
    .SE(w2[15]),
    .SI(n_127));
 SDFHx1_ASAP7_75t_R \text_out_reg[48]  (.CLK(clk),
    .QN(\text_out[48]_3088 ),
    .D(n_7450),
    .SE(w2[16]),
    .SI(n_7451));
 SDFHx1_ASAP7_75t_R \text_out_reg[49]  (.CLK(clk),
    .QN(\text_out[49]_3089 ),
    .D(n_363),
    .SE(w2[17]),
    .SI(n_8319));
 SDFHx1_ASAP7_75t_R \text_out_reg[4]  (.CLK(clk),
    .QN(\text_out[4]_3164 ),
    .D(n_47),
    .SE(n_8629),
    .SI(n_8345));
 SDFHx1_ASAP7_75t_R \text_out_reg[50]  (.CLK(clk),
    .QN(\text_out[50]_3090 ),
    .D(n_187),
    .SE(w2[18]),
    .SI(n_8318));
 SDFHx1_ASAP7_75t_R \text_out_reg[51]  (.CLK(clk),
    .QN(\text_out[51]_3091 ),
    .D(n_8225),
    .SE(w2[19]),
    .SI(n_7560));
 SDFHx1_ASAP7_75t_R \text_out_reg[52]  (.CLK(clk),
    .QN(\text_out[52]_3092 ),
    .D(n_239),
    .SE(w2[20]),
    .SI(n_8317));
 SDFHx1_ASAP7_75t_R \text_out_reg[53]  (.CLK(clk),
    .QN(\text_out[53]_3093 ),
    .D(n_7548),
    .SE(w2[21]),
    .SI(n_7549));
 SDFHx1_ASAP7_75t_R \text_out_reg[54]  (.CLK(clk),
    .QN(\text_out[54]_3094 ),
    .D(n_8273),
    .SE(w2[22]),
    .SI(n_351));
 SDFHx1_ASAP7_75t_R \text_out_reg[55]  (.CLK(clk),
    .QN(\text_out[55]_3095 ),
    .D(n_8247),
    .SE(w2[23]),
    .SI(n_330));
 SDFHx1_ASAP7_75t_R \text_out_reg[56]  (.CLK(clk),
    .QN(\text_out[56]_3056 ),
    .D(n_8285),
    .SE(w2[24]),
    .SI(n_229));
 SDFHx1_ASAP7_75t_R \text_out_reg[57]  (.CLK(clk),
    .QN(\text_out[57]_3057 ),
    .D(n_8771),
    .SE(w2[25]),
    .SI(n_8770));
 SDFHx1_ASAP7_75t_R \text_out_reg[58]  (.CLK(clk),
    .QN(\text_out[58]_3058 ),
    .D(n_53),
    .SE(w2[26]),
    .SI(n_169));
 SDFHx1_ASAP7_75t_R \text_out_reg[59]  (.CLK(clk),
    .QN(\text_out[59]_3059 ),
    .D(n_8733),
    .SE(w2[27]),
    .SI(n_8732));
 SDFHx1_ASAP7_75t_R \text_out_reg[5]  (.CLK(clk),
    .QN(\text_out[5]_3165 ),
    .D(n_8266),
    .SE(w3[5]),
    .SI(n_190));
 SDFHx1_ASAP7_75t_R \text_out_reg[60]  (.CLK(clk),
    .QN(\text_out[60]_3060 ),
    .D(n_191),
    .SE(w2[28]),
    .SI(n_8305));
 SDFHx1_ASAP7_75t_R \text_out_reg[61]  (.CLK(clk),
    .QN(\text_out[61]_3061 ),
    .D(n_7588),
    .SE(w2[29]),
    .SI(n_7589));
 SDFHx1_ASAP7_75t_R \text_out_reg[62]  (.CLK(clk),
    .QN(\text_out[62]_3062 ),
    .D(n_8269),
    .SE(w2[30]),
    .SI(n_151));
 SDFHx1_ASAP7_75t_R \text_out_reg[63]  (.CLK(clk),
    .QN(\text_out[63]_3063 ),
    .D(n_8783),
    .SE(w2[31]),
    .SI(n_8785));
 SDFHx1_ASAP7_75t_R \text_out_reg[64]  (.CLK(clk),
    .QN(\text_out[64]_3144 ),
    .D(n_8296),
    .SE(w1[0]),
    .SI(n_177));
 SDFHx1_ASAP7_75t_R \text_out_reg[65]  (.CLK(clk),
    .QN(\text_out[65]_3145 ),
    .D(n_7507),
    .SE(w1[1]),
    .SI(n_8340));
 SDFHx1_ASAP7_75t_R \text_out_reg[66]  (.CLK(clk),
    .QN(\text_out[66]_3146 ),
    .D(n_7533),
    .SE(w1[2]),
    .SI(n_8339));
 SDFHx1_ASAP7_75t_R \text_out_reg[67]  (.CLK(clk),
    .QN(\text_out[67]_3147 ),
    .D(n_8232),
    .SE(w1[3]),
    .SI(n_7550));
 SDFHx1_ASAP7_75t_R \text_out_reg[68]  (.CLK(clk),
    .QN(\text_out[68]_3148 ),
    .D(n_134),
    .SE(w1[4]),
    .SI(n_8338));
 SDFHx1_ASAP7_75t_R \text_out_reg[69]  (.CLK(clk),
    .QN(\text_out[69]_3149 ),
    .D(n_8262),
    .SE(w1[5]),
    .SI(n_143));
 SDFHx1_ASAP7_75t_R \text_out_reg[6]  (.CLK(clk),
    .QN(\text_out[6]_3166 ),
    .D(n_1800),
    .SE(w3[6]),
    .SI(n_7602));
 SDFHx1_ASAP7_75t_R \text_out_reg[70]  (.CLK(clk),
    .QN(\text_out[70]_3150 ),
    .D(n_8280),
    .SE(w1[6]),
    .SI(n_8723));
 SDFHx1_ASAP7_75t_R \text_out_reg[71]  (.CLK(clk),
    .QN(\text_out[71]_3151 ),
    .D(n_8932),
    .SE(w1[7]),
    .SI(n_8933));
 SDFHx1_ASAP7_75t_R \text_out_reg[72]  (.CLK(clk),
    .QN(\text_out[72]_3112 ),
    .D(n_207),
    .SE(w1[8]),
    .SI(n_206));
 SDFHx1_ASAP7_75t_R \text_out_reg[73]  (.CLK(clk),
    .QN(\text_out[73]_3113 ),
    .D(n_217),
    .SE(w1[9]),
    .SI(n_8328));
 SDFHx1_ASAP7_75t_R \text_out_reg[74]  (.CLK(clk),
    .QN(\text_out[74]_3114 ),
    .D(n_346),
    .SE(w1[10]),
    .SI(n_8327));
 SDFHx1_ASAP7_75t_R \text_out_reg[75]  (.CLK(clk),
    .QN(\text_out[75]_3115 ),
    .D(n_8228),
    .SE(w1[11]),
    .SI(n_202));
 SDFHx1_ASAP7_75t_R \text_out_reg[76]  (.CLK(clk),
    .QN(\text_out[76]_3116 ),
    .D(n_230),
    .SE(w1[12]),
    .SI(n_8326));
 SDFHx1_ASAP7_75t_R \text_out_reg[77]  (.CLK(clk),
    .QN(\text_out[77]_3117 ),
    .D(n_8254),
    .SE(w1[13]),
    .SI(n_135));
 SDFHx1_ASAP7_75t_R \text_out_reg[78]  (.CLK(clk),
    .QN(\text_out[78]_3118 ),
    .D(n_8276),
    .SE(w1[14]),
    .SI(n_165));
 SDFHx1_ASAP7_75t_R \text_out_reg[79]  (.CLK(clk),
    .QN(\text_out[79]_3119 ),
    .D(n_8766),
    .SE(w1[15]),
    .SI(n_8760));
 SDFHx1_ASAP7_75t_R \text_out_reg[7]  (.CLK(clk),
    .QN(\text_out[7]_3167 ),
    .D(n_117),
    .SE(w3[7]),
    .SI(n_116));
 SDFHx1_ASAP7_75t_R \text_out_reg[80]  (.CLK(clk),
    .QN(\text_out[80]_3080 ),
    .D(n_37),
    .SE(w1[16]),
    .SI(n_167));
 SDFHx1_ASAP7_75t_R \text_out_reg[81]  (.CLK(clk),
    .QN(\text_out[81]_3081 ),
    .D(n_283),
    .SE(w1[17]),
    .SI(n_8316));
 SDFHx1_ASAP7_75t_R \text_out_reg[82]  (.CLK(clk),
    .QN(\text_out[82]_3082 ),
    .D(n_232),
    .SE(w1[18]),
    .SI(n_8315));
 SDFHx1_ASAP7_75t_R \text_out_reg[83]  (.CLK(clk),
    .QN(\text_out[83]_3083 ),
    .D(n_8224),
    .SE(w1[19]),
    .SI(n_234));
 SDFHx1_ASAP7_75t_R \text_out_reg[84]  (.CLK(clk),
    .QN(\text_out[84]_3084 ),
    .D(n_371),
    .SE(w1[20]),
    .SI(n_8314));
 SDFHx1_ASAP7_75t_R \text_out_reg[85]  (.CLK(clk),
    .QN(\text_out[85]_3085 ),
    .D(n_7573),
    .SE(w1[21]),
    .SI(n_7574));
 SDFHx1_ASAP7_75t_R \text_out_reg[86]  (.CLK(clk),
    .QN(\text_out[86]_3086 ),
    .D(n_8272),
    .SE(w1[22]),
    .SI(n_199));
 SDFHx1_ASAP7_75t_R \text_out_reg[87]  (.CLK(clk),
    .QN(\text_out[87]_3087 ),
    .D(n_8245),
    .SE(w1[23]),
    .SI(n_8679));
 SDFHx1_ASAP7_75t_R \text_out_reg[88]  (.CLK(clk),
    .QN(\text_out[88]_3048 ),
    .D(n_7474),
    .SE(w1[24]),
    .SI(n_7475));
 SDFHx1_ASAP7_75t_R \text_out_reg[89]  (.CLK(clk),
    .QN(\text_out[89]_3049 ),
    .D(n_348),
    .SE(w1[25]),
    .SI(n_8304));
 SDFHx1_ASAP7_75t_R \text_out_reg[8]  (.CLK(clk),
    .QN(\text_out[8]_3128 ),
    .D(n_7513),
    .SE(n_11401),
    .SI(n_7514));
 SDFHx1_ASAP7_75t_R \text_out_reg[90]  (.CLK(clk),
    .QN(\text_out[90]_3050 ),
    .D(n_237),
    .SE(w1[26]),
    .SI(n_8303));
 SDFHx1_ASAP7_75t_R \text_out_reg[91]  (.CLK(clk),
    .QN(\text_out[91]_3051 ),
    .D(n_8220),
    .SE(w1[27]),
    .SI(n_168));
 SDFHx1_ASAP7_75t_R \text_out_reg[92]  (.CLK(clk),
    .QN(\text_out[92]_3052 ),
    .D(n_345),
    .SE(w1[28]),
    .SI(n_8302));
 SDFHx1_ASAP7_75t_R \text_out_reg[93]  (.CLK(clk),
    .QN(\text_out[93]_3053 ),
    .D(n_8238),
    .SE(w1[29]),
    .SI(n_209));
 SDFHx1_ASAP7_75t_R \text_out_reg[94]  (.CLK(clk),
    .QN(\text_out[94]_3054 ),
    .D(n_8268),
    .SE(w1[30]),
    .SI(n_172));
 SDFHx1_ASAP7_75t_R \text_out_reg[95]  (.CLK(clk),
    .QN(\text_out[95]_3055 ),
    .D(n_131),
    .SE(w1[31]),
    .SI(n_130));
 SDFHx1_ASAP7_75t_R \text_out_reg[96]  (.CLK(clk),
    .QN(\text_out[96]_3136 ),
    .D(n_8295),
    .SE(w0[0]),
    .SI(n_175));
 SDFHx1_ASAP7_75t_R \text_out_reg[97]  (.CLK(clk),
    .QN(\text_out[97]_3137 ),
    .D(n_340),
    .SE(w0[1]),
    .SI(n_8337));
 SDFHx1_ASAP7_75t_R \text_out_reg[98]  (.CLK(clk),
    .QN(\text_out[98]_3138 ),
    .D(n_233),
    .SE(w0[2]),
    .SI(n_8336));
 SDFHx1_ASAP7_75t_R \text_out_reg[99]  (.CLK(clk),
    .QN(\text_out[99]_3139 ),
    .D(n_8231),
    .SE(w0[3]),
    .SI(n_186));
 SDFHx1_ASAP7_75t_R \text_out_reg[9]  (.CLK(clk),
    .QN(\text_out[9]_3129 ),
    .D(n_362),
    .SE(n_8856),
    .SI(n_8334));
 INVx1_ASAP7_75t_R u0_drc_bufs (.A(u0_n_32835),
    .Y(u0_n_32834));
 INVx2_ASAP7_75t_R u0_drc_bufs64517 (.A(u0_n_32835),
    .Y(u0_n_32843));
 INVxp67_ASAP7_75t_R u0_drc_bufs64518 (.A(u0_n_32835),
    .Y(u0_n_32851));
 INVx2_ASAP7_75t_SL u0_drc_bufs64519 (.A(ld),
    .Y(u0_n_32835));
 INVx1_ASAP7_75t_R u0_drc_bufs64528 (.A(u0_n_32836),
    .Y(u0_n_32966));
 INVxp33_ASAP7_75t_R u0_drc_bufs64529 (.A(u0_n_32836),
    .Y(u0_n_32967));
 INVxp67_ASAP7_75t_R u0_drc_bufs64533 (.A(u0_n_32836),
    .Y(u0_n_32971));
 INVx1_ASAP7_75t_R u0_drc_bufs64545 (.A(u0_n_32834),
    .Y(u0_n_32983));
 INVxp67_ASAP7_75t_R u0_drc_bufs64552 (.A(u0_n_32835),
    .Y(u0_n_32990));
 INVxp33_ASAP7_75t_R u0_drc_bufs64553 (.A(u0_n_32835),
    .Y(u0_n_32991));
 HB1xp67_ASAP7_75t_L u0_drc_bufs64638 (.A(\u0_w[3] [27]),
    .Y(w3[27]));
 HB1xp67_ASAP7_75t_R u0_drc_bufs64644 (.A(u0_n_32825),
    .Y(u0_n_33110));
 BUFx2_ASAP7_75t_L u0_drc_bufs64652 (.A(\u0_w[3] [12]),
    .Y(w3[12]));
 HB1xp67_ASAP7_75t_R u0_drc_bufs64658 (.A(\u0_w[3] [16]),
    .Y(w3[16]));
 INVx1_ASAP7_75t_L u0_fopt1 (.A(u0_n_33008),
    .Y(u0_n_33001));
 INVx1_ASAP7_75t_R u0_fopt12 (.A(w3[22]),
    .Y(u0_n_33008));
 BUFx3_ASAP7_75t_SL u0_fopt14 (.A(\u0_w[3] [22]),
    .Y(w3[22]));
 INVx1_ASAP7_75t_L u0_fopt64580 (.A(u0_n_33030),
    .Y(u0_n_33033));
 INVxp67_ASAP7_75t_R u0_fopt64581 (.A(w3[30]),
    .Y(u0_n_33030));
 BUFx2_ASAP7_75t_L u0_fopt64582 (.A(\u0_w[3] [30]),
    .Y(w3[30]));
 INVx2_ASAP7_75t_L u0_fopt64679 (.A(w3[20]),
    .Y(u0_n_33138));
 INVxp67_ASAP7_75t_R u0_fopt8 (.A(u0_n_33008),
    .Y(u0_n_33004));
 AO221x1_ASAP7_75t_L u0_g2 (.A1(u0_n_31272),
    .A2(u0_n_32012),
    .B1(u0_n_31240),
    .B2(u0_n_32260),
    .C(u0_n_30967),
    .Y(u0_n_33149));
 AOI22xp5_ASAP7_75t_SL u0_g61910 (.A1(u0_n_29305),
    .A2(u0_n_32924),
    .B1(key[56]),
    .B2(u0_n_32843),
    .Y(u0_n_29279));
 AO21x1_ASAP7_75t_SL u0_g61911 (.A1(key[13]),
    .A2(u0_n_32836),
    .B(u0_n_29281),
    .Y(u0_n_29280));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g61933 (.A1(w3[13]),
    .A2(u0_n_29394),
    .B(u0_n_29322),
    .C(u0_n_32843),
    .Y(u0_n_29281));
 AOI22xp33_ASAP7_75t_L u0_g61934 (.A1(u0_n_32924),
    .A2(u0_n_29368),
    .B1(key[62]),
    .B2(u0_n_32934),
    .Y(u0_n_29283));
 AOI22xp5_ASAP7_75t_SL u0_g61935 (.A1(u0_n_32924),
    .A2(u0_n_29350),
    .B1(key[36]),
    .B2(u0_n_32934),
    .Y(u0_n_29284));
 AOI22xp5_ASAP7_75t_SL u0_g61936 (.A1(u0_n_32924),
    .A2(u0_n_29345),
    .B1(key[34]),
    .B2(u0_n_32934),
    .Y(u0_n_29285));
 AOI22xp33_ASAP7_75t_SL u0_g61937 (.A1(u0_n_32835),
    .A2(u0_n_29364),
    .B1(key[94]),
    .B2(u0_n_32843),
    .Y(u0_n_29286));
 AOI22xp5_ASAP7_75t_SL u0_g61949 (.A1(u0_n_32924),
    .A2(u0_n_29414),
    .B1(key[43]),
    .B2(u0_n_32836),
    .Y(u0_n_29287));
 AOI22xp5_ASAP7_75t_SL u0_g61950 (.A1(u0_n_32839),
    .A2(u0_n_29436),
    .B1(key[90]),
    .B2(u0_n_32843),
    .Y(u0_n_29288));
 AO21x1_ASAP7_75t_SL u0_g61951 (.A1(key[29]),
    .A2(u0_n_32836),
    .B(u0_n_29330),
    .Y(u0_n_29289));
 AOI22xp5_ASAP7_75t_SL u0_g61968 (.A1(u0_n_32839),
    .A2(u0_n_29418),
    .B1(key[50]),
    .B2(u0_n_32942),
    .Y(u0_n_29290));
 AOI22xp5_ASAP7_75t_SL u0_g61969 (.A1(u0_n_32924),
    .A2(u0_n_29440),
    .B1(key[58]),
    .B2(u0_n_32934),
    .Y(u0_n_29291));
 AOI22xp5_ASAP7_75t_SL u0_g61970 (.A1(u0_n_32971),
    .A2(u0_n_29421),
    .B1(key[59]),
    .B2(u0_n_32942),
    .Y(u0_n_29292));
 AOI22xp5_ASAP7_75t_R u0_g61971 (.A1(u0_n_32875),
    .A2(u0_n_29424),
    .B1(key[61]),
    .B2(u0_n_32942),
    .Y(u0_n_29293));
 AOI22xp5_ASAP7_75t_SL u0_g61972 (.A1(u0_n_32839),
    .A2(u0_n_29426),
    .B1(key[63]),
    .B2(u0_n_32934),
    .Y(u0_n_29294));
 AO21x1_ASAP7_75t_SL u0_g61973 (.A1(key[5]),
    .A2(u0_n_32834),
    .B(u0_n_29332),
    .Y(u0_n_29295));
 AO21x1_ASAP7_75t_SL u0_g61974 (.A1(key[26]),
    .A2(u0_n_32836),
    .B(u0_n_29331),
    .Y(u0_n_29296));
 AOI22xp33_ASAP7_75t_R u0_g61975 (.A1(u0_n_32983),
    .A2(u0_n_29396),
    .B1(key[88]),
    .B2(u0_n_32845),
    .Y(u0_n_29297));
 AOI22xp33_ASAP7_75t_R u0_g61976 (.A1(u0_n_32879),
    .A2(u0_n_29395),
    .B1(key[32]),
    .B2(u0_n_32991),
    .Y(u0_n_29298));
 AOI22xp33_ASAP7_75t_R u0_g61977 (.A1(u0_n_32983),
    .A2(u0_n_29391),
    .B1(key[40]),
    .B2(u0_n_33110),
    .Y(u0_n_29299));
 AOI22xp33_ASAP7_75t_SL u0_g61978 (.A1(u0_n_32983),
    .A2(u0_n_29393),
    .B1(key[45]),
    .B2(u0_n_32990),
    .Y(u0_n_29300));
 AOI22xp33_ASAP7_75t_L u0_g61979 (.A1(u0_n_32875),
    .A2(n_8847),
    .B1(key[48]),
    .B2(u0_n_32845),
    .Y(u0_n_29301));
 AOI22xp33_ASAP7_75t_R u0_g61980 (.A1(u0_n_32877),
    .A2(u0_n_29392),
    .B1(key[53]),
    .B2(u0_n_32991),
    .Y(u0_n_29302));
 AOI322xp5_ASAP7_75t_SL u0_g61981 (.A1(u0_n_29477),
    .A2(w2[28]),
    .A3(u0_n_32835),
    .B1(u0_n_32571),
    .B2(u0_n_29372),
    .C1(key[60]),
    .C2(u0_n_32843),
    .Y(u0_n_29303));
 XOR2xp5_ASAP7_75t_SL u0_g61982 (.A(u0_n_29396),
    .B(w2[24]),
    .Y(u0_n_29305));
 XNOR2xp5_ASAP7_75t_SL u0_g61983 (.A(u0_n_29395),
    .B(w3[0]),
    .Y(u0_n_29308));
 XNOR2xp5_ASAP7_75t_SL u0_g61984 (.A(u0_n_29391),
    .B(n_11401),
    .Y(u0_n_29311));
 AOI22xp5_ASAP7_75t_SL u0_g61985 (.A1(\u0_w[3] [16]),
    .A2(u0_n_29390),
    .B1(u0_n_32753),
    .B2(n_8847),
    .Y(u0_n_29314));
 XNOR2xp5_ASAP7_75t_SL u0_g61986 (.A(u0_n_29392),
    .B(w3[21]),
    .Y(u0_n_29317));
 XNOR2xp5_ASAP7_75t_L u0_g61987 (.A(u0_n_29397),
    .B(u0_n_31722),
    .Y(u0_n_29320));
 AOI22xp33_ASAP7_75t_L u0_g61988 (.A1(u0_n_32839),
    .A2(u0_n_29500),
    .B1(key[70]),
    .B2(u0_n_32825),
    .Y(u0_n_29321));
 NAND2xp5_ASAP7_75t_SL u0_g61989 (.A(u0_n_29394),
    .B(w3[13]),
    .Y(u0_n_29322));
 XNOR2xp5_ASAP7_75t_SL u0_g62018 (.A(u0_n_29468),
    .B(u0_n_32774),
    .Y(u0_n_29324));
 AOI21xp5_ASAP7_75t_R u0_g62019 (.A1(key[92]),
    .A2(u0_n_32834),
    .B(u0_n_29372),
    .Y(u0_n_29326));
 AOI22xp33_ASAP7_75t_L u0_g62020 (.A1(u0_n_32879),
    .A2(u0_n_29506),
    .B1(key[47]),
    .B2(u0_n_32942),
    .Y(u0_n_29328));
 AOI22xp5_ASAP7_75t_L u0_g62021 (.A1(u0_n_32879),
    .A2(u0_n_29498),
    .B1(key[52]),
    .B2(u0_n_32934),
    .Y(u0_n_29329));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62022 (.A1(u0_n_31574),
    .A2(u0_n_29563),
    .B(u0_n_29463),
    .C(u0_n_32836),
    .Y(u0_n_29330));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62023 (.A1(u0_n_30904),
    .A2(u0_n_29521),
    .B(u0_n_29465),
    .C(u0_n_32836),
    .Y(u0_n_29331));
 AOI221xp5_ASAP7_75t_SL u0_g62024 (.A1(u0_n_29550),
    .A2(u0_n_32691),
    .B1(w3[5]),
    .B2(u0_n_29549),
    .C(u0_n_32843),
    .Y(u0_n_29332));
 AOI22xp33_ASAP7_75t_R u0_g62025 (.A1(u0_n_32877),
    .A2(u0_n_29482),
    .B1(key[126]),
    .B2(u0_n_32845),
    .Y(u0_n_29334));
 AOI22xp33_ASAP7_75t_R u0_g62026 (.A1(u0_n_32983),
    .A2(u0_n_29480),
    .B1(key[66]),
    .B2(u0_n_32990),
    .Y(u0_n_29335));
 AOI22xp33_ASAP7_75t_R u0_g62027 (.A1(u0_n_32983),
    .A2(u0_n_29478),
    .B1(key[68]),
    .B2(u0_n_32991),
    .Y(u0_n_29336));
 AOI22xp33_ASAP7_75t_L u0_g62028 (.A1(u0_n_32877),
    .A2(u0_n_29475),
    .B1(key[79]),
    .B2(u0_n_32836),
    .Y(u0_n_29337));
 AOI22xp33_ASAP7_75t_L u0_g62029 (.A1(u0_n_32967),
    .A2(u0_n_29473),
    .B1(key[33]),
    .B2(u0_n_32991),
    .Y(u0_n_29338));
 AOI22xp33_ASAP7_75t_R u0_g62030 (.A1(u0_n_32967),
    .A2(u0_n_29468),
    .B1(key[38]),
    .B2(u0_n_32991),
    .Y(u0_n_29339));
 AOI22xp33_ASAP7_75t_L u0_g62031 (.A1(u0_n_32966),
    .A2(u0_n_29469),
    .B1(key[39]),
    .B2(u0_n_32845),
    .Y(u0_n_29341));
 AOI22xp33_ASAP7_75t_R u0_g62032 (.A1(u0_n_32877),
    .A2(u0_n_29471),
    .B1(key[41]),
    .B2(u0_n_32990),
    .Y(u0_n_29342));
 AOI22xp33_ASAP7_75t_R u0_g62033 (.A1(u0_n_32879),
    .A2(u0_n_29472),
    .B1(key[44]),
    .B2(u0_n_32991),
    .Y(u0_n_29343));
 XNOR2xp5_ASAP7_75t_L u0_g62034 (.A(u0_n_29481),
    .B(u0_n_31076),
    .Y(u0_n_29344));
 XOR2xp5_ASAP7_75t_L u0_g62035 (.A(u0_n_29480),
    .B(w2[2]),
    .Y(u0_n_29345));
 XNOR2xp5_ASAP7_75t_SL u0_g62036 (.A(u0_n_31727),
    .B(u0_n_29477),
    .Y(u0_n_29348));
 XOR2xp5_ASAP7_75t_SL u0_g62037 (.A(u0_n_29478),
    .B(w2[4]),
    .Y(u0_n_29350));
 XOR2xp5_ASAP7_75t_SL u0_g62038 (.A(u0_n_29474),
    .B(n_8748),
    .Y(u0_n_29353));
 XNOR2xp5_ASAP7_75t_SL u0_g62039 (.A(u0_n_29480),
    .B(u0_n_31720),
    .Y(u0_n_29355));
 XNOR2xp5_ASAP7_75t_R u0_g62040 (.A(u0_n_29479),
    .B(u0_n_31724),
    .Y(u0_n_29356));
 XNOR2xp5_ASAP7_75t_SL u0_g62041 (.A(u0_n_29471),
    .B(n_8856),
    .Y(u0_n_29357));
 XNOR2xp5_ASAP7_75t_SL u0_g62042 (.A(u0_n_29472),
    .B(\u0_w[3] [12]),
    .Y(u0_n_29360));
 XOR2xp5_ASAP7_75t_SL u0_g62043 (.A(u0_n_29476),
    .B(u0_n_31715),
    .Y(u0_n_29363));
 OAI22xp5_ASAP7_75t_SL u0_g62044 (.A1(u0_n_32676),
    .A2(u0_n_29482),
    .B1(w1[30]),
    .B2(u0_n_29481),
    .Y(u0_n_29364));
 XOR2xp5_ASAP7_75t_L u0_g62045 (.A(u0_n_29481),
    .B(u0_n_31709),
    .Y(u0_n_29368));
 XOR2xp5_ASAP7_75t_L u0_g62046 (.A(u0_n_29470),
    .B(w3[7]),
    .Y(u0_n_29369));
 AOI22xp33_ASAP7_75t_R u0_g62047 (.A1(u0_n_32966),
    .A2(u0_n_29503),
    .B1(key[71]),
    .B2(u0_n_32934),
    .Y(u0_n_29371));
 AOI22xp5_ASAP7_75t_R u0_g62048 (.A1(u0_n_32967),
    .A2(u0_n_29524),
    .B1(key[121]),
    .B2(u0_n_32942),
    .Y(u0_n_29373));
 AOI22xp33_ASAP7_75t_R u0_g62049 (.A1(u0_n_32877),
    .A2(u0_n_29551),
    .B1(key[80]),
    .B2(u0_n_32991),
    .Y(u0_n_29374));
 AOI22xp33_ASAP7_75t_R u0_g62050 (.A1(u0_n_32877),
    .A2(u0_n_29552),
    .B1(key[77]),
    .B2(u0_n_32825),
    .Y(u0_n_29375));
 AOI22xp33_ASAP7_75t_L u0_g62051 (.A1(u0_n_32971),
    .A2(u0_n_29561),
    .B1(key[75]),
    .B2(u0_n_32942),
    .Y(u0_n_29376));
 AOI22xp33_ASAP7_75t_R u0_g62052 (.A1(u0_n_32966),
    .A2(u0_n_29562),
    .B1(key[72]),
    .B2(u0_n_32991),
    .Y(u0_n_29377));
 AOI22xp33_ASAP7_75t_R u0_g62053 (.A1(u0_n_32966),
    .A2(u0_n_29547),
    .B1(key[64]),
    .B2(u0_n_32991),
    .Y(u0_n_29378));
 AOI22xp33_ASAP7_75t_L u0_g62054 (.A1(u0_n_32967),
    .A2(u0_n_29522),
    .B1(key[122]),
    .B2(u0_n_32990),
    .Y(u0_n_29379));
 AOI22xp33_ASAP7_75t_R u0_g62055 (.A1(u0_n_32879),
    .A2(u0_n_29520),
    .B1(key[120]),
    .B2(u0_n_32991),
    .Y(u0_n_29380));
 AO21x1_ASAP7_75t_SL u0_g62056 (.A1(key[10]),
    .A2(u0_n_32836),
    .B(u0_n_29467),
    .Y(u0_n_29381));
 AOI22xp5_ASAP7_75t_SL u0_g62057 (.A1(u0_n_32839),
    .A2(u0_n_33150),
    .B1(key[46]),
    .B2(u0_n_32942),
    .Y(u0_n_29382));
 AOI22xp33_ASAP7_75t_L u0_g62058 (.A1(u0_n_32875),
    .A2(u0_n_29579),
    .B1(key[42]),
    .B2(u0_n_32942),
    .Y(u0_n_29383));
 AOI22xp33_ASAP7_75t_R u0_g62059 (.A1(u0_n_32924),
    .A2(u0_n_29584),
    .B1(key[86]),
    .B2(u0_n_32942),
    .Y(u0_n_29384));
 AOI22xp33_ASAP7_75t_R u0_g62060 (.A1(u0_n_32924),
    .A2(u0_n_29587),
    .B1(key[83]),
    .B2(u0_n_32942),
    .Y(u0_n_29385));
 AOI22xp5_ASAP7_75t_SL u0_g62061 (.A1(u0_n_32966),
    .A2(u0_n_29582),
    .B1(key[78]),
    .B2(u0_n_32843),
    .Y(u0_n_29386));
 AOI22xp33_ASAP7_75t_R u0_g62062 (.A1(u0_n_32967),
    .A2(u0_n_29571),
    .B1(key[69]),
    .B2(u0_n_32843),
    .Y(u0_n_29387));
 AOI22xp33_ASAP7_75t_R u0_g62063 (.A1(u0_n_32967),
    .A2(u0_n_29574),
    .B1(key[67]),
    .B2(u0_n_32934),
    .Y(u0_n_29388));
 NOR2xp67_ASAP7_75t_SL u0_g62064 (.A(u0_n_32851),
    .B(u0_n_29477),
    .Y(u0_n_29372));
 INVxp33_ASAP7_75t_R u0_g62081 (.A(u0_n_29394),
    .Y(u0_n_29393));
 INVx1_ASAP7_75t_SL u0_g62082 (.A(u0_n_29397),
    .Y(u0_n_29396));
 AOI22xp33_ASAP7_75t_R u0_g62083 (.A1(u0_n_32875),
    .A2(u0_n_29560),
    .B1(key[85]),
    .B2(u0_n_32825),
    .Y(u0_n_29398));
 AOI22xp33_ASAP7_75t_R u0_g62084 (.A1(u0_n_32967),
    .A2(u0_n_29566),
    .B1(key[91]),
    .B2(u0_n_32825),
    .Y(u0_n_29399));
 AOI22xp33_ASAP7_75t_R u0_g62085 (.A1(u0_n_32966),
    .A2(u0_n_29563),
    .B1(key[93]),
    .B2(u0_n_32990),
    .Y(u0_n_29400));
 AOI22xp33_ASAP7_75t_R u0_g62086 (.A1(u0_n_32877),
    .A2(u0_n_29564),
    .B1(key[95]),
    .B2(u0_n_32851),
    .Y(u0_n_29402));
 AOI22xp33_ASAP7_75t_R u0_g62087 (.A1(u0_n_32983),
    .A2(u0_n_29548),
    .B1(key[35]),
    .B2(u0_n_32825),
    .Y(u0_n_29403));
 AOI22xp33_ASAP7_75t_R u0_g62088 (.A1(u0_n_32877),
    .A2(u0_n_29549),
    .B1(key[37]),
    .B2(u0_n_32991),
    .Y(u0_n_29404));
 AOI22xp33_ASAP7_75t_L u0_g62089 (.A1(u0_n_32983),
    .A2(u0_n_29553),
    .B1(key[49]),
    .B2(u0_n_32851),
    .Y(u0_n_29406));
 AOI22xp33_ASAP7_75t_R u0_g62090 (.A1(u0_n_32966),
    .A2(u0_n_29555),
    .B1(key[51]),
    .B2(u0_n_32934),
    .Y(u0_n_29407));
 AOI22xp33_ASAP7_75t_R u0_g62091 (.A1(u0_n_32983),
    .A2(u0_n_29557),
    .B1(key[54]),
    .B2(u0_n_32991),
    .Y(u0_n_29408));
 AOI22xp33_ASAP7_75t_SL u0_g62092 (.A1(u0_n_32877),
    .A2(u0_n_29558),
    .B1(key[57]),
    .B2(u0_n_32851),
    .Y(u0_n_29409));
 XNOR2xp5_ASAP7_75t_L u0_g62093 (.A(u0_n_29565),
    .B(u0_n_31717),
    .Y(u0_n_29410));
 XNOR2xp5_ASAP7_75t_SL u0_g62094 (.A(u0_n_29557),
    .B(u0_n_33004),
    .Y(u0_n_29411));
 XOR2xp5_ASAP7_75t_SL u0_g62095 (.A(u0_n_29561),
    .B(w2[11]),
    .Y(u0_n_29414));
 AOI22xp33_ASAP7_75t_R u0_g62096 (.A1(u0_n_32879),
    .A2(u0_n_29568),
    .B1(key[82]),
    .B2(u0_n_32851),
    .Y(u0_n_29417));
 XOR2xp5_ASAP7_75t_SL u0_g62097 (.A(u0_n_29568),
    .B(w2[18]),
    .Y(u0_n_29418));
 XOR2xp5_ASAP7_75t_SL u0_g62098 (.A(u0_n_29566),
    .B(w2[27]),
    .Y(u0_n_29421));
 XOR2xp5_ASAP7_75t_L u0_g62099 (.A(u0_n_29563),
    .B(w2[29]),
    .Y(u0_n_29424));
 XOR2xp5_ASAP7_75t_SL u0_g62100 (.A(u0_n_29564),
    .B(w2[31]),
    .Y(u0_n_29426));
 XOR2xp5_ASAP7_75t_SL u0_g62101 (.A(u0_n_29554),
    .B(w3[17]),
    .Y(u0_n_29429));
 XNOR2xp5_ASAP7_75t_L u0_g62102 (.A(u0_n_29569),
    .B(u0_n_31721),
    .Y(u0_n_29431));
 XOR2xp5_ASAP7_75t_SL u0_g62103 (.A(u0_n_29559),
    .B(u0_n_32704),
    .Y(u0_n_29432));
 XNOR2xp5_ASAP7_75t_L u0_g62104 (.A(u0_n_29567),
    .B(u0_n_31723),
    .Y(u0_n_29434));
 XOR2xp5_ASAP7_75t_SL u0_g62105 (.A(u0_n_29590),
    .B(u0_n_31693),
    .Y(u0_n_29435));
 OAI22xp5_ASAP7_75t_SL u0_g62106 (.A1(u0_n_32675),
    .A2(u0_n_29522),
    .B1(w1[26]),
    .B2(u0_n_29521),
    .Y(u0_n_29436));
 OAI22xp5_ASAP7_75t_SL u0_g62107 (.A1(u0_n_31571),
    .A2(u0_n_29522),
    .B1(u0_n_31572),
    .B2(u0_n_29521),
    .Y(u0_n_29440));
 XNOR2xp5_ASAP7_75t_SL u0_g62108 (.A(u0_n_29548),
    .B(w3[3]),
    .Y(u0_n_29441));
 AOI22xp33_ASAP7_75t_L u0_g62109 (.A1(n_8668),
    .A2(u0_n_29556),
    .B1(n_8656),
    .B2(u0_n_29555),
    .Y(u0_n_29444));
 XNOR2xp5_ASAP7_75t_SL u0_g62110 (.A(w2[16]),
    .B(u0_n_29551),
    .Y(u0_n_29390));
 XOR2xp5_ASAP7_75t_SL u0_g62111 (.A(w2[8]),
    .B(u0_n_29562),
    .Y(u0_n_29391));
 XOR2xp5_ASAP7_75t_SL u0_g62112 (.A(u0_n_32528),
    .B(u0_n_29560),
    .Y(u0_n_29392));
 XNOR2xp5_ASAP7_75t_SL u0_g62113 (.A(w2[13]),
    .B(u0_n_29552),
    .Y(u0_n_29394));
 XOR2xp5_ASAP7_75t_SL u0_g62114 (.A(w2[0]),
    .B(u0_n_29547),
    .Y(u0_n_29395));
 XNOR2xp5_ASAP7_75t_SL u0_g62115 (.A(w1[24]),
    .B(u0_n_29520),
    .Y(u0_n_29397));
 AOI22xp33_ASAP7_75t_R u0_g62116 (.A1(u0_n_32966),
    .A2(u0_n_29621),
    .B1(key[105]),
    .B2(u0_n_32942),
    .Y(u0_n_29459));
 AOI22xp33_ASAP7_75t_R u0_g62117 (.A1(u0_n_32967),
    .A2(u0_n_29646),
    .B1(key[87]),
    .B2(u0_n_32942),
    .Y(u0_n_29460));
 AOI22xp33_ASAP7_75t_R u0_g62118 (.A1(u0_n_32924),
    .A2(u0_n_29643),
    .B1(key[97]),
    .B2(u0_n_32942),
    .Y(u0_n_29461));
 AOI22xp33_ASAP7_75t_R u0_g62119 (.A1(u0_n_32924),
    .A2(u0_n_29625),
    .B1(key[108]),
    .B2(u0_n_32934),
    .Y(u0_n_29462));
 NAND2xp33_ASAP7_75t_L u0_g62120 (.A(u0_n_29563),
    .B(u0_n_31574),
    .Y(u0_n_29463));
 NAND2xp33_ASAP7_75t_SL u0_g62121 (.A(u0_n_30904),
    .B(u0_n_29521),
    .Y(u0_n_29465));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62122 (.A1(u0_n_30906),
    .A2(u0_n_29661),
    .B(u0_n_29627),
    .C(u0_n_32851),
    .Y(u0_n_29467));
 INVxp33_ASAP7_75t_L u0_g62143 (.A(u0_n_29470),
    .Y(u0_n_29469));
 INVxp67_ASAP7_75t_L u0_g62144 (.A(u0_n_29474),
    .Y(u0_n_29473));
 INVxp33_ASAP7_75t_SL u0_g62145 (.A(u0_n_29476),
    .Y(u0_n_29475));
 INVxp67_ASAP7_75t_SL u0_g62146 (.A(u0_n_29479),
    .Y(u0_n_29478));
 INVxp67_ASAP7_75t_L u0_g62147 (.A(u0_n_29481),
    .Y(u0_n_29482));
 AOI22xp33_ASAP7_75t_R u0_g62148 (.A1(u0_n_32879),
    .A2(u0_n_29619),
    .B1(key[124]),
    .B2(u0_n_32990),
    .Y(u0_n_29483));
 AOI22xp33_ASAP7_75t_R u0_g62149 (.A1(u0_n_32879),
    .A2(u0_n_29617),
    .B1(key[98]),
    .B2(u0_n_32825),
    .Y(u0_n_29484));
 AOI22xp33_ASAP7_75t_R u0_g62150 (.A1(u0_n_32971),
    .A2(u0_n_29616),
    .B1(key[100]),
    .B2(u0_n_32825),
    .Y(u0_n_29485));
 AOI22xp33_ASAP7_75t_R u0_g62151 (.A1(u0_n_32966),
    .A2(u0_n_29620),
    .B1(key[65]),
    .B2(u0_n_32942),
    .Y(u0_n_29486));
 AOI22xp33_ASAP7_75t_R u0_g62152 (.A1(u0_n_32966),
    .A2(u0_n_29635),
    .B1(key[73]),
    .B2(u0_n_32990),
    .Y(u0_n_29487));
 AOI22xp33_ASAP7_75t_R u0_g62153 (.A1(u0_n_32967),
    .A2(u0_n_29632),
    .B1(key[76]),
    .B2(u0_n_32834),
    .Y(u0_n_29488));
 AOI22xp33_ASAP7_75t_R u0_g62154 (.A1(u0_n_32924),
    .A2(u0_n_29639),
    .B1(key[111]),
    .B2(u0_n_32843),
    .Y(u0_n_29489));
 AOI22xp33_ASAP7_75t_R u0_g62155 (.A1(u0_n_32967),
    .A2(u0_n_29642),
    .B1(key[84]),
    .B2(u0_n_32990),
    .Y(u0_n_29490));
 AOI22xp33_ASAP7_75t_R u0_g62156 (.A1(u0_n_32924),
    .A2(u0_n_29637),
    .B1(key[102]),
    .B2(u0_n_32942),
    .Y(u0_n_29491));
 AOI22xp33_ASAP7_75t_SL u0_g62157 (.A1(u0_n_32875),
    .A2(u0_n_29633),
    .B1(key[55]),
    .B2(u0_n_32825),
    .Y(u0_n_29492));
 AOI22xp33_ASAP7_75t_R u0_g62158 (.A1(u0_n_32971),
    .A2(u0_n_29641),
    .B1(key[103]),
    .B2(u0_n_32825),
    .Y(u0_n_29493));
 XOR2xp5_ASAP7_75t_SL u0_g62159 (.A(u0_n_29634),
    .B(n_8831),
    .Y(u0_n_29494));
 XNOR2xp5_ASAP7_75t_SL u0_g62160 (.A(u0_n_29642),
    .B(u0_n_31726),
    .Y(u0_n_29496));
 XOR2xp5_ASAP7_75t_SL u0_g62161 (.A(u0_n_29642),
    .B(w2[20]),
    .Y(u0_n_29498));
 XOR2xp5_ASAP7_75t_SL u0_g62162 (.A(u0_n_29637),
    .B(w1[6]),
    .Y(u0_n_29500));
 XOR2xp5_ASAP7_75t_R u0_g62163 (.A(u0_n_29641),
    .B(w1[7]),
    .Y(u0_n_29503));
 XOR2xp5_ASAP7_75t_L u0_g62164 (.A(u0_n_29640),
    .B(u0_n_31740),
    .Y(u0_n_29506));
 XOR2xp5_ASAP7_75t_SL u0_g62165 (.A(u0_n_31700),
    .B(u0_n_29638),
    .Y(u0_n_29468));
 XNOR2x1_ASAP7_75t_SL u0_g62166 (.B(u0_n_29641),
    .Y(u0_n_29470),
    .A(u0_n_31702));
 XNOR2xp5_ASAP7_75t_SL u0_g62167 (.A(u0_n_29636),
    .B(w2[9]),
    .Y(u0_n_29471));
 XOR2xp5_ASAP7_75t_SL u0_g62168 (.A(u0_n_29632),
    .B(w2[12]),
    .Y(u0_n_29472));
 XNOR2x1_ASAP7_75t_SL u0_g62169 (.B(u0_n_29620),
    .Y(u0_n_29474),
    .A(w2[1]));
 XNOR2xp5_ASAP7_75t_SL u0_g62170 (.A(u0_n_29639),
    .B(w1[15]),
    .Y(u0_n_29476));
 XNOR2xp5_ASAP7_75t_SL u0_g62171 (.A(w1[28]),
    .B(u0_n_29619),
    .Y(u0_n_29477));
 XNOR2x1_ASAP7_75t_SL u0_g62172 (.B(u0_n_29616),
    .Y(u0_n_29479),
    .A(w1[4]));
 XNOR2x1_ASAP7_75t_SL u0_g62173 (.B(u0_n_29618),
    .Y(u0_n_29480),
    .A(w1[2]));
 XNOR2x1_ASAP7_75t_SL u0_g62174 (.B(u0_n_29649),
    .Y(u0_n_29481),
    .A(w0[30]));
 INVxp67_ASAP7_75t_SL u0_g62175 (.A(u0_n_29521),
    .Y(u0_n_29522));
 AOI22xp33_ASAP7_75t_R u0_g62176 (.A1(u0_n_32924),
    .A2(u0_n_29682),
    .B1(key[101]),
    .B2(u0_n_32934),
    .Y(u0_n_29523));
 XNOR2xp5_ASAP7_75t_L u0_g62177 (.A(u0_n_29688),
    .B(w0[25]),
    .Y(u0_n_29524));
 AOI22xp33_ASAP7_75t_R u0_g62178 (.A1(u0_n_32924),
    .A2(u0_n_29684),
    .B1(key[113]),
    .B2(u0_n_32934),
    .Y(u0_n_29526));
 AOI22xp33_ASAP7_75t_R u0_g62179 (.A1(u0_n_32983),
    .A2(u0_n_29663),
    .B1(key[114]),
    .B2(u0_n_32990),
    .Y(u0_n_29527));
 AOI22xp33_ASAP7_75t_R u0_g62180 (.A1(u0_n_32877),
    .A2(u0_n_29657),
    .B1(key[104]),
    .B2(u0_n_33110),
    .Y(u0_n_29528));
 AOI22xp33_ASAP7_75t_R u0_g62181 (.A1(u0_n_32983),
    .A2(u0_n_29679),
    .B1(key[115]),
    .B2(u0_n_32851),
    .Y(u0_n_29529));
 AOI22xp33_ASAP7_75t_R u0_g62182 (.A1(u0_n_32983),
    .A2(u0_n_29659),
    .B1(key[117]),
    .B2(u0_n_32990),
    .Y(u0_n_29530));
 AOI22xp33_ASAP7_75t_R u0_g62183 (.A1(u0_n_32877),
    .A2(u0_n_29678),
    .B1(key[118]),
    .B2(u0_n_32851),
    .Y(u0_n_29531));
 AOI22xp33_ASAP7_75t_R u0_g62184 (.A1(u0_n_32877),
    .A2(u0_n_29683),
    .B1(key[99]),
    .B2(u0_n_33110),
    .Y(u0_n_29532));
 AOI22xp33_ASAP7_75t_L u0_g62185 (.A1(u0_n_32983),
    .A2(u0_n_29660),
    .B1(key[106]),
    .B2(u0_n_32990),
    .Y(u0_n_29533));
 AOI22xp33_ASAP7_75t_R u0_g62186 (.A1(u0_n_32971),
    .A2(u0_n_29680),
    .B1(key[107]),
    .B2(u0_n_32990),
    .Y(u0_n_29534));
 AOI22xp33_ASAP7_75t_R u0_g62187 (.A1(u0_n_32924),
    .A2(u0_n_29662),
    .B1(key[123]),
    .B2(u0_n_32825),
    .Y(u0_n_29535));
 AOI22xp33_ASAP7_75t_R u0_g62188 (.A1(u0_n_32924),
    .A2(u0_n_29676),
    .B1(key[112]),
    .B2(u0_n_32942),
    .Y(u0_n_29536));
 AOI22xp33_ASAP7_75t_R u0_g62189 (.A1(u0_n_32879),
    .A2(u0_n_29668),
    .B1(key[125]),
    .B2(u0_n_32934),
    .Y(u0_n_29537));
 AOI22xp33_ASAP7_75t_R u0_g62190 (.A1(u0_n_32879),
    .A2(u0_n_29677),
    .B1(key[109]),
    .B2(u0_n_32825),
    .Y(u0_n_29538));
 AOI22xp33_ASAP7_75t_R u0_g62191 (.A1(u0_n_32879),
    .A2(u0_n_29681),
    .B1(key[110]),
    .B2(u0_n_32851),
    .Y(u0_n_29539));
 AOI22xp33_ASAP7_75t_R u0_g62192 (.A1(u0_n_32967),
    .A2(u0_n_29664),
    .B1(key[127]),
    .B2(u0_n_32934),
    .Y(u0_n_29540));
 AOI22xp33_ASAP7_75t_R u0_g62193 (.A1(u0_n_32966),
    .A2(u0_n_29665),
    .B1(key[74]),
    .B2(u0_n_32934),
    .Y(u0_n_29541));
 AOI22xp33_ASAP7_75t_R u0_g62194 (.A1(u0_n_32879),
    .A2(u0_n_29666),
    .B1(key[81]),
    .B2(u0_n_32825),
    .Y(u0_n_29542));
 AOI22xp33_ASAP7_75t_R u0_g62195 (.A1(u0_n_32966),
    .A2(u0_n_29667),
    .B1(key[89]),
    .B2(u0_n_32825),
    .Y(u0_n_29543));
 AOI22xp33_ASAP7_75t_R u0_g62196 (.A1(u0_n_32875),
    .A2(u0_n_29658),
    .B1(key[96]),
    .B2(u0_n_32851),
    .Y(u0_n_29544));
 XOR2xp5_ASAP7_75t_SL u0_g62198 (.A(u0_n_29690),
    .B(w0[24]),
    .Y(u0_n_29520));
 XNOR2xp5_ASAP7_75t_SL u0_g62200 (.A(w0[26]),
    .B(u0_n_29687),
    .Y(u0_n_29521));
 INVx1_ASAP7_75t_L u0_g62201 (.A(u0_n_29550),
    .Y(u0_n_29549));
 INVxp67_ASAP7_75t_R u0_g62202 (.A(u0_n_29554),
    .Y(u0_n_29553));
 INVx1_ASAP7_75t_SL u0_g62203 (.A(u0_n_29556),
    .Y(u0_n_29555));
 INVxp67_ASAP7_75t_R u0_g62204 (.A(u0_n_29559),
    .Y(u0_n_29558));
 INVx1_ASAP7_75t_SL u0_g62205 (.A(u0_n_29565),
    .Y(u0_n_29564));
 INVx1_ASAP7_75t_SL u0_g62206 (.A(u0_n_29567),
    .Y(u0_n_29566));
 INVxp67_ASAP7_75t_SL u0_g62207 (.A(u0_n_29569),
    .Y(u0_n_29568));
 XNOR2xp5_ASAP7_75t_SL u0_g62208 (.A(u0_n_29669),
    .B(u0_n_31642),
    .Y(u0_n_29570));
 XOR2xp5_ASAP7_75t_R u0_g62209 (.A(u0_n_29682),
    .B(w1[5]),
    .Y(u0_n_29571));
 XOR2xp5_ASAP7_75t_R u0_g62210 (.A(u0_n_29683),
    .B(w1[3]),
    .Y(u0_n_29574));
 XOR2xp5_ASAP7_75t_L u0_g62212 (.A(u0_n_29665),
    .B(w2[10]),
    .Y(u0_n_29579));
 XOR2xp5_ASAP7_75t_SL u0_g62213 (.A(u0_n_29681),
    .B(w1[14]),
    .Y(u0_n_29582));
 XOR2xp5_ASAP7_75t_R u0_g62214 (.A(u0_n_29678),
    .B(w1[22]),
    .Y(u0_n_29584));
 XOR2xp5_ASAP7_75t_R u0_g62215 (.A(u0_n_29679),
    .B(w1[19]),
    .Y(u0_n_29587));
 XNOR2xp5_ASAP7_75t_L u0_g62216 (.A(u0_n_29680),
    .B(w3[11]),
    .Y(u0_n_29590));
 XOR2xp5_ASAP7_75t_SL u0_g62217 (.A(w1[0]),
    .B(u0_n_29658),
    .Y(u0_n_29547));
 XNOR2x1_ASAP7_75t_SL u0_g62218 (.B(u0_n_29683),
    .Y(u0_n_29548),
    .A(u0_n_31734));
 XNOR2xp5_ASAP7_75t_SL u0_g62219 (.A(u0_n_29682),
    .B(u0_n_31738),
    .Y(u0_n_29550));
 XOR2xp5_ASAP7_75t_SL u0_g62220 (.A(u0_n_29676),
    .B(w1[16]),
    .Y(u0_n_29551));
 XOR2xp5_ASAP7_75t_SL u0_g62221 (.A(w1[13]),
    .B(u0_n_29677),
    .Y(u0_n_29552));
 XNOR2xp5_ASAP7_75t_SL u0_g62222 (.A(w2[17]),
    .B(u0_n_29666),
    .Y(u0_n_29554));
 XOR2xp5_ASAP7_75t_SL u0_g62223 (.A(u0_n_29679),
    .B(u0_n_31698),
    .Y(u0_n_29556));
 XOR2xp5_ASAP7_75t_SL u0_g62224 (.A(u0_n_31704),
    .B(u0_n_29678),
    .Y(u0_n_29557));
 XNOR2xp5_ASAP7_75t_SL u0_g62225 (.A(w2[25]),
    .B(u0_n_29667),
    .Y(u0_n_29559));
 XOR2xp5_ASAP7_75t_SL u0_g62226 (.A(u0_n_29659),
    .B(w1[21]),
    .Y(u0_n_29560));
 XOR2xp5_ASAP7_75t_SL u0_g62227 (.A(w1[11]),
    .B(u0_n_29680),
    .Y(u0_n_29561));
 XOR2xp5_ASAP7_75t_SL u0_g62228 (.A(w1[8]),
    .B(u0_n_29657),
    .Y(u0_n_29562));
 XOR2x2_ASAP7_75t_SL u0_g62229 (.A(u0_n_29668),
    .B(w1[29]),
    .Y(u0_n_29563));
 XNOR2xp5_ASAP7_75t_SL u0_g62230 (.A(u0_n_29664),
    .B(w1[31]),
    .Y(u0_n_29565));
 XNOR2xp5_ASAP7_75t_SL u0_g62231 (.A(w1[27]),
    .B(u0_n_29662),
    .Y(u0_n_29567));
 XNOR2xp5_ASAP7_75t_SL u0_g62232 (.A(w1[18]),
    .B(u0_n_29663),
    .Y(u0_n_29569));
 INVxp33_ASAP7_75t_R u0_g62233 (.A(u0_n_29618),
    .Y(u0_n_29617));
 XNOR2xp5_ASAP7_75t_R u0_g62234 (.A(u0_n_29701),
    .B(w0[9]),
    .Y(u0_n_29621));
 AOI22xp33_ASAP7_75t_R u0_g62235 (.A1(u0_n_32971),
    .A2(u0_n_29709),
    .B1(key[119]),
    .B2(u0_n_32834),
    .Y(u0_n_29623));
 AOI22xp33_ASAP7_75t_R u0_g62236 (.A1(u0_n_32967),
    .A2(u0_n_29708),
    .B1(key[116]),
    .B2(u0_n_32934),
    .Y(u0_n_29624));
 XNOR2xp5_ASAP7_75t_R u0_g62237 (.A(u0_n_29702),
    .B(w0[12]),
    .Y(u0_n_29625));
 NAND2xp5_ASAP7_75t_L u0_g62238 (.A(u0_n_30906),
    .B(u0_n_29661),
    .Y(u0_n_29627));
 XNOR2xp5_ASAP7_75t_SL u0_g62239 (.A(w0[4]),
    .B(u0_n_29706),
    .Y(u0_n_29616));
 XOR2xp5_ASAP7_75t_SL u0_g62240 (.A(u0_n_29704),
    .B(w0[2]),
    .Y(u0_n_29618));
 XOR2xp5_ASAP7_75t_SL u0_g62241 (.A(u0_n_29712),
    .B(u0_n_29763),
    .Y(u0_n_29619));
 XOR2xp5_ASAP7_75t_SL u0_g62242 (.A(u0_n_29700),
    .B(u0_n_31707),
    .Y(u0_n_29620));
 INVxp33_ASAP7_75t_SL u0_g62243 (.A(u0_n_29634),
    .Y(u0_n_29633));
 INVxp33_ASAP7_75t_R u0_g62244 (.A(u0_n_29636),
    .Y(u0_n_29635));
 INVxp67_ASAP7_75t_L u0_g62245 (.A(u0_n_29638),
    .Y(u0_n_29637));
 INVxp67_ASAP7_75t_L u0_g62246 (.A(u0_n_29639),
    .Y(u0_n_29640));
 XOR2xp5_ASAP7_75t_R u0_g62247 (.A(u0_n_29700),
    .B(w0[1]),
    .Y(u0_n_29643));
 XOR2xp5_ASAP7_75t_L u0_g62248 (.A(u0_n_29709),
    .B(w1[23]),
    .Y(u0_n_29646));
 XOR2xp5_ASAP7_75t_SL u0_g62249 (.A(u0_rcon[30]),
    .B(u0_n_29710),
    .Y(u0_n_29649));
 XNOR2xp5_ASAP7_75t_SL u0_g62250 (.A(u0_n_29702),
    .B(u0_n_31696),
    .Y(u0_n_29632));
 XNOR2xp5_ASAP7_75t_SL u0_g62251 (.A(u0_n_29709),
    .B(u0_n_31736),
    .Y(u0_n_29634));
 XOR2xp5_ASAP7_75t_SL u0_g62252 (.A(u0_n_29701),
    .B(u0_n_31694),
    .Y(u0_n_29636));
 XNOR2xp5_ASAP7_75t_SL u0_g62253 (.A(w0[6]),
    .B(u0_n_29711),
    .Y(u0_n_29638));
 XOR2x2_ASAP7_75t_SL u0_g62254 (.A(w0[15]),
    .B(u0_n_29703),
    .Y(u0_n_29639));
 XNOR2x1_ASAP7_75t_SL u0_g62255 (.B(u0_n_29714),
    .Y(u0_n_29641),
    .A(w0[7]));
 XOR2x2_ASAP7_75t_SL u0_g62256 (.A(u0_n_29708),
    .B(w1[20]),
    .Y(u0_n_29642));
 INVxp33_ASAP7_75t_R u0_g62257 (.A(u0_n_29661),
    .Y(u0_n_29660));
 XNOR2xp5_ASAP7_75t_SL u0_g62258 (.A(u0_n_29728),
    .B(u0_n_31729),
    .Y(u0_n_29669));
 XOR2xp5_ASAP7_75t_SL u0_g62259 (.A(w0[8]),
    .B(u0_n_29726),
    .Y(u0_n_29657));
 XNOR2xp5_ASAP7_75t_SL u0_g62260 (.A(w0[0]),
    .B(u0_n_29721),
    .Y(u0_n_29658));
 XNOR2xp5_ASAP7_75t_SL u0_g62261 (.A(u0_n_29731),
    .B(w0[21]),
    .Y(u0_n_29659));
 XOR2xp5_ASAP7_75t_SL u0_g62262 (.A(u0_n_29718),
    .B(w0[10]),
    .Y(u0_n_29661));
 XOR2xp5_ASAP7_75t_SL u0_g62263 (.A(u0_n_29761),
    .B(u0_n_29724),
    .Y(u0_n_29662));
 XNOR2xp5_ASAP7_75t_SL u0_g62264 (.A(w0[18]),
    .B(u0_n_29734),
    .Y(u0_n_29663));
 XOR2xp5_ASAP7_75t_SL u0_g62265 (.A(u0_n_29720),
    .B(u0_n_29813),
    .Y(u0_n_29664));
 XNOR2xp5_ASAP7_75t_L u0_g62266 (.A(u0_n_29718),
    .B(u0_n_31706),
    .Y(u0_n_29665));
 XOR2xp5_ASAP7_75t_SL u0_g62267 (.A(u0_n_29717),
    .B(u0_n_31718),
    .Y(u0_n_29666));
 XOR2xp5_ASAP7_75t_SL u0_g62268 (.A(u0_n_29727),
    .B(u0_n_29815),
    .Y(u0_n_29667));
 XNOR2xp5_ASAP7_75t_SL u0_g62269 (.A(u0_n_29765),
    .B(u0_n_29730),
    .Y(u0_n_29668));
 XOR2xp5_ASAP7_75t_R u0_g62270 (.A(u0_n_29717),
    .B(w0[17]),
    .Y(u0_n_29684));
 XOR2xp5_ASAP7_75t_SL u0_g62271 (.A(u0_n_29722),
    .B(u0_rcon[26]),
    .Y(u0_n_29687));
 XNOR2xp5_ASAP7_75t_L u0_g62272 (.A(u0_n_29727),
    .B(u0_rcon[25]),
    .Y(u0_n_29688));
 XOR2xp5_ASAP7_75t_SL u0_g62273 (.A(u0_n_29725),
    .B(u0_rcon[24]),
    .Y(u0_n_29690));
 XOR2xp5_ASAP7_75t_SL u0_g62274 (.A(u0_n_29719),
    .B(w0[16]),
    .Y(u0_n_29676));
 XOR2xp5_ASAP7_75t_SL u0_g62275 (.A(w0[13]),
    .B(u0_n_29739),
    .Y(u0_n_29677));
 XOR2x2_ASAP7_75t_SL u0_g62276 (.A(w0[22]),
    .B(u0_n_29723),
    .Y(u0_n_29678));
 XNOR2x2_ASAP7_75t_SL u0_g62277 (.A(w0[19]),
    .B(u0_n_29738),
    .Y(u0_n_29679));
 XOR2xp5_ASAP7_75t_SL u0_g62278 (.A(w0[11]),
    .B(u0_n_29733),
    .Y(u0_n_29680));
 XOR2x2_ASAP7_75t_SL u0_g62279 (.A(w0[14]),
    .B(u0_n_29728),
    .Y(u0_n_29681));
 XOR2x2_ASAP7_75t_SL u0_g62280 (.A(u0_n_29735),
    .B(w0[5]),
    .Y(u0_n_29682));
 XOR2x2_ASAP7_75t_SL u0_g62281 (.A(u0_n_29736),
    .B(w0[3]),
    .Y(u0_n_29683));
 AOI211xp5_ASAP7_75t_SL u0_g62282 (.A1(u0_n_29806),
    .A2(w3[5]),
    .B(u0_n_29742),
    .C(u0_n_30255),
    .Y(u0_n_29703));
 AOI221x1_ASAP7_75t_SL u0_g62283 (.A1(u0_n_29804),
    .A2(u0_n_32689),
    .B1(w3[29]),
    .B2(u0_n_29777),
    .C(u0_n_30009),
    .Y(u0_n_29704));
 AOI21xp5_ASAP7_75t_SL u0_g62284 (.A1(u0_n_29754),
    .A2(w3[29]),
    .B(u0_n_29828),
    .Y(u0_n_29706));
 NAND4xp25_ASAP7_75t_SL u0_g62285 (.A(u0_n_29729),
    .B(u0_n_29922),
    .C(u0_n_29981),
    .D(u0_n_29896),
    .Y(u0_n_29700));
 AOI221x1_ASAP7_75t_SL u0_g62286 (.A1(w3[5]),
    .A2(u0_n_29785),
    .B1(u0_n_32691),
    .B2(u0_n_29796),
    .C(u0_n_30068),
    .Y(u0_n_29701));
 AOI221x1_ASAP7_75t_SL u0_g62287 (.A1(u0_n_31761),
    .A2(u0_n_29900),
    .B1(w3[5]),
    .B2(u0_n_29746),
    .C(u0_n_29940),
    .Y(u0_n_29702));
 AOI21xp5_ASAP7_75t_SL u0_g62288 (.A1(u0_n_29755),
    .A2(u0_n_32731),
    .B(u0_n_29759),
    .Y(u0_n_29710));
 AOI221xp5_ASAP7_75t_SL u0_g62289 (.A1(u0_n_30180),
    .A2(u0_n_31516),
    .B1(w3[29]),
    .B2(u0_n_29798),
    .C(u0_n_29745),
    .Y(u0_n_29711));
 OAI21xp5_ASAP7_75t_SL u0_g62290 (.A1(u0_n_32731),
    .A2(u0_n_29744),
    .B(u0_n_29811),
    .Y(u0_n_29712));
 NAND4xp25_ASAP7_75t_SL u0_g62291 (.A(u0_n_30214),
    .B(u0_n_30258),
    .C(u0_n_29838),
    .D(u0_n_29748),
    .Y(u0_n_29714));
 XNOR2xp5_ASAP7_75t_SL u0_g62292 (.A(w0[20]),
    .B(u0_n_29752),
    .Y(u0_n_29708));
 XOR2x2_ASAP7_75t_SL u0_g62293 (.A(w0[23]),
    .B(u0_n_29751),
    .Y(u0_n_29709));
 AOI211x1_ASAP7_75t_SL u0_g62294 (.A1(u0_n_30039),
    .A2(u0_n_31447),
    .B(u0_n_29864),
    .C(u0_n_29780),
    .Y(u0_n_29719));
 AOI321xp33_ASAP7_75t_SL u0_g62295 (.A1(u0_n_29987),
    .A2(u0_n_29963),
    .A3(u0_n_31759),
    .B1(u0_n_29787),
    .B2(w3[21]),
    .C(u0_n_30004),
    .Y(u0_n_29720));
 OAI31xp33_ASAP7_75t_SL u0_g62296 (.A1(u0_n_29881),
    .A2(u0_n_30431),
    .A3(u0_n_30428),
    .B(u0_n_29747),
    .Y(u0_n_29721));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62297 (.A1(u0_n_29948),
    .A2(u0_n_29837),
    .B(u0_n_32731),
    .C(u0_n_29808),
    .Y(u0_n_29722));
 AOI21xp5_ASAP7_75t_SL u0_g62298 (.A1(u0_n_29786),
    .A2(w3[13]),
    .B(u0_n_29757),
    .Y(u0_n_29723));
 O2A1O1Ixp5_ASAP7_75t_SL u0_g62299 (.A1(u0_n_30092),
    .A2(u0_n_29958),
    .B(u0_n_32731),
    .C(u0_n_29756),
    .Y(u0_n_29724));
 AOI211x1_ASAP7_75t_SL u0_g62300 (.A1(u0_n_29852),
    .A2(u0_n_31909),
    .B(u0_n_29850),
    .C(u0_n_29773),
    .Y(u0_n_29725));
 NOR4xp25_ASAP7_75t_SL u0_g62301 (.A(u0_n_29822),
    .B(u0_n_29844),
    .C(u0_n_30082),
    .D(u0_n_29887),
    .Y(u0_n_29726));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62302 (.A1(u0_n_30033),
    .A2(u0_n_29825),
    .B(u0_n_32685),
    .C(u0_n_29778),
    .Y(u0_n_29717));
 O2A1O1Ixp5_ASAP7_75t_SL u0_g62303 (.A1(u0_n_29891),
    .A2(u0_n_29857),
    .B(w3[5]),
    .C(u0_n_29790),
    .Y(u0_n_29718));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62304 (.A1(u0_n_31940),
    .A2(u0_n_30370),
    .B(u0_n_29797),
    .C(w3[29]),
    .Y(u0_n_29729));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62305 (.A1(u0_n_29923),
    .A2(u0_n_29872),
    .B(u0_n_32731),
    .C(u0_n_29795),
    .Y(u0_n_29730));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62306 (.A1(u0_n_29874),
    .A2(u0_n_29994),
    .B(u0_n_32685),
    .C(u0_n_29775),
    .Y(u0_n_29731));
 AOI221xp5_ASAP7_75t_SL u0_g62307 (.A1(u0_n_32691),
    .A2(u0_n_29794),
    .B1(u0_n_29935),
    .B2(u0_n_31912),
    .C(u0_n_29866),
    .Y(u0_n_29733));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62308 (.A1(u0_n_29928),
    .A2(u0_n_29835),
    .B(w3[13]),
    .C(u0_n_29750),
    .Y(u0_n_29734));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62309 (.A1(u0_n_29871),
    .A2(u0_n_29933),
    .B(w3[29]),
    .C(u0_n_29776),
    .Y(u0_n_29735));
 AOI21xp5_ASAP7_75t_SL u0_g62310 (.A1(u0_n_29789),
    .A2(u0_n_32689),
    .B(u0_n_29753),
    .Y(u0_n_29736));
 OAI221xp5_ASAP7_75t_SL u0_g62311 (.A1(w3[13]),
    .A2(u0_n_29781),
    .B1(u0_n_29846),
    .B2(u0_n_31914),
    .C(u0_n_29861),
    .Y(u0_n_29738));
 AOI221xp5_ASAP7_75t_SL u0_g62312 (.A1(u0_n_29783),
    .A2(w3[5]),
    .B1(u0_n_30062),
    .B2(u0_n_31514),
    .C(u0_n_29821),
    .Y(u0_n_29739));
 OAI321xp33_ASAP7_75t_SL u0_g62313 (.A1(u0_n_29910),
    .A2(u0_n_32753),
    .A3(w3[21]),
    .B1(u0_n_32731),
    .B2(u0_n_29801),
    .C(u0_n_29903),
    .Y(u0_n_29727));
 AOI221xp5_ASAP7_75t_SL u0_g62314 (.A1(w3[5]),
    .A2(u0_n_29802),
    .B1(u0_n_30146),
    .B2(u0_n_31514),
    .C(u0_n_29774),
    .Y(u0_n_29728));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62315 (.A1(w3[2]),
    .A2(u0_n_30296),
    .B(u0_n_29868),
    .C(u0_n_30138),
    .Y(u0_n_29742));
 AOI221xp5_ASAP7_75t_SL u0_g62316 (.A1(u0_n_32741),
    .A2(u0_n_29908),
    .B1(u0_n_30101),
    .B2(u0_n_31957),
    .C(u0_n_29976),
    .Y(u0_n_29744));
 OAI22xp5_ASAP7_75t_SL u0_g62317 (.A1(u0_n_31768),
    .A2(u0_n_29870),
    .B1(u0_n_31458),
    .B2(u0_n_30443),
    .Y(u0_n_29745));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62318 (.A1(u0_n_30569),
    .A2(u0_n_30357),
    .B(u0_n_31789),
    .C(u0_n_29782),
    .Y(u0_n_29746));
 AOI311xp33_ASAP7_75t_SL u0_g62319 (.A1(u0_n_30099),
    .A2(u0_n_30081),
    .A3(u0_n_31751),
    .B(u0_n_29869),
    .C(u0_n_30096),
    .Y(u0_n_29747));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62320 (.A1(u0_n_31940),
    .A2(u0_n_30235),
    .B(u0_n_29859),
    .C(w3[29]),
    .Y(u0_n_29748));
 OAI211xp5_ASAP7_75t_SL u0_g62321 (.A1(u0_n_31521),
    .A2(u0_n_30018),
    .B(u0_n_29772),
    .C(u0_n_29975),
    .Y(u0_n_29750));
 AOI21xp5_ASAP7_75t_SL u0_g62322 (.A1(u0_n_29855),
    .A2(w3[13]),
    .B(u0_n_29807),
    .Y(u0_n_29751));
 AOI211xp5_ASAP7_75t_SL u0_g62323 (.A1(u0_n_29909),
    .A2(u0_n_31757),
    .B(u0_n_29791),
    .C(u0_n_29863),
    .Y(u0_n_29752));
 OAI221xp5_ASAP7_75t_SL u0_g62324 (.A1(u0_n_29842),
    .A2(u0_n_31910),
    .B1(u0_n_29997),
    .B2(u0_n_31406),
    .C(u0_n_29969),
    .Y(u0_n_29753));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62325 (.A1(u0_n_30565),
    .A2(u0_n_30352),
    .B(u0_n_31797),
    .C(u0_n_29800),
    .Y(u0_n_29754));
 OAI221xp5_ASAP7_75t_SL u0_g62326 (.A1(u0_n_29848),
    .A2(\u0_w[3] [16]),
    .B1(u0_n_30176),
    .B2(u0_n_31787),
    .C(u0_n_30132),
    .Y(u0_n_29755));
 OAI221xp5_ASAP7_75t_SL u0_g62327 (.A1(u0_n_30024),
    .A2(u0_n_31432),
    .B1(u0_n_29992),
    .B2(u0_n_31389),
    .C(u0_n_29770),
    .Y(u0_n_29756));
 OAI221xp5_ASAP7_75t_SL u0_g62328 (.A1(u0_n_30141),
    .A2(u0_n_31521),
    .B1(u0_n_30450),
    .B2(u0_n_31451),
    .C(u0_n_29767),
    .Y(u0_n_29757));
 OAI321xp33_ASAP7_75t_SL u0_g62329 (.A1(u0_n_30266),
    .A2(u0_n_31949),
    .A3(u0_n_32731),
    .B1(u0_n_31432),
    .B2(u0_n_30064),
    .C(u0_n_29810),
    .Y(u0_n_29759));
 XOR2xp5_ASAP7_75t_R u0_g62330 (.A(w0[27]),
    .B(u0_rcon[27]),
    .Y(u0_n_29761));
 XOR2xp5_ASAP7_75t_R u0_g62331 (.A(w0[28]),
    .B(u0_rcon[28]),
    .Y(u0_n_29763));
 XOR2xp5_ASAP7_75t_R u0_g62332 (.A(w0[29]),
    .B(u0_rcon[29]),
    .Y(u0_n_29765));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62333 (.A1(w3[10]),
    .A2(u0_n_30013),
    .B(u0_n_30104),
    .C(u0_n_31757),
    .Y(u0_n_29767));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62334 (.A1(u0_n_30908),
    .A2(u0_n_30182),
    .B(u0_n_29951),
    .C(u0_n_31909),
    .Y(u0_n_29770));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62335 (.A1(u0_n_31444),
    .A2(u0_n_30753),
    .B(u0_n_29957),
    .C(u0_n_31764),
    .Y(u0_n_29772));
 OAI22xp5_ASAP7_75t_SL u0_g62336 (.A1(u0_n_30195),
    .A2(u0_n_29877),
    .B1(u0_n_30054),
    .B2(u0_n_31432),
    .Y(u0_n_29773));
 NAND2xp33_ASAP7_75t_L u0_g62337 (.A(u0_n_30122),
    .B(u0_n_29840),
    .Y(u0_n_29774));
 AOI211xp5_ASAP7_75t_SL u0_g62338 (.A1(u0_n_30123),
    .A2(u0_n_31479),
    .B(u0_n_29912),
    .C(u0_n_29959),
    .Y(u0_n_29775));
 OAI211xp5_ASAP7_75t_SL u0_g62339 (.A1(u0_n_31454),
    .A2(u0_n_30124),
    .B(u0_n_29950),
    .C(u0_n_29913),
    .Y(u0_n_29776));
 NAND4xp25_ASAP7_75t_SL u0_g62340 (.A(u0_n_30044),
    .B(u0_n_29924),
    .C(u0_n_29999),
    .D(u0_n_29973),
    .Y(u0_n_29777));
 AOI221xp5_ASAP7_75t_SL u0_g62341 (.A1(u0_n_30498),
    .A2(u0_n_30419),
    .B1(u0_n_30072),
    .B2(u0_n_31479),
    .C(u0_n_29936),
    .Y(u0_n_29778));
 OAI31xp33_ASAP7_75t_SL u0_g62342 (.A1(u0_n_30080),
    .A2(u0_n_30144),
    .A3(u0_n_31765),
    .B(u0_n_29911),
    .Y(u0_n_29780));
 AOI311xp33_ASAP7_75t_SL u0_g62343 (.A1(u0_n_30358),
    .A2(u0_n_30457),
    .A3(u0_n_30477),
    .B(u0_n_29930),
    .C(u0_n_30078),
    .Y(u0_n_29781));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62344 (.A1(u0_n_30286),
    .A2(u0_n_30021),
    .B(u0_n_32695),
    .C(u0_n_29968),
    .Y(u0_n_29782));
 OAI321xp33_ASAP7_75t_SL u0_g62345 (.A1(u0_n_30353),
    .A2(u0_n_30341),
    .A3(u0_n_30722),
    .B1(u0_n_31789),
    .B2(u0_n_30032),
    .C(u0_n_29934),
    .Y(u0_n_29783));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62346 (.A1(u0_n_30686),
    .A2(u0_n_30367),
    .B(u0_n_31941),
    .C(u0_n_29824),
    .Y(u0_n_29785));
 OAI221xp5_ASAP7_75t_SL u0_g62347 (.A1(u0_n_30031),
    .A2(u0_n_31783),
    .B1(u0_n_30267),
    .B2(u0_n_31932),
    .C(u0_n_29832),
    .Y(u0_n_29786));
 OAI221xp5_ASAP7_75t_SL u0_g62348 (.A1(u0_n_30233),
    .A2(u0_n_31958),
    .B1(u0_n_30108),
    .B2(u0_n_31949),
    .C(u0_n_29819),
    .Y(u0_n_29787));
 OAI211xp5_ASAP7_75t_SL u0_g62349 (.A1(u0_n_30159),
    .A2(u0_n_30350),
    .B(u0_n_29932),
    .C(u0_n_30087),
    .Y(u0_n_29789));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62350 (.A1(u0_n_30178),
    .A2(u0_n_30016),
    .B(u0_n_31755),
    .C(u0_n_29817),
    .Y(u0_n_29790));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62351 (.A1(u0_n_30648),
    .A2(u0_n_30358),
    .B(u0_n_31451),
    .C(u0_n_29818),
    .Y(u0_n_29791));
 OAI211xp5_ASAP7_75t_SL u0_g62352 (.A1(u0_n_30349),
    .A2(u0_n_30161),
    .B(u0_n_29931),
    .C(u0_n_30083),
    .Y(u0_n_29794));
 AOI221x1_ASAP7_75t_SL u0_g62353 (.A1(u0_n_30058),
    .A2(u0_n_30155),
    .B1(u0_n_30059),
    .B2(u0_n_31512),
    .C(u0_n_30223),
    .Y(u0_n_29795));
 OAI21xp5_ASAP7_75t_SL u0_g62354 (.A1(u0_n_32747),
    .A2(u0_n_29894),
    .B(u0_n_30090),
    .Y(u0_n_29796));
 OAI211xp5_ASAP7_75t_SL u0_g62355 (.A1(u0_n_31939),
    .A2(u0_n_30668),
    .B(u0_n_30190),
    .C(u0_n_29853),
    .Y(u0_n_29797));
 OAI211xp5_ASAP7_75t_SL u0_g62356 (.A1(u0_n_31797),
    .A2(u0_n_30035),
    .B(u0_n_29833),
    .C(u0_n_29962),
    .Y(u0_n_29798));
 AOI22xp5_ASAP7_75t_L u0_g62357 (.A1(u0_n_29929),
    .A2(u0_n_32687),
    .B1(u0_n_30204),
    .B2(u0_n_31973),
    .Y(u0_n_29800));
 AOI211xp5_ASAP7_75t_SL u0_g62358 (.A1(u0_n_30273),
    .A2(u0_n_31770),
    .B(u0_n_29983),
    .C(u0_n_29831),
    .Y(u0_n_29801));
 OAI221xp5_ASAP7_75t_SL u0_g62359 (.A1(u0_n_30028),
    .A2(u0_n_31789),
    .B1(u0_n_30263),
    .B2(u0_n_31941),
    .C(u0_n_29826),
    .Y(u0_n_29802));
 OAI22xp5_ASAP7_75t_SL u0_g62360 (.A1(u0_n_29919),
    .A2(w3[26]),
    .B1(u0_n_29889),
    .B2(u0_n_31797),
    .Y(u0_n_29804));
 OAI211xp5_ASAP7_75t_L u0_g62361 (.A1(u0_n_31941),
    .A2(u0_n_30257),
    .B(u0_n_29941),
    .C(u0_n_29938),
    .Y(u0_n_29806));
 NAND3xp33_ASAP7_75t_SL u0_g62362 (.A(u0_n_30201),
    .B(u0_n_29845),
    .C(u0_n_30249),
    .Y(u0_n_29807));
 AOI221xp5_ASAP7_75t_SL u0_g62363 (.A1(u0_n_29944),
    .A2(u0_n_31760),
    .B1(u0_n_30094),
    .B2(u0_n_31512),
    .C(u0_n_30252),
    .Y(u0_n_29808));
 OAI211xp5_ASAP7_75t_SL u0_g62364 (.A1(u0_n_29984),
    .A2(u0_n_29952),
    .B(u0_n_32753),
    .C(w3[21]),
    .Y(u0_n_29810));
 AOI221xp5_ASAP7_75t_SL u0_g62365 (.A1(u0_n_30425),
    .A2(u0_n_31512),
    .B1(u0_n_31759),
    .B2(u0_n_29926),
    .C(u0_n_30001),
    .Y(u0_n_29811));
 XOR2xp5_ASAP7_75t_R u0_g62366 (.A(w0[31]),
    .B(u0_rcon[31]),
    .Y(u0_n_29813));
 XNOR2xp5_ASAP7_75t_R u0_g62367 (.A(u0_n_31730),
    .B(u0_rcon[25]),
    .Y(u0_n_29815));
 AOI21xp5_ASAP7_75t_L u0_g62368 (.A1(u0_n_30056),
    .A2(u0_n_31514),
    .B(u0_n_30250),
    .Y(u0_n_29817));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62369 (.A1(u0_n_30472),
    .A2(u0_n_30115),
    .B(u0_n_30268),
    .C(u0_n_31915),
    .Y(u0_n_29818));
 A2O1A1O1Ixp25_ASAP7_75t_SL u0_g62370 (.A1(u0_n_31650),
    .A2(u0_n_32021),
    .B(u0_n_30644),
    .C(u0_n_31770),
    .D(u0_n_29901),
    .Y(u0_n_29819));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62371 (.A1(u0_n_31443),
    .A2(u0_n_30760),
    .B(u0_n_29970),
    .C(u0_n_30183),
    .Y(u0_n_29821));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62372 (.A1(u0_n_30409),
    .A2(u0_n_30134),
    .B(u0_n_32747),
    .C(u0_n_30126),
    .Y(u0_n_29822));
 AOI221xp5_ASAP7_75t_SL u0_g62373 (.A1(u0_n_30121),
    .A2(u0_n_31779),
    .B1(u0_n_30602),
    .B2(u0_n_31790),
    .C(u0_n_29960),
    .Y(u0_n_29824));
 AOI221xp5_ASAP7_75t_SL u0_g62374 (.A1(u0_n_30120),
    .A2(u0_n_31777),
    .B1(u0_n_30536),
    .B2(u0_n_31784),
    .C(u0_n_29916),
    .Y(u0_n_29825));
 AOI22xp5_ASAP7_75t_L u0_g62375 (.A1(u0_n_31967),
    .A2(u0_n_29964),
    .B1(u0_n_31779),
    .B2(u0_n_30211),
    .Y(u0_n_29826));
 OAI322xp33_ASAP7_75t_SL u0_g62376 (.A1(u0_n_31768),
    .A2(u0_n_30269),
    .A3(u0_n_29989),
    .B1(u0_n_31458),
    .B2(u0_n_30109),
    .C1(u0_n_31517),
    .C2(u0_n_30422),
    .Y(u0_n_29828));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62377 (.A1(u0_n_30597),
    .A2(u0_n_30372),
    .B(u0_n_31949),
    .C(u0_n_29878),
    .Y(u0_n_29831));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62378 (.A1(u0_n_30293),
    .A2(u0_n_30356),
    .B(u0_n_31955),
    .C(u0_n_30006),
    .Y(u0_n_29832));
 AOI22xp33_ASAP7_75t_SL u0_g62379 (.A1(u0_n_31973),
    .A2(u0_n_29966),
    .B1(u0_n_31774),
    .B2(u0_n_30209),
    .Y(u0_n_29833));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62380 (.A1(u0_n_30615),
    .A2(u0_n_30355),
    .B(u0_n_31783),
    .C(u0_n_29883),
    .Y(u0_n_29835));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62381 (.A1(u0_n_30310),
    .A2(u0_n_30371),
    .B(u0_n_31950),
    .C(u0_n_30037),
    .Y(u0_n_29837));
 OAI21xp33_ASAP7_75t_L u0_g62382 (.A1(u0_n_32687),
    .A2(u0_n_30168),
    .B(u0_n_29886),
    .Y(u0_n_29838));
 OAI21xp33_ASAP7_75t_L u0_g62383 (.A1(u0_n_30224),
    .A2(u0_n_30076),
    .B(u0_n_31761),
    .Y(u0_n_29840));
 AOI322xp5_ASAP7_75t_SL u0_g62388 (.A1(u0_n_30504),
    .A2(u0_n_30721),
    .A3(u0_n_30782),
    .B1(u0_n_32743),
    .B2(u0_n_30279),
    .C1(u0_n_31440),
    .C2(n_8942),
    .Y(u0_n_29842));
 OAI321xp33_ASAP7_75t_SL u0_g62389 (.A1(u0_n_30382),
    .A2(u0_n_31292),
    .A3(u0_n_31403),
    .B1(u0_n_30242),
    .B2(u0_n_30864),
    .C(u0_n_30298),
    .Y(u0_n_29844));
 OAI211xp5_ASAP7_75t_L u0_g62390 (.A1(w3[10]),
    .A2(u0_n_30194),
    .B(u0_n_30008),
    .C(u0_n_31757),
    .Y(u0_n_29845));
 AOI221xp5_ASAP7_75t_SL u0_g62391 (.A1(u0_n_30276),
    .A2(u0_n_32745),
    .B1(u0_n_31444),
    .B2(w3[12]),
    .C(u0_n_30321),
    .Y(u0_n_29846));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62392 (.A1(u0_n_30360),
    .A2(u0_n_30217),
    .B(w3[18]),
    .C(u0_n_30136),
    .Y(u0_n_29848));
 OAI331xp33_ASAP7_75t_SL u0_g62393 (.A1(u0_n_30529),
    .A2(u0_n_31308),
    .A3(u0_n_31389),
    .B1(u0_n_30869),
    .B2(u0_n_30629),
    .B3(u0_n_31510),
    .C1(u0_n_30289),
    .Y(u0_n_29850));
 AOI211xp5_ASAP7_75t_SL u0_g62394 (.A1(u0_n_30052),
    .A2(u0_n_32753),
    .B(u0_n_30445),
    .C(u0_n_31006),
    .Y(u0_n_29852));
 AOI322xp5_ASAP7_75t_SL u0_g62395 (.A1(u0_n_31331),
    .A2(u0_n_31774),
    .A3(u0_n_32304),
    .B1(u0_n_31798),
    .B2(u0_n_30544),
    .C1(u0_n_31973),
    .C2(u0_n_30049),
    .Y(u0_n_29853));
 OAI221xp5_ASAP7_75t_SL u0_g62396 (.A1(u0_n_30200),
    .A2(u0_n_31956),
    .B1(u0_n_30247),
    .B2(u0_n_31932),
    .C(u0_n_29937),
    .Y(u0_n_29855));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62397 (.A1(u0_n_30314),
    .A2(u0_n_30367),
    .B(u0_n_31941),
    .C(u0_n_30029),
    .Y(u0_n_29857));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62398 (.A1(u0_n_30721),
    .A2(u0_n_30339),
    .B(u0_n_31974),
    .C(u0_n_29946),
    .Y(u0_n_29859));
 AOI22xp33_ASAP7_75t_SL u0_g62399 (.A1(u0_n_31447),
    .A2(u0_n_30102),
    .B1(u0_n_31412),
    .B2(u0_n_29991),
    .Y(u0_n_29861));
 OAI221xp5_ASAP7_75t_SL u0_g62400 (.A1(u0_n_30423),
    .A2(u0_n_31521),
    .B1(u0_n_30156),
    .B2(u0_n_31411),
    .C(u0_n_29978),
    .Y(u0_n_29863));
 AOI211xp5_ASAP7_75t_SL u0_g62401 (.A1(u0_n_30066),
    .A2(u0_n_32745),
    .B(u0_n_30435),
    .C(u0_n_30578),
    .Y(u0_n_29864));
 OAI22xp5_ASAP7_75t_SL u0_g62402 (.A1(u0_n_31405),
    .A2(u0_n_30014),
    .B1(u0_n_31403),
    .B2(u0_n_29990),
    .Y(u0_n_29866));
 OAI221xp5_ASAP7_75t_SL u0_g62403 (.A1(u0_n_29971),
    .A2(w3[2]),
    .B1(u0_n_31426),
    .B2(u0_n_31583),
    .C(u0_n_31761),
    .Y(u0_n_29868));
 OAI221xp5_ASAP7_75t_SL u0_g62404 (.A1(u0_n_30041),
    .A2(u0_n_31408),
    .B1(u0_n_31311),
    .B2(u0_n_30463),
    .C(u0_n_30270),
    .Y(u0_n_29869));
 AOI22xp33_ASAP7_75t_SL u0_g62405 (.A1(w3[26]),
    .A2(u0_n_30043),
    .B1(u0_n_32687),
    .B2(u0_n_30375),
    .Y(u0_n_29870));
 OAI211xp5_ASAP7_75t_SL u0_g62406 (.A1(u0_n_31797),
    .A2(u0_n_30346),
    .B(u0_n_30003),
    .C(u0_n_30332),
    .Y(u0_n_29871));
 AOI221x1_ASAP7_75t_SL u0_g62407 (.A1(u0_n_33149),
    .A2(u0_n_31788),
    .B1(u0_n_30193),
    .B2(u0_n_31950),
    .C(u0_n_30330),
    .Y(u0_n_29872));
 AOI221xp5_ASAP7_75t_SL u0_g62408 (.A1(u0_n_30051),
    .A2(u0_n_31784),
    .B1(u0_n_30158),
    .B2(u0_n_31933),
    .C(u0_n_30323),
    .Y(u0_n_29874));
 OAI221xp5_ASAP7_75t_L u0_g62409 (.A1(u0_n_31237),
    .A2(u0_n_31468),
    .B1(u0_n_31409),
    .B2(u0_n_31935),
    .C(u0_n_30137),
    .Y(u0_n_29877));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62410 (.A1(u0_n_32021),
    .A2(u0_n_31153),
    .B(u0_n_30148),
    .C(u0_n_31957),
    .Y(u0_n_29878));
 A2O1A1O1Ixp25_ASAP7_75t_SL u0_g62411 (.A1(u0_n_31491),
    .A2(u0_n_31184),
    .B(u0_n_32053),
    .C(u0_n_30218),
    .D(w3[24]),
    .Y(u0_n_29881));
 AOI22xp33_ASAP7_75t_SL u0_g62412 (.A1(u0_n_31955),
    .A2(u0_n_30232),
    .B1(u0_n_31777),
    .B2(u0_n_30237),
    .Y(u0_n_29883));
 AOI21xp5_ASAP7_75t_L u0_g62413 (.A1(u0_n_32687),
    .A2(u0_n_30187),
    .B(u0_n_31768),
    .Y(u0_n_29886));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62414 (.A1(u0_n_32763),
    .A2(u0_n_30570),
    .B(u0_n_30658),
    .C(u0_n_31405),
    .Y(u0_n_29887));
 AOI211xp5_ASAP7_75t_L u0_g62415 (.A1(u0_n_31236),
    .A2(u0_n_32063),
    .B(u0_n_30768),
    .C(u0_n_30324),
    .Y(u0_n_29889));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62416 (.A1(u0_n_30733),
    .A2(u0_n_30373),
    .B(u0_n_30098),
    .C(u0_n_32839),
    .Y(u0_n_29890));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62417 (.A1(u0_n_30766),
    .A2(u0_n_30705),
    .B(u0_n_31968),
    .C(u0_n_29972),
    .Y(u0_n_29891));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62418 (.A1(u0_n_30733),
    .A2(u0_n_30369),
    .B(u0_n_31110),
    .C(u0_n_32835),
    .Y(u0_n_29892));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62419 (.A1(u0_n_31422),
    .A2(u0_n_30353),
    .B(w3[2]),
    .C(u0_n_29988),
    .Y(u0_n_29894));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62420 (.A1(u0_n_32040),
    .A2(u0_n_31148),
    .B(u0_n_30280),
    .C(u0_n_31455),
    .Y(u0_n_29896));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62421 (.A1(u0_n_30734),
    .A2(u0_n_30373),
    .B(u0_n_30506),
    .C(u0_n_32839),
    .Y(u0_n_29898));
 OAI21xp5_ASAP7_75t_L u0_g62422 (.A1(w3[2]),
    .A2(u0_n_30160),
    .B(u0_n_30284),
    .Y(u0_n_29900));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62423 (.A1(u0_n_32795),
    .A2(u0_n_31272),
    .B(u0_n_30165),
    .C(u0_n_31787),
    .Y(u0_n_29901));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62424 (.A1(u0_n_32242),
    .A2(u0_n_31312),
    .B(u0_n_30274),
    .C(u0_n_30070),
    .Y(u0_n_29903));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62425 (.A1(u0_n_30734),
    .A2(u0_n_30369),
    .B(u0_n_30098),
    .C(u0_n_32839),
    .Y(u0_n_29904));
 OAI321xp33_ASAP7_75t_SL u0_g62426 (.A1(u0_n_30963),
    .A2(u0_n_30215),
    .A3(\u0_w[3] [16]),
    .B1(u0_n_31917),
    .B2(u0_n_30910),
    .C(u0_n_30608),
    .Y(u0_n_29908));
 OAI22xp33_ASAP7_75t_L u0_g62427 (.A1(u0_n_30166),
    .A2(w3[10]),
    .B1(u0_n_30240),
    .B2(u0_n_32683),
    .Y(u0_n_29909));
 AOI221xp5_ASAP7_75t_L u0_g62428 (.A1(u0_n_30365),
    .A2(w3[18]),
    .B1(u0_n_30441),
    .B2(u0_n_30715),
    .C(u0_n_30192),
    .Y(u0_n_29910));
 AOI331xp33_ASAP7_75t_SL u0_g62429 (.A1(u0_n_30811),
    .A2(u0_n_31038),
    .A3(u0_n_31299),
    .B1(u0_n_30843),
    .B2(u0_n_30418),
    .B3(u0_n_31520),
    .C1(u0_n_30283),
    .Y(u0_n_29911));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62430 (.A1(u0_n_32185),
    .A2(u0_n_30728),
    .B(u0_n_30302),
    .C(u0_n_31521),
    .Y(u0_n_29912));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62431 (.A1(u0_n_32320),
    .A2(u0_n_30735),
    .B(u0_n_30299),
    .C(u0_n_31516),
    .Y(u0_n_29913));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62432 (.A1(u0_n_32194),
    .A2(u0_n_31120),
    .B(u0_n_30153),
    .C(u0_n_31956),
    .Y(u0_n_29916));
 AOI221xp5_ASAP7_75t_SL u0_g62436 (.A1(u0_n_30594),
    .A2(u0_n_32743),
    .B1(u0_n_30769),
    .B2(u0_n_31440),
    .C(u0_n_30191),
    .Y(u0_n_29919));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62437 (.A1(u0_n_30605),
    .A2(u0_n_30514),
    .B(u0_n_31516),
    .C(u0_n_30185),
    .Y(u0_n_29922));
 OAI211xp5_ASAP7_75t_R u0_g62438 (.A1(u0_n_32209),
    .A2(u0_n_31181),
    .B(u0_n_30343),
    .C(u0_n_30366),
    .Y(u0_n_29923));
 OAI21xp5_ASAP7_75t_L u0_g62439 (.A1(u0_n_30304),
    .A2(u0_n_30370),
    .B(u0_n_31940),
    .Y(u0_n_29924));
 OAI221xp5_ASAP7_75t_SL u0_g62440 (.A1(u0_n_31312),
    .A2(u0_n_31417),
    .B1(u0_n_31553),
    .B2(u0_n_31752),
    .C(u0_n_30011),
    .Y(u0_n_29926));
 AOI21xp5_ASAP7_75t_R u0_g62441 (.A1(u0_n_30368),
    .A2(u0_n_30317),
    .B(u0_n_31932),
    .Y(u0_n_29928));
 OAI321xp33_ASAP7_75t_SL u0_g62442 (.A1(u0_n_30362),
    .A2(u0_n_30899),
    .A3(u0_n_30488),
    .B1(u0_n_31769),
    .B2(u0_n_30903),
    .C(u0_n_30676),
    .Y(u0_n_29929));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62443 (.A1(u0_n_32353),
    .A2(u0_n_31303),
    .B(u0_n_30405),
    .C(u0_n_30020),
    .Y(u0_n_29930));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62444 (.A1(u0_n_31886),
    .A2(u0_n_31266),
    .B(u0_n_30530),
    .C(u0_n_30022),
    .Y(u0_n_29931));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62445 (.A1(u0_n_32290),
    .A2(u0_n_31277),
    .B(u0_n_30395),
    .C(u0_n_30027),
    .Y(u0_n_29932));
 AOI211xp5_ASAP7_75t_R u0_g62446 (.A1(u0_n_31173),
    .A2(u0_n_32040),
    .B(u0_n_30170),
    .C(u0_n_30726),
    .Y(u0_n_29933));
 AOI21xp5_ASAP7_75t_SL u0_g62447 (.A1(u0_n_30196),
    .A2(u0_n_31942),
    .B(u0_n_30334),
    .Y(u0_n_29934));
 OAI32xp33_ASAP7_75t_L u0_g62448 (.A1(u0_n_30404),
    .A2(u0_n_30727),
    .A3(u0_n_30788),
    .B1(n_11482),
    .B2(u0_n_30199),
    .Y(u0_n_29935));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62449 (.A1(u0_n_30589),
    .A2(u0_n_30359),
    .B(u0_n_31521),
    .C(u0_n_30221),
    .Y(u0_n_29936));
 AOI21xp33_ASAP7_75t_L u0_g62450 (.A1(u0_n_30524),
    .A2(u0_n_31777),
    .B(u0_n_30017),
    .Y(u0_n_29937));
 AOI22xp33_ASAP7_75t_R u0_g62451 (.A1(u0_n_31790),
    .A2(u0_n_30229),
    .B1(u0_n_31779),
    .B2(u0_n_30540),
    .Y(u0_n_29938));
 OAI22xp5_ASAP7_75t_L u0_g62452 (.A1(u0_n_31420),
    .A2(u0_n_30111),
    .B1(u0_n_31515),
    .B2(u0_n_30420),
    .Y(u0_n_29940));
 OAI21xp33_ASAP7_75t_R u0_g62453 (.A1(u0_n_30727),
    .A2(u0_n_30326),
    .B(u0_n_31967),
    .Y(u0_n_29941));
 OAI322xp33_ASAP7_75t_SL u0_g62454 (.A1(u0_n_30961),
    .A2(u0_n_31196),
    .A3(u0_n_30469),
    .B1(\u0_w[3] [16]),
    .B2(u0_n_30598),
    .C1(u0_n_30772),
    .C2(u0_n_31409),
    .Y(u0_n_29944));
 AOI22xp5_ASAP7_75t_SL u0_g62455 (.A1(u0_n_31798),
    .A2(u0_n_30197),
    .B1(u0_n_31774),
    .B2(u0_n_30503),
    .Y(u0_n_29946));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62456 (.A1(u0_n_30623),
    .A2(u0_n_30354),
    .B(u0_n_31788),
    .C(u0_n_29980),
    .Y(u0_n_29948));
 OAI221xp5_ASAP7_75t_SL u0_g62457 (.A1(u0_n_30765),
    .A2(u0_n_31438),
    .B1(u0_n_30729),
    .B2(u0_n_30541),
    .C(u0_n_30114),
    .Y(u0_n_29950));
 OAI22xp5_ASAP7_75t_SL u0_g62458 (.A1(\u0_w[3] [16]),
    .A2(u0_n_30277),
    .B1(u0_n_33138),
    .B2(u0_n_31409),
    .Y(u0_n_29951));
 OAI322xp33_ASAP7_75t_SL u0_g62459 (.A1(u0_n_31317),
    .A2(u0_n_32249),
    .A3(u0_n_32741),
    .B1(u0_n_31752),
    .B2(u0_n_30385),
    .C1(u0_n_30771),
    .C2(u0_n_31417),
    .Y(u0_n_29952));
 AOI22xp33_ASAP7_75t_SL u0_g62460 (.A1(n_11401),
    .A2(u0_n_30292),
    .B1(u0_n_32745),
    .B2(u0_n_30704),
    .Y(u0_n_29957));
 OAI221xp5_ASAP7_75t_SL u0_g62461 (.A1(u0_n_30163),
    .A2(u0_n_30351),
    .B1(u0_n_30659),
    .B2(u0_n_30491),
    .C(u0_n_30207),
    .Y(u0_n_29958));
 AOI211xp5_ASAP7_75t_SL u0_g62462 (.A1(u0_n_30757),
    .A2(u0_n_31442),
    .B(u0_n_30172),
    .C(u0_n_30244),
    .Y(u0_n_29959));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62463 (.A1(u0_n_31842),
    .A2(u0_n_31161),
    .B(u0_n_30150),
    .C(u0_n_31968),
    .Y(u0_n_29960));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62464 (.A1(u0_n_32052),
    .A2(u0_n_31671),
    .B(u0_n_30582),
    .C(u0_n_31940),
    .Y(u0_n_29962));
 NAND2xp33_ASAP7_75t_R u0_g62465 (.A(u0_n_32741),
    .B(u0_n_30271),
    .Y(u0_n_29963));
 OAI211xp5_ASAP7_75t_L u0_g62466 (.A1(u0_n_32141),
    .A2(u0_n_31314),
    .B(u0_n_30357),
    .C(u0_n_30413),
    .Y(u0_n_29964));
 OAI211xp5_ASAP7_75t_SL u0_g62467 (.A1(u0_n_32385),
    .A2(u0_n_31318),
    .B(u0_n_30352),
    .C(u0_n_30465),
    .Y(u0_n_29966));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62468 (.A1(w3[7]),
    .A2(u0_n_31633),
    .B(u0_n_30572),
    .C(u0_n_31968),
    .Y(u0_n_29968));
 OAI21xp33_ASAP7_75t_L u0_g62469 (.A1(u0_n_30909),
    .A2(u0_n_30549),
    .B(u0_n_31407),
    .Y(u0_n_29969));
 OAI21xp5_ASAP7_75t_SL u0_g62470 (.A1(u0_n_30720),
    .A2(u0_n_30532),
    .B(u0_n_30105),
    .Y(u0_n_29970));
 A2O1A1O1Ixp25_ASAP7_75t_R u0_g62471 (.A1(u0_n_32773),
    .A2(u0_n_31673),
    .B(u0_n_30762),
    .C(u0_n_31837),
    .D(u0_n_30560),
    .Y(u0_n_29971));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62472 (.A1(w3[3]),
    .A2(u0_n_31547),
    .B(u0_n_30561),
    .C(u0_n_31779),
    .Y(u0_n_29972));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62473 (.A1(\u0_w[3] [27]),
    .A2(u0_n_31549),
    .B(u0_n_30575),
    .C(u0_n_31774),
    .Y(u0_n_29973));
 OAI31xp33_ASAP7_75t_L u0_g62474 (.A1(u0_n_30577),
    .A2(u0_n_31350),
    .A3(u0_n_31624),
    .B(u0_n_31479),
    .Y(u0_n_29975));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62475 (.A1(u0_n_32023),
    .A2(u0_n_30771),
    .B(u0_n_30563),
    .C(u0_n_31787),
    .Y(u0_n_29976));
 OAI21xp33_ASAP7_75t_L u0_g62476 (.A1(u0_n_30567),
    .A2(u0_n_30356),
    .B(u0_n_31447),
    .Y(u0_n_29978));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62477 (.A1(u0_n_33004),
    .A2(u0_n_31489),
    .B(u0_n_30573),
    .C(u0_n_31771),
    .Y(u0_n_29980));
 OAI211xp5_ASAP7_75t_R u0_g62478 (.A1(u0_n_32387),
    .A2(u0_n_31548),
    .B(u0_n_30133),
    .C(u0_n_30741),
    .Y(u0_n_29981));
 NOR2xp33_ASAP7_75t_R u0_g62479 (.A(u0_n_31787),
    .B(u0_n_30261),
    .Y(u0_n_29983));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62480 (.A1(u0_n_32221),
    .A2(u0_n_30739),
    .B(u0_n_30611),
    .C(w3[18]),
    .Y(u0_n_29984));
 NAND3xp33_ASAP7_75t_R u0_g62481 (.A(u0_n_30369),
    .B(u0_n_30731),
    .C(u0_n_32839),
    .Y(u0_n_29986));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62482 (.A1(u0_n_32021),
    .A2(u0_n_30764),
    .B(u0_n_30599),
    .C(w3[18]),
    .Y(u0_n_29987));
 OAI332xp33_ASAP7_75t_SL u0_g62483 (.A1(u0_n_30890),
    .A2(u0_n_30391),
    .A3(u0_n_31346),
    .B1(u0_n_31410),
    .B2(u0_n_31533),
    .B3(u0_n_31924),
    .C1(u0_n_31132),
    .C2(u0_n_31758),
    .Y(u0_n_29988));
 NOR3xp33_ASAP7_75t_L u0_g62484 (.A(u0_n_30411),
    .B(u0_n_30550),
    .C(w3[26]),
    .Y(u0_n_29989));
 AOI322xp5_ASAP7_75t_R u0_g62485 (.A1(u0_n_31095),
    .A2(u0_n_32080),
    .A3(u0_n_31977),
    .B1(u0_n_31874),
    .B2(u0_n_31136),
    .C1(u0_n_31187),
    .C2(u0_n_30474),
    .Y(u0_n_29990));
 OAI322xp33_ASAP7_75t_L u0_g62486 (.A1(u0_n_31097),
    .A2(u0_n_32108),
    .A3(u0_n_31982),
    .B1(u0_n_31182),
    .B2(u0_n_30478),
    .C1(u0_n_31142),
    .C2(u0_n_32338),
    .Y(u0_n_29991));
 AOI322xp5_ASAP7_75t_R u0_g62487 (.A1(u0_n_31098),
    .A2(u0_n_31986),
    .A3(u0_n_31985),
    .B1(u0_n_32226),
    .B2(u0_n_31130),
    .C1(u0_n_30480),
    .C2(u0_n_31181),
    .Y(u0_n_29992));
 OAI211xp5_ASAP7_75t_L u0_g62488 (.A1(u0_n_32338),
    .A2(u0_n_31183),
    .B(u0_n_30337),
    .C(u0_n_30359),
    .Y(u0_n_29994));
 AOI322xp5_ASAP7_75t_R u0_g62489 (.A1(u0_n_31102),
    .A2(u0_n_32040),
    .A3(u0_n_31976),
    .B1(u0_n_32273),
    .B2(u0_n_31133),
    .C1(u0_n_30482),
    .C2(u0_n_31184),
    .Y(u0_n_29997));
 OAI21xp33_ASAP7_75t_R u0_g62490 (.A1(u0_n_30618),
    .A2(u0_n_30909),
    .B(u0_n_31798),
    .Y(u0_n_29999));
 OA21x2_ASAP7_75t_SL u0_g62491 (.A1(u0_n_30351),
    .A2(u0_n_30521),
    .B(u0_n_31390),
    .Y(u0_n_30001));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62492 (.A1(u0_n_32320),
    .A2(u0_n_31239),
    .B(u0_n_30453),
    .C(u0_n_31940),
    .Y(u0_n_30003));
 OAI33xp33_ASAP7_75t_SL u0_g62493 (.A1(u0_n_30941),
    .A2(u0_n_30922),
    .A3(u0_n_30371),
    .B1(u0_n_30535),
    .B2(u0_n_30926),
    .B3(u0_n_31115),
    .Y(u0_n_30004));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62494 (.A1(u0_n_32338),
    .A2(u0_n_30728),
    .B(u0_n_30667),
    .C(u0_n_31778),
    .Y(u0_n_30006));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62495 (.A1(u0_n_32184),
    .A2(u0_n_30756),
    .B(u0_n_30692),
    .C(w3[10]),
    .Y(u0_n_30008));
 AOI21xp33_ASAP7_75t_R u0_g62496 (.A1(u0_n_30900),
    .A2(u0_n_30592),
    .B(u0_n_31454),
    .Y(u0_n_30009));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62497 (.A1(u0_n_32260),
    .A2(u0_n_30772),
    .B(u0_n_32741),
    .C(u0_n_30119),
    .Y(u0_n_30011));
 OAI211xp5_ASAP7_75t_L u0_g62498 (.A1(u0_n_32410),
    .A2(u0_n_31091),
    .B(u0_n_30364),
    .C(u0_n_30380),
    .Y(u0_n_30013));
 AOI211xp5_ASAP7_75t_SL u0_g62499 (.A1(u0_n_31320),
    .A2(u0_n_32084),
    .B(u0_n_30348),
    .C(u0_n_30452),
    .Y(u0_n_30014));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62500 (.A1(u0_n_31841),
    .A2(u0_n_30761),
    .B(u0_n_30702),
    .C(u0_n_32747),
    .Y(u0_n_30016));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62501 (.A1(n_8801),
    .A2(u0_n_31166),
    .B(u0_n_30525),
    .C(u0_n_31783),
    .Y(u0_n_30017));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62502 (.A1(u0_n_31539),
    .A2(u0_n_31177),
    .B(u0_n_32353),
    .C(u0_n_30290),
    .Y(u0_n_30018));
 OAI311xp33_ASAP7_75t_L u0_g62503 (.A1(u0_n_31125),
    .A2(u0_n_31528),
    .A3(u0_n_32194),
    .B1(u0_n_30798),
    .C1(u0_n_30400),
    .Y(u0_n_30020));
 AOI211xp5_ASAP7_75t_L u0_g62504 (.A1(u0_n_30776),
    .A2(u0_n_32763),
    .B(u0_n_30969),
    .C(u0_n_30486),
    .Y(u0_n_30021));
 AOI311xp33_ASAP7_75t_SL u0_g62505 (.A1(u0_n_31163),
    .A2(u0_n_31841),
    .A3(u0_n_31531),
    .B(u0_n_30810),
    .C(u0_n_30398),
    .Y(u0_n_30022));
 AOI211xp5_ASAP7_75t_SL u0_g62506 (.A1(u0_n_31312),
    .A2(u0_n_31986),
    .B(u0_n_30354),
    .C(u0_n_30460),
    .Y(u0_n_30024));
 AOI311xp33_ASAP7_75t_R u0_g62507 (.A1(u0_n_31170),
    .A2(u0_n_31536),
    .A3(u0_n_32308),
    .B(u0_n_30814),
    .C(u0_n_30402),
    .Y(u0_n_30027));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62508 (.A1(u0_n_31175),
    .A2(u0_n_31186),
    .B(u0_n_32142),
    .C(u0_n_30198),
    .Y(u0_n_30028));
 OAI21xp33_ASAP7_75t_R u0_g62509 (.A1(u0_n_30626),
    .A2(u0_n_30348),
    .B(u0_n_31790),
    .Y(u0_n_30029));
 AOI211xp5_ASAP7_75t_L u0_g62510 (.A1(u0_n_30738),
    .A2(u0_n_32407),
    .B(u0_n_30717),
    .C(u0_n_30377),
    .Y(u0_n_30031));
 AOI21xp5_ASAP7_75t_SL u0_g62511 (.A1(u0_n_31123),
    .A2(u0_n_31841),
    .B(u0_n_30169),
    .Y(u0_n_30032));
 AO21x1_ASAP7_75t_R u0_g62512 (.A1(u0_n_30653),
    .A2(u0_n_30368),
    .B(u0_n_31932),
    .Y(u0_n_30033));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62513 (.A1(u0_n_31185),
    .A2(u0_n_31173),
    .B(u0_n_32386),
    .C(u0_n_30189),
    .Y(u0_n_30035));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62514 (.A1(u0_n_32221),
    .A2(u0_n_31178),
    .B(u0_n_30708),
    .C(u0_n_31958),
    .Y(u0_n_30037));
 OAI221xp5_ASAP7_75t_L u0_g62515 (.A1(u0_n_31162),
    .A2(u0_n_32338),
    .B1(u0_n_31392),
    .B2(u0_n_32108),
    .C(u0_n_30131),
    .Y(u0_n_30039));
 AOI221xp5_ASAP7_75t_SL u0_g62516 (.A1(u0_n_31141),
    .A2(u0_n_32273),
    .B1(u0_n_31569),
    .B2(u0_n_32063),
    .C(u0_n_30129),
    .Y(u0_n_30041));
 OAI211xp5_ASAP7_75t_L u0_g62517 (.A1(u0_n_32385),
    .A2(u0_n_31088),
    .B(u0_n_30361),
    .C(u0_n_30542),
    .Y(u0_n_30043));
 OAI21xp33_ASAP7_75t_R u0_g62518 (.A1(u0_n_30711),
    .A2(u0_n_30768),
    .B(u0_n_31973),
    .Y(u0_n_30044));
 OR3x1_ASAP7_75t_R u0_g62519 (.A(u0_n_30373),
    .B(u0_n_30725),
    .C(u0_n_32845),
    .Y(u0_n_30046));
 NAND3xp33_ASAP7_75t_R u0_g62520 (.A(u0_n_30373),
    .B(u0_n_30731),
    .C(u0_n_32835),
    .Y(u0_n_30047));
 AO21x1_ASAP7_75t_SL u0_g62521 (.A1(u0_n_32308),
    .A2(u0_n_31148),
    .B(u0_n_30140),
    .Y(u0_n_30049));
 NAND5xp2_ASAP7_75t_SL u0_g62522 (.A(u0_n_30876),
    .B(u0_n_31243),
    .C(u0_n_30997),
    .D(u0_n_31646),
    .E(u0_n_31425),
    .Y(u0_n_30051));
 OAI211xp5_ASAP7_75t_L u0_g62523 (.A1(u0_n_32017),
    .A2(u0_n_31149),
    .B(u0_n_30427),
    .C(u0_n_30408),
    .Y(u0_n_30052));
 AOI221xp5_ASAP7_75t_SL u0_g62524 (.A1(u0_n_31150),
    .A2(u0_n_32208),
    .B1(u0_n_31391),
    .B2(u0_n_31986),
    .C(u0_n_30128),
    .Y(u0_n_30054));
 OAI211xp5_ASAP7_75t_R u0_g62525 (.A1(u0_n_32774),
    .A2(u0_n_30905),
    .B(u0_n_30697),
    .C(u0_n_30766),
    .Y(u0_n_30056));
 AOI211xp5_ASAP7_75t_SL u0_g62526 (.A1(u0_n_30763),
    .A2(u0_n_31435),
    .B(u0_n_30586),
    .C(u0_n_30826),
    .Y(u0_n_30058));
 OAI221xp5_ASAP7_75t_SL u0_g62527 (.A1(u0_n_30739),
    .A2(u0_n_32017),
    .B1(u0_n_31289),
    .B2(u0_n_32795),
    .C(u0_n_30531),
    .Y(u0_n_30059));
 OAI21xp33_ASAP7_75t_L u0_g62528 (.A1(u0_n_31842),
    .A2(u0_n_30732),
    .B(u0_n_30309),
    .Y(u0_n_30062));
 AOI211xp5_ASAP7_75t_SL u0_g62529 (.A1(u0_n_30736),
    .A2(u0_n_32241),
    .B(u0_n_30723),
    .C(u0_n_30527),
    .Y(u0_n_30064));
 NAND5xp2_ASAP7_75t_L u0_g62530 (.A(u0_n_30406),
    .B(u0_n_30745),
    .C(u0_n_30872),
    .D(u0_n_31581),
    .E(u0_n_31425),
    .Y(u0_n_30066));
 OAI221xp5_ASAP7_75t_R u0_g62531 (.A1(u0_n_31131),
    .A2(u0_n_31161),
    .B1(u0_n_31139),
    .B2(u0_n_31145),
    .C(u0_n_30650),
    .Y(u0_n_30068));
 OAI221xp5_ASAP7_75t_SL u0_g62532 (.A1(u0_n_31147),
    .A2(u0_n_31152),
    .B1(u0_n_31157),
    .B2(u0_n_31149),
    .C(u0_n_30520),
    .Y(u0_n_30070));
 OAI221xp5_ASAP7_75t_R u0_g62533 (.A1(u0_n_31120),
    .A2(u0_n_32121),
    .B1(u0_n_31162),
    .B2(u0_n_32409),
    .C(u0_n_30683),
    .Y(u0_n_30072));
 OAI22xp33_ASAP7_75t_L u0_g62534 (.A1(u0_n_30467),
    .A2(w3[2]),
    .B1(u0_n_30775),
    .B2(u0_n_31758),
    .Y(u0_n_30076));
 AOI221xp5_ASAP7_75t_L u0_g62535 (.A1(u0_n_31106),
    .A2(u0_n_32353),
    .B1(u0_n_30757),
    .B2(u0_n_32113),
    .C(u0_n_30584),
    .Y(u0_n_30078));
 OAI211xp5_ASAP7_75t_R u0_g62536 (.A1(u0_n_31474),
    .A2(u0_n_31233),
    .B(u0_n_30438),
    .C(u0_n_31192),
    .Y(u0_n_30080));
 AOI211xp5_ASAP7_75t_R u0_g62537 (.A1(u0_n_31440),
    .A2(u0_n_31923),
    .B(u0_n_30799),
    .C(u0_n_30449),
    .Y(u0_n_30081));
 AOI221xp5_ASAP7_75t_SL u0_g62538 (.A1(u0_n_31234),
    .A2(u0_n_31460),
    .B1(u0_n_30489),
    .B2(u0_n_32747),
    .C(u0_n_30388),
    .Y(u0_n_30082));
 AO221x1_ASAP7_75t_SL u0_g62539 (.A1(u0_n_30760),
    .A2(u0_n_32073),
    .B1(u0_n_31320),
    .B2(u0_n_32166),
    .C(u0_n_30654),
    .Y(u0_n_30083));
 OAI221xp5_ASAP7_75t_R u0_g62540 (.A1(u0_n_30765),
    .A2(u0_n_32042),
    .B1(u0_n_31323),
    .B2(u0_n_32387),
    .C(u0_n_30663),
    .Y(u0_n_30087));
 OAI221xp5_ASAP7_75t_R u0_g62541 (.A1(u0_n_31291),
    .A2(u0_n_31964),
    .B1(u0_n_31320),
    .B2(u0_n_32141),
    .C(u0_n_30674),
    .Y(u0_n_30090));
 AOI221xp5_ASAP7_75t_L u0_g62542 (.A1(u0_n_31312),
    .A2(u0_n_32241),
    .B1(u0_n_30763),
    .B2(u0_n_31998),
    .C(u0_n_30670),
    .Y(u0_n_30092));
 OAI221xp5_ASAP7_75t_L u0_g62543 (.A1(u0_n_30910),
    .A2(u0_n_33004),
    .B1(u0_n_30853),
    .B2(u0_n_32209),
    .C(u0_n_30849),
    .Y(u0_n_30094));
 AOI211xp5_ASAP7_75t_L u0_g62544 (.A1(u0_n_31311),
    .A2(u0_n_31830),
    .B(u0_n_30640),
    .C(u0_n_31454),
    .Y(u0_n_30096));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62545 (.A1(u0_n_32040),
    .A2(u0_n_31549),
    .B(u0_n_30740),
    .C(u0_n_32743),
    .Y(u0_n_30099));
 OAI221xp5_ASAP7_75t_R u0_g62546 (.A1(u0_n_31632),
    .A2(n_8831),
    .B1(u0_n_31600),
    .B2(u0_n_32242),
    .C(u0_n_31068),
    .Y(u0_n_30101));
 OAI211xp5_ASAP7_75t_SL u0_g62547 (.A1(u0_n_32108),
    .A2(u0_n_31322),
    .B(u0_n_30355),
    .C(u0_n_30789),
    .Y(u0_n_30102));
 AOI31xp33_ASAP7_75t_L u0_g62548 (.A1(u0_n_31260),
    .A2(u0_n_30953),
    .A3(u0_n_31355),
    .B(w3[10]),
    .Y(u0_n_30104));
 A2O1A1O1Ixp25_ASAP7_75t_SL u0_g62549 (.A1(u0_n_31810),
    .A2(u0_n_31874),
    .B(u0_n_31422),
    .C(w3[0]),
    .D(u0_n_30546),
    .Y(u0_n_30105));
 NOR2xp33_ASAP7_75t_R u0_g62550 (.A(u0_n_30576),
    .B(u0_n_30743),
    .Y(u0_n_30108));
 NOR4xp25_ASAP7_75t_R u0_g62551 (.A(u0_n_30350),
    .B(u0_n_30824),
    .C(u0_n_31119),
    .D(u0_n_31247),
    .Y(u0_n_30109));
 AOI211xp5_ASAP7_75t_L u0_g62552 (.A1(u0_n_31132),
    .A2(u0_n_32073),
    .B(u0_n_30349),
    .C(u0_n_30854),
    .Y(u0_n_30111));
 AOI211xp5_ASAP7_75t_R u0_g62553 (.A1(u0_n_31275),
    .A2(u0_n_31478),
    .B(u0_n_30828),
    .C(u0_n_30822),
    .Y(u0_n_30114));
 A2O1A1O1Ixp25_ASAP7_75t_SL u0_g62554 (.A1(n_8801),
    .A2(u0_n_31970),
    .B(u0_n_32407),
    .C(u0_n_31166),
    .D(u0_n_30363),
    .Y(u0_n_30115));
 OAI211xp5_ASAP7_75t_SL u0_g62555 (.A1(u0_n_31988),
    .A2(u0_n_31294),
    .B(u0_n_30464),
    .C(u0_n_31027),
    .Y(u0_n_30119));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62556 (.A1(u0_n_32425),
    .A2(u0_n_31324),
    .B(u0_n_30875),
    .C(u0_n_30915),
    .Y(u0_n_30120));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62557 (.A1(u0_n_32141),
    .A2(u0_n_31327),
    .B(u0_n_30777),
    .C(u0_n_30820),
    .Y(u0_n_30121));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62558 (.A1(u0_n_32774),
    .A2(u0_n_31144),
    .B(u0_n_30837),
    .C(u0_n_31419),
    .Y(u0_n_30122));
 OAI211xp5_ASAP7_75t_SL u0_g62559 (.A1(u0_n_32409),
    .A2(u0_n_31612),
    .B(u0_n_31070),
    .C(u0_n_31297),
    .Y(u0_n_30123));
 AOI211xp5_ASAP7_75t_R u0_g62560 (.A1(u0_n_31606),
    .A2(u0_n_32373),
    .B(u0_n_31036),
    .C(u0_n_31295),
    .Y(u0_n_30124));
 OAI221xp5_ASAP7_75t_L u0_g62561 (.A1(u0_n_31327),
    .A2(u0_n_31766),
    .B1(u0_n_31459),
    .B2(u0_n_31434),
    .C(u0_n_30484),
    .Y(u0_n_30126));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62562 (.A1(w3[19]),
    .A2(u0_n_31264),
    .B(u0_n_30802),
    .C(u0_n_33001),
    .Y(u0_n_30128));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62563 (.A1(\u0_w[3] [27]),
    .A2(u0_n_31281),
    .B(u0_n_30804),
    .C(w3[30]),
    .Y(u0_n_30129));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62564 (.A1(w3[11]),
    .A2(u0_n_31285),
    .B(u0_n_30806),
    .C(n_8801),
    .Y(u0_n_30131));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62565 (.A1(u0_n_33004),
    .A2(u0_n_31143),
    .B(u0_n_30835),
    .C(u0_n_31950),
    .Y(u0_n_30132));
 AOI211xp5_ASAP7_75t_R u0_g62566 (.A1(u0_n_31274),
    .A2(u0_n_32063),
    .B(u0_n_31458),
    .C(u0_n_31254),
    .Y(u0_n_30133));
 OAI211xp5_ASAP7_75t_L u0_g62567 (.A1(u0_n_31842),
    .A2(u0_n_31145),
    .B(u0_n_30747),
    .C(u0_n_31353),
    .Y(u0_n_30134));
 AOI211xp5_ASAP7_75t_L u0_g62568 (.A1(u0_n_31347),
    .A2(u0_n_33004),
    .B(u0_n_31004),
    .C(w3[18]),
    .Y(u0_n_30136));
 AOI321xp33_ASAP7_75t_L u0_g62569 (.A1(u0_n_31662),
    .A2(\u0_w[3] [16]),
    .A3(w3[19]),
    .B1(u0_n_31822),
    .B2(u0_n_32208),
    .C(u0_n_30845),
    .Y(u0_n_30137));
 NAND4xp25_ASAP7_75t_L u0_g62570 (.A(u0_n_30367),
    .B(u0_n_31043),
    .C(u0_n_31082),
    .D(u0_n_31419),
    .Y(u0_n_30138));
 OAI221xp5_ASAP7_75t_SL u0_g62571 (.A1(u0_n_32042),
    .A2(u0_n_31256),
    .B1(u0_n_32372),
    .B2(u0_n_31683),
    .C(u0_n_30737),
    .Y(u0_n_30140));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62572 (.A1(u0_n_31817),
    .A2(u0_n_31177),
    .B(u0_n_32109),
    .C(u0_n_30558),
    .Y(u0_n_30141));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62573 (.A1(u0_n_32121),
    .A2(u0_n_31541),
    .B(u0_n_30745),
    .C(n_11401),
    .Y(u0_n_30144));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62574 (.A1(u0_n_31837),
    .A2(u0_n_31174),
    .B(u0_n_32075),
    .C(u0_n_30555),
    .Y(u0_n_30146));
 OAI221xp5_ASAP7_75t_SL u0_g62575 (.A1(u0_n_31250),
    .A2(u0_n_31988),
    .B1(u0_n_32254),
    .B2(u0_n_31535),
    .C(u0_n_30742),
    .Y(u0_n_30148));
 AOI221xp5_ASAP7_75t_SL u0_g62576 (.A1(u0_n_31255),
    .A2(u0_n_32084),
    .B1(u0_n_31533),
    .B2(u0_n_32142),
    .C(u0_n_30762),
    .Y(u0_n_30150));
 AOI221xp5_ASAP7_75t_SL u0_g62577 (.A1(u0_n_31251),
    .A2(u0_n_32122),
    .B1(u0_n_31539),
    .B2(u0_n_32407),
    .C(u0_n_30744),
    .Y(u0_n_30153));
 OAI211xp5_ASAP7_75t_L u0_g62578 (.A1(u0_n_32023),
    .A2(u0_n_31287),
    .B(u0_n_30921),
    .C(u0_n_30724),
    .Y(u0_n_30155));
 AOI221xp5_ASAP7_75t_R u0_g62579 (.A1(u0_n_31612),
    .A2(u0_n_32407),
    .B1(u0_n_31636),
    .B2(u0_n_32714),
    .C(u0_n_31061),
    .Y(u0_n_30156));
 OAI311xp33_ASAP7_75t_L u0_g62580 (.A1(u0_n_31686),
    .A2(u0_n_31674),
    .A3(u0_n_32194),
    .B1(u0_n_31014),
    .C1(u0_n_31118),
    .Y(u0_n_30158));
 OAI211xp5_ASAP7_75t_R u0_g62581 (.A1(u0_n_32321),
    .A2(u0_n_31135),
    .B(u0_n_30461),
    .C(u0_n_31774),
    .Y(u0_n_30159));
 AOI211xp5_ASAP7_75t_R u0_g62582 (.A1(u0_n_31276),
    .A2(u0_n_32073),
    .B(u0_n_30501),
    .C(u0_n_31023),
    .Y(u0_n_30160));
 OAI211xp5_ASAP7_75t_R u0_g62583 (.A1(u0_n_31842),
    .A2(u0_n_31144),
    .B(u0_n_30454),
    .C(u0_n_31779),
    .Y(u0_n_30161));
 OAI221xp5_ASAP7_75t_R u0_g62584 (.A1(u0_n_30754),
    .A2(u0_n_30958),
    .B1(u0_n_31143),
    .B2(u0_n_32023),
    .C(u0_n_31770),
    .Y(u0_n_30163));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62585 (.A1(u0_n_31799),
    .A2(u0_n_32208),
    .B(u0_n_30996),
    .C(u0_n_31089),
    .Y(u0_n_30165));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62586 (.A1(u0_n_31825),
    .A2(u0_n_31125),
    .B(u0_n_32416),
    .C(u0_n_30551),
    .Y(u0_n_30166));
 AOI21xp33_ASAP7_75t_R u0_g62587 (.A1(u0_n_32320),
    .A2(u0_n_30765),
    .B(u0_n_30595),
    .Y(u0_n_30168));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62588 (.A1(u0_n_31689),
    .A2(u0_n_31677),
    .B(u0_n_32165),
    .C(u0_n_30459),
    .Y(u0_n_30169));
 OAI211xp5_ASAP7_75t_R u0_g62589 (.A1(u0_n_33033),
    .A2(u0_n_30755),
    .B(u0_n_30741),
    .C(u0_n_31774),
    .Y(u0_n_30170));
 AOI211xp5_ASAP7_75t_SL u0_g62590 (.A1(u0_n_31303),
    .A2(u0_n_32193),
    .B(u0_n_30717),
    .C(u0_n_30938),
    .Y(u0_n_30172));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62591 (.A1(u0_n_31822),
    .A2(u0_n_31179),
    .B(u0_n_31998),
    .C(u0_n_30553),
    .Y(u0_n_30176));
 OAI211xp5_ASAP7_75t_R u0_g62592 (.A1(u0_n_31484),
    .A2(u0_n_31633),
    .B(u0_n_30964),
    .C(u0_n_30471),
    .Y(u0_n_30178));
 A2O1A1Ixp33_ASAP7_75t_SL u0_g62593 (.A1(u0_n_31830),
    .A2(u0_n_31172),
    .B(u0_n_32042),
    .C(u0_n_30557),
    .Y(u0_n_30180));
 AOI21xp33_ASAP7_75t_R u0_g62594 (.A1(u0_n_32021),
    .A2(u0_n_30751),
    .B(u0_n_31005),
    .Y(u0_n_30182));
 AOI221xp5_ASAP7_75t_SL u0_g62595 (.A1(u0_n_31121),
    .A2(u0_n_31583),
    .B1(u0_n_31138),
    .B2(u0_n_31809),
    .C(u0_n_30632),
    .Y(u0_n_30183));
 AOI221xp5_ASAP7_75t_SL u0_g62596 (.A1(u0_n_31311),
    .A2(u0_n_31959),
    .B1(u0_n_31323),
    .B2(u0_n_32386),
    .C(u0_n_30492),
    .Y(u0_n_30185));
 OAI222xp33_ASAP7_75t_R u0_g62597 (.A1(u0_n_31318),
    .A2(u0_n_31335),
    .B1(u0_n_31273),
    .B2(u0_n_33033),
    .C1(u0_n_31805),
    .C2(u0_n_32387),
    .Y(u0_n_30187));
 OAI211xp5_ASAP7_75t_L u0_g62598 (.A1(u0_n_31792),
    .A2(u0_n_31279),
    .B(u0_n_30730),
    .C(u0_n_30978),
    .Y(u0_n_30189));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62599 (.A1(u0_n_32373),
    .A2(u0_n_31330),
    .B(u0_n_30778),
    .C(u0_n_31774),
    .Y(u0_n_30190));
 AOI221xp5_ASAP7_75t_SL u0_g62600 (.A1(u0_n_31634),
    .A2(u0_n_31651),
    .B1(u0_n_31278),
    .B2(u0_n_31823),
    .C(u0_n_30988),
    .Y(u0_n_30191));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62601 (.A1(u0_n_31916),
    .A2(u0_n_31167),
    .B(u0_n_31752),
    .C(u0_n_30928),
    .Y(u0_n_30192));
 OAI211xp5_ASAP7_75t_L u0_g62602 (.A1(u0_n_32017),
    .A2(u0_n_31240),
    .B(u0_n_31011),
    .C(u0_n_31092),
    .Y(u0_n_30193));
 AOI221xp5_ASAP7_75t_R u0_g62603 (.A1(u0_n_31263),
    .A2(n_8801),
    .B1(u0_n_32416),
    .B2(u0_n_31801),
    .C(u0_n_30784),
    .Y(u0_n_30194));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62604 (.A1(u0_n_31988),
    .A2(u0_n_31544),
    .B(u0_n_30911),
    .C(\u0_w[3] [16]),
    .Y(u0_n_30195));
 OAI311xp33_ASAP7_75t_SL u0_g62605 (.A1(u0_n_31688),
    .A2(u0_n_31676),
    .A3(u0_n_31842),
    .B1(u0_n_31016),
    .C1(u0_n_31096),
    .Y(u0_n_30196));
 OAI21xp33_ASAP7_75t_SL u0_g62606 (.A1(u0_n_32793),
    .A2(u0_n_31269),
    .B(u0_n_30390),
    .Y(u0_n_30197));
 OAI211xp5_ASAP7_75t_SL u0_g62607 (.A1(u0_n_31796),
    .A2(u0_n_31241),
    .B(u0_n_30719),
    .C(u0_n_30985),
    .Y(u0_n_30198));
 AOI221xp5_ASAP7_75t_L u0_g62608 (.A1(u0_n_31144),
    .A2(u0_n_31874),
    .B1(u0_n_31602),
    .B2(u0_n_32073),
    .C(u0_n_30493),
    .Y(u0_n_30199));
 AOI211xp5_ASAP7_75t_L u0_g62609 (.A1(u0_n_31363),
    .A2(u0_n_32339),
    .B(u0_n_30652),
    .C(u0_n_30718),
    .Y(u0_n_30200));
 NAND4xp25_ASAP7_75t_L u0_g62610 (.A(u0_n_30368),
    .B(u0_n_31045),
    .C(u0_n_31452),
    .D(u0_n_31083),
    .Y(u0_n_30201));
 NOR3xp33_ASAP7_75t_R u0_g62612 (.A(u0_n_30773),
    .B(u0_n_30725),
    .C(u0_r0_rcnt[0]),
    .Y(u0_n_30098));
 OAI221xp5_ASAP7_75t_R u0_g62614 (.A1(u0_n_31635),
    .A2(u0_n_32717),
    .B1(u0_n_31606),
    .B2(u0_n_32372),
    .C(u0_n_31063),
    .Y(u0_n_30204));
 OAI221xp5_ASAP7_75t_L u0_g62615 (.A1(u0_n_31489),
    .A2(u0_n_32017),
    .B1(u0_n_32249),
    .B2(u0_n_31609),
    .C(u0_n_30679),
    .Y(u0_n_30207));
 AO21x1_ASAP7_75t_L u0_g62616 (.A1(u0_n_32289),
    .A2(u0_n_30735),
    .B(u0_n_30614),
    .Y(u0_n_30209));
 OAI21xp33_ASAP7_75t_L u0_g62617 (.A1(u0_n_31886),
    .A2(u0_n_30732),
    .B(u0_n_30672),
    .Y(u0_n_30211));
 OR4x1_ASAP7_75t_R u0_g62618 (.A(u0_n_30370),
    .B(u0_n_31041),
    .C(u0_n_31458),
    .D(u0_n_31087),
    .Y(u0_n_30214));
 AO21x1_ASAP7_75t_SL u0_g62619 (.A1(u0_n_31998),
    .A2(u0_n_31257),
    .B(u0_n_30360),
    .Y(u0_n_30215));
 OAI221xp5_ASAP7_75t_L u0_g62620 (.A1(u0_n_31081),
    .A2(u0_n_31988),
    .B1(u0_n_31821),
    .B2(u0_n_32017),
    .C(u0_n_30980),
    .Y(u0_n_30217));
 AOI211xp5_ASAP7_75t_SL u0_g62621 (.A1(u0_n_31141),
    .A2(u0_n_32320),
    .B(u0_n_30740),
    .C(u0_n_31198),
    .Y(u0_n_30218));
 OAI211xp5_ASAP7_75t_SL u0_g62622 (.A1(u0_n_31969),
    .A2(u0_n_31299),
    .B(u0_n_30591),
    .C(u0_n_30998),
    .Y(u0_n_30221));
 OAI221xp5_ASAP7_75t_SL u0_g62623 (.A1(u0_n_31128),
    .A2(u0_n_31691),
    .B1(u0_n_31159),
    .B2(u0_n_31808),
    .C(u0_n_30647),
    .Y(u0_n_30223));
 OAI322xp33_ASAP7_75t_R u0_g62624 (.A1(u0_n_31258),
    .A2(u0_n_32075),
    .A3(u0_n_32695),
    .B1(u0_n_31426),
    .B2(u0_n_31195),
    .C1(u0_n_31410),
    .C2(u0_n_31837),
    .Y(u0_n_30224));
 OAI21xp33_ASAP7_75t_R u0_g62625 (.A1(u0_n_32773),
    .A2(u0_n_31123),
    .B(u0_n_30392),
    .Y(u0_n_30229));
 OAI21xp33_ASAP7_75t_SL u0_g62626 (.A1(u0_n_32121),
    .A2(u0_n_31305),
    .B(u0_n_30685),
    .Y(u0_n_30232));
 AOI221xp5_ASAP7_75t_SL u0_g62627 (.A1(u0_n_31103),
    .A2(u0_n_32012),
    .B1(u0_n_32260),
    .B2(u0_n_31287),
    .C(u0_n_30415),
    .Y(u0_n_30233));
 OAI211xp5_ASAP7_75t_L u0_g62628 (.A1(u0_n_32385),
    .A2(u0_n_31117),
    .B(u0_n_30690),
    .C(u0_n_30737),
    .Y(u0_n_30235));
 OAI221xp5_ASAP7_75t_R u0_g62629 (.A1(u0_n_31541),
    .A2(u0_n_32749),
    .B1(u0_n_31502),
    .B2(n_8820),
    .C(u0_n_31000),
    .Y(u0_n_30237));
 AOI221xp5_ASAP7_75t_R u0_g62630 (.A1(u0_n_31322),
    .A2(u0_n_32193),
    .B1(u0_n_30752),
    .B2(u0_n_32416),
    .C(u0_n_31334),
    .Y(u0_n_30240));
 OAI321xp33_ASAP7_75t_L u0_g62631 (.A1(u0_n_31653),
    .A2(u0_n_31526),
    .A3(u0_n_32075),
    .B1(n_8629),
    .B2(u0_n_31875),
    .C(u0_n_30791),
    .Y(u0_n_30242));
 OAI211xp5_ASAP7_75t_SL u0_g62632 (.A1(u0_n_31474),
    .A2(u0_n_31286),
    .B(u0_n_31764),
    .C(u0_n_30476),
    .Y(u0_n_30244));
 AOI211xp5_ASAP7_75t_R u0_g62633 (.A1(u0_n_31116),
    .A2(u0_n_32416),
    .B(u0_n_30744),
    .C(u0_n_30695),
    .Y(u0_n_30247));
 OAI211xp5_ASAP7_75t_R u0_g62634 (.A1(u0_n_32194),
    .A2(u0_n_31313),
    .B(u0_n_30495),
    .C(u0_n_30793),
    .Y(u0_n_30249));
 OAI211xp5_ASAP7_75t_L u0_g62635 (.A1(n_8748),
    .A2(u0_n_31139),
    .B(u0_n_30396),
    .C(u0_n_30808),
    .Y(u0_n_30250));
 OAI221xp5_ASAP7_75t_L u0_g62636 (.A1(u0_n_31147),
    .A2(u0_n_31692),
    .B1(u0_n_31157),
    .B2(w3[17]),
    .C(u0_n_30522),
    .Y(u0_n_30252));
 NOR4xp25_ASAP7_75t_R u0_g62637 (.A(u0_n_30538),
    .B(u0_n_31252),
    .C(u0_n_31114),
    .D(u0_n_31515),
    .Y(u0_n_30255));
 AOI211xp5_ASAP7_75t_R u0_g62638 (.A1(u0_n_31109),
    .A2(u0_n_32142),
    .B(u0_n_30762),
    .C(u0_n_30698),
    .Y(u0_n_30257));
 OR4x1_ASAP7_75t_R u0_g62639 (.A(u0_n_31370),
    .B(u0_n_30543),
    .C(u0_n_31119),
    .D(u0_n_31517),
    .Y(u0_n_30258));
 AOI221xp5_ASAP7_75t_R u0_g62640 (.A1(u0_n_31619),
    .A2(u0_n_32021),
    .B1(u0_n_32208),
    .B2(u0_n_31650),
    .C(u0_n_31001),
    .Y(u0_n_30261));
 AOI221xp5_ASAP7_75t_R u0_g62641 (.A1(u0_n_31850),
    .A2(u0_n_31526),
    .B1(u0_n_32073),
    .B2(u0_n_31677),
    .C(u0_n_31064),
    .Y(u0_n_30263));
 AOI221xp5_ASAP7_75t_R u0_g62642 (.A1(u0_n_32012),
    .A2(u0_n_31522),
    .B1(u0_n_31678),
    .B2(u0_n_31986),
    .C(u0_n_31072),
    .Y(u0_n_30266));
 AOI221xp5_ASAP7_75t_R u0_g62643 (.A1(u0_n_32184),
    .A2(u0_n_31524),
    .B1(u0_n_31675),
    .B2(u0_n_32109),
    .C(u0_n_31065),
    .Y(u0_n_30267));
 OAI21xp33_ASAP7_75t_L u0_g62644 (.A1(u0_n_31762),
    .A2(u0_n_30907),
    .B(u0_n_30606),
    .Y(u0_n_30268));
 AOI221xp5_ASAP7_75t_R u0_g62645 (.A1(u0_n_31323),
    .A2(u0_n_32308),
    .B1(u0_n_30770),
    .B2(u0_n_32373),
    .C(u0_n_31019),
    .Y(u0_n_30269));
 OAI211xp5_ASAP7_75t_SL u0_g62646 (.A1(w3[30]),
    .A2(u0_n_31054),
    .B(u0_n_30831),
    .C(u0_n_31516),
    .Y(u0_n_30270));
 OAI322xp33_ASAP7_75t_R u0_g62647 (.A1(u0_n_31317),
    .A2(u0_n_31354),
    .A3(u0_n_32795),
    .B1(u0_n_31283),
    .B2(u0_n_33004),
    .C1(u0_n_32242),
    .C2(u0_n_31812),
    .Y(u0_n_30271));
 OAI211xp5_ASAP7_75t_L u0_g62648 (.A1(u0_n_32023),
    .A2(u0_n_31329),
    .B(u0_n_30796),
    .C(u0_n_30868),
    .Y(u0_n_30273));
 AOI221xp5_ASAP7_75t_R u0_g62649 (.A1(u0_n_31308),
    .A2(u0_n_31965),
    .B1(u0_n_31328),
    .B2(u0_n_31998),
    .C(u0_n_31002),
    .Y(u0_n_30274));
 OAI222xp33_ASAP7_75t_L u0_g62650 (.A1(u0_n_31151),
    .A2(u0_n_32338),
    .B1(u0_n_31304),
    .B2(n_8820),
    .C1(u0_n_31599),
    .C2(u0_n_32121),
    .Y(u0_n_30276));
 AOI222xp33_ASAP7_75t_SL u0_g62651 (.A1(u0_n_32208),
    .A2(u0_n_31143),
    .B1(u0_n_31619),
    .B2(u0_n_31998),
    .C1(u0_n_31306),
    .C2(u0_n_32795),
    .Y(u0_n_30277));
 OAI21xp33_ASAP7_75t_L u0_g62652 (.A1(w3[30]),
    .A2(u0_n_31310),
    .B(u0_n_30688),
    .Y(u0_n_30279));
 OAI221xp5_ASAP7_75t_R u0_g62653 (.A1(u0_n_31137),
    .A2(u0_n_32272),
    .B1(u0_n_32306),
    .B2(u0_n_31824),
    .C(u0_n_30858),
    .Y(u0_n_30280));
 AOI321xp33_ASAP7_75t_SL u0_g62654 (.A1(u0_n_31665),
    .A2(u0_n_31525),
    .A3(u0_n_32113),
    .B1(u0_n_31300),
    .B2(u0_n_31818),
    .C(u0_n_30914),
    .Y(u0_n_30283));
 OA222x2_ASAP7_75t_L u0_g62655 (.A1(u0_n_30761),
    .A2(u0_n_31426),
    .B1(u0_n_31320),
    .B2(u0_n_31410),
    .C1(u0_n_31551),
    .C2(u0_n_31758),
    .Y(u0_n_30284));
 OAI21xp33_ASAP7_75t_L u0_g62656 (.A1(u0_n_31766),
    .A2(u0_n_30905),
    .B(u0_n_30680),
    .Y(u0_n_30286));
 OAI211xp5_ASAP7_75t_SL u0_g62657 (.A1(u0_n_31059),
    .A2(u0_n_33001),
    .B(u0_n_30983),
    .C(u0_n_31512),
    .Y(u0_n_30289));
 OAI21xp33_ASAP7_75t_L u0_g62658 (.A1(w3[14]),
    .A2(u0_n_30907),
    .B(u0_n_30851),
    .Y(u0_n_30290));
 OAI221xp5_ASAP7_75t_SL u0_g62659 (.A1(u0_n_31270),
    .A2(u0_n_32108),
    .B1(u0_n_31637),
    .B2(u0_n_31470),
    .C(u0_n_30959),
    .Y(u0_n_30292));
 OAI321xp33_ASAP7_75t_L u0_g62660 (.A1(u0_n_31686),
    .A2(u0_n_32121),
    .A3(u0_n_31794),
    .B1(u0_n_32410),
    .B2(u0_n_31313),
    .C(u0_n_30976),
    .Y(u0_n_30293));
 OAI221xp5_ASAP7_75t_R u0_g62661 (.A1(u0_n_30760),
    .A2(u0_n_31842),
    .B1(u0_n_31302),
    .B2(u0_n_31886),
    .C(u0_n_31096),
    .Y(u0_n_30296));
 OAI321xp33_ASAP7_75t_L u0_g62662 (.A1(u0_n_31644),
    .A2(u0_n_31499),
    .A3(u0_n_31550),
    .B1(u0_n_32763),
    .B2(u0_n_31050),
    .C(u0_n_31514),
    .Y(u0_n_30298));
 OAI221xp5_ASAP7_75t_SL u0_g62663 (.A1(u0_n_32793),
    .A2(u0_n_31262),
    .B1(u0_n_32272),
    .B2(u0_n_31792),
    .C(u0_n_30971),
    .Y(u0_n_30299));
 AOI221xp5_ASAP7_75t_SL u0_g62664 (.A1(u0_n_31270),
    .A2(w3[14]),
    .B1(u0_n_32353),
    .B2(u0_n_31793),
    .C(u0_n_30972),
    .Y(u0_n_30302));
 AO332x1_ASAP7_75t_L u0_g62665 (.A1(u0_n_31102),
    .A2(u0_n_32304),
    .A3(u0_n_31976),
    .B1(u0_n_31519),
    .B2(u0_n_31683),
    .B3(u0_n_32373),
    .C1(u0_n_31137),
    .C2(u0_n_32040),
    .Y(u0_n_30304));
 AOI221xp5_ASAP7_75t_L u0_g62666 (.A1(u0_n_31268),
    .A2(u0_n_32774),
    .B1(u0_n_31874),
    .B2(u0_n_31795),
    .C(u0_n_30975),
    .Y(u0_n_30309));
 AO332x1_ASAP7_75t_L u0_g62667 (.A1(u0_n_31098),
    .A2(u0_n_32012),
    .A3(u0_n_31985),
    .B1(u0_n_31523),
    .B2(u0_n_31535),
    .B3(u0_n_32241),
    .C1(u0_n_31164),
    .C2(u0_n_31998),
    .Y(u0_n_30310));
 AOI332xp33_ASAP7_75t_R u0_g62668 (.A1(u0_n_31095),
    .A2(u0_n_31850),
    .A3(u0_n_31977),
    .B1(u0_n_31532),
    .B2(u0_n_32166),
    .B3(u0_n_31527),
    .C1(u0_n_31155),
    .C2(u0_n_32073),
    .Y(u0_n_30314));
 OA332x1_ASAP7_75t_L u0_g62669 (.A1(u0_n_31097),
    .A2(u0_n_32185),
    .A3(u0_n_31982),
    .B1(u0_n_31539),
    .B2(u0_n_31524),
    .B3(u0_n_32409),
    .C1(u0_n_31156),
    .C2(u0_n_32108),
    .Y(u0_n_30317));
 AOI211xp5_ASAP7_75t_L u0_g62670 (.A1(u0_n_30750),
    .A2(u0_n_32184),
    .B(u0_n_30718),
    .C(u0_n_30786),
    .Y(u0_n_30321));
 AOI221xp5_ASAP7_75t_L u0_g62671 (.A1(u0_n_31541),
    .A2(u0_n_32113),
    .B1(u0_n_31270),
    .B2(u0_n_32339),
    .C(u0_n_31057),
    .Y(u0_n_30323));
 OAI22xp33_ASAP7_75t_L u0_g62672 (.A1(w3[30]),
    .A2(u0_n_30903),
    .B1(u0_n_31683),
    .B2(u0_n_32272),
    .Y(u0_n_30324));
 OAI322xp33_ASAP7_75t_R u0_g62673 (.A1(u0_n_31546),
    .A2(u0_n_31886),
    .A3(u0_n_31838),
    .B1(u0_n_31267),
    .B2(u0_n_32141),
    .C1(u0_n_31105),
    .C2(u0_n_31842),
    .Y(u0_n_30326));
 AOI221xp5_ASAP7_75t_R u0_g62675 (.A1(u0_n_31544),
    .A2(u0_n_31998),
    .B1(u0_n_31290),
    .B2(u0_n_32226),
    .C(u0_n_31069),
    .Y(u0_n_30330));
 OAI221xp5_ASAP7_75t_R u0_g62676 (.A1(u0_n_31262),
    .A2(u0_n_32272),
    .B1(u0_n_31549),
    .B2(u0_n_32053),
    .C(u0_n_31073),
    .Y(u0_n_30332));
 AOI221xp5_ASAP7_75t_L u0_g62677 (.A1(u0_n_31546),
    .A2(u0_n_32084),
    .B1(u0_n_31268),
    .B2(u0_n_31874),
    .C(u0_n_31066),
    .Y(u0_n_30334));
 AOI211xp5_ASAP7_75t_SL u0_g62678 (.A1(u0_n_31177),
    .A2(u0_n_32109),
    .B(u0_n_31778),
    .C(u0_n_30746),
    .Y(u0_n_30337));
 AOI322xp5_ASAP7_75t_L u0_g62679 (.A1(u0_n_31549),
    .A2(u0_n_31830),
    .A3(u0_n_32289),
    .B1(u0_n_32304),
    .B2(u0_n_31113),
    .C1(u0_n_31277),
    .C2(u0_n_32386),
    .Y(u0_n_30339));
 OAI221xp5_ASAP7_75t_R u0_g62680 (.A1(u0_n_31174),
    .A2(u0_n_32083),
    .B1(u0_n_31100),
    .B2(u0_n_31842),
    .C(u0_n_31779),
    .Y(u0_n_30341));
 AOI211xp5_ASAP7_75t_R u0_g62681 (.A1(u0_n_31179),
    .A2(u0_n_31998),
    .B(u0_n_30913),
    .C(u0_n_31771),
    .Y(u0_n_30343));
 AOI211xp5_ASAP7_75t_L u0_g62682 (.A1(u0_n_31269),
    .A2(u0_n_32320),
    .B(u0_n_30992),
    .C(u0_n_30847),
    .Y(u0_n_30346));
 INVxp33_ASAP7_75t_R u0_g62683 (.A(u0_n_30362),
    .Y(u0_n_30361));
 INVx1_ASAP7_75t_SL u0_g62684 (.A(u0_n_30364),
    .Y(u0_n_30363));
 INVxp33_ASAP7_75t_R u0_g62685 (.A(u0_n_30366),
    .Y(u0_n_30365));
 INVxp67_ASAP7_75t_L u0_g62686 (.A(u0_n_30372),
    .Y(u0_n_30371));
 OAI321xp33_ASAP7_75t_L u0_g62687 (.A1(u0_n_32306),
    .A2(u0_n_31823),
    .A3(n_8942),
    .B1(u0_n_32387),
    .B2(u0_n_31413),
    .C(u0_n_30952),
    .Y(u0_n_30375));
 OAI21xp33_ASAP7_75t_R u0_g62688 (.A1(u0_n_31794),
    .A2(u0_n_31243),
    .B(u0_n_30986),
    .Y(u0_n_30377));
 OAI21xp33_ASAP7_75t_R u0_g62689 (.A1(u0_n_31818),
    .A2(u0_n_32184),
    .B(u0_n_30932),
    .Y(u0_n_30380));
 OAI211xp5_ASAP7_75t_R u0_g62690 (.A1(u0_n_32165),
    .A2(u0_n_31467),
    .B(u0_n_31232),
    .C(u0_n_31352),
    .Y(u0_n_30382));
 OR2x2_ASAP7_75t_R u0_g62691 (.A(u0_n_32845),
    .B(u0_n_30773),
    .Y(u0_n_30383));
 AOI32xp33_ASAP7_75t_SL u0_g62692 (.A1(u0_n_31685),
    .A2(u0_n_31799),
    .A3(n_8656),
    .B1(u0_n_31344),
    .B2(w3[19]),
    .Y(u0_n_30385));
 OAI321xp33_ASAP7_75t_L u0_g62693 (.A1(u0_n_31653),
    .A2(u0_n_32747),
    .A3(u0_n_32737),
    .B1(u0_n_31837),
    .B2(u0_n_31900),
    .C(u0_n_30833),
    .Y(u0_n_30388));
 AOI211xp5_ASAP7_75t_SL u0_g62694 (.A1(u0_n_31791),
    .A2(u0_n_32373),
    .B(u0_n_30779),
    .C(u0_n_31578),
    .Y(u0_n_30390));
 OAI21xp33_ASAP7_75t_L u0_g62695 (.A1(u0_n_32083),
    .A2(u0_n_31259),
    .B(u0_n_30935),
    .Y(u0_n_30391));
 AOI221xp5_ASAP7_75t_R u0_g62696 (.A1(u0_n_31484),
    .A2(u0_n_31841),
    .B1(u0_n_32142),
    .B2(u0_n_31795),
    .C(u0_n_31349),
    .Y(u0_n_30392));
 AOI211xp5_ASAP7_75t_L u0_g62697 (.A1(u0_n_31414),
    .A2(u0_n_32040),
    .B(u0_n_30950),
    .C(u0_n_31797),
    .Y(u0_n_30395));
 AOI21xp33_ASAP7_75t_R u0_g62698 (.A1(u0_n_31121),
    .A2(u0_n_31464),
    .B(u0_n_30931),
    .Y(u0_n_30396));
 AO21x1_ASAP7_75t_SL u0_g62699 (.A1(u0_n_32142),
    .A2(u0_n_31255),
    .B(u0_n_31231),
    .Y(u0_n_30398));
 AOI21xp5_ASAP7_75t_L u0_g62700 (.A1(u0_n_31251),
    .A2(u0_n_32407),
    .B(u0_n_31298),
    .Y(u0_n_30400));
 OAI21xp33_ASAP7_75t_R u0_g62701 (.A1(u0_n_32385),
    .A2(u0_n_31256),
    .B(u0_n_31296),
    .Y(u0_n_30402));
 NOR2xp33_ASAP7_75t_R u0_g62702 (.A(u0_n_31842),
    .B(u0_n_30748),
    .Y(u0_n_30404));
 OAI211xp5_ASAP7_75t_L u0_g62703 (.A1(u0_n_32121),
    .A2(u0_n_31433),
    .B(u0_n_30901),
    .C(u0_n_31784),
    .Y(u0_n_30405));
 OAI21xp33_ASAP7_75t_R u0_g62704 (.A1(u0_n_31507),
    .A2(u0_n_31182),
    .B(u0_n_32113),
    .Y(u0_n_30406));
 OAI21xp33_ASAP7_75t_R u0_g62705 (.A1(u0_n_31501),
    .A2(u0_n_31180),
    .B(u0_n_31998),
    .Y(u0_n_30408));
 AOI21xp33_ASAP7_75t_R u0_g62706 (.A1(u0_n_31187),
    .A2(u0_n_31504),
    .B(u0_n_32075),
    .Y(u0_n_30409));
 AOI21xp33_ASAP7_75t_R u0_g62707 (.A1(u0_n_31170),
    .A2(u0_n_31823),
    .B(u0_n_32385),
    .Y(u0_n_30411));
 AOI32xp33_ASAP7_75t_R u0_g62708 (.A1(u0_n_31689),
    .A2(u0_n_32073),
    .A3(u0_n_31795),
    .B1(u0_n_31191),
    .B2(u0_n_31874),
    .Y(u0_n_30413));
 OAI21xp33_ASAP7_75t_R u0_g62709 (.A1(u0_n_32209),
    .A2(u0_n_31257),
    .B(u0_n_30908),
    .Y(u0_n_30415));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62710 (.A1(w3[11]),
    .A2(u0_n_31582),
    .B(u0_n_31193),
    .C(n_8801),
    .Y(u0_n_30418));
 AOI211xp5_ASAP7_75t_R u0_g62711 (.A1(u0_n_31540),
    .A2(u0_n_32416),
    .B(u0_n_31238),
    .C(u0_n_31451),
    .Y(u0_n_30419));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62712 (.A1(u0_n_31503),
    .A2(u0_n_31688),
    .B(w3[3]),
    .C(u0_n_31030),
    .Y(u0_n_30420));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62713 (.A1(u0_n_31492),
    .A2(u0_n_31680),
    .B(\u0_w[3] [27]),
    .C(u0_n_31009),
    .Y(u0_n_30422));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62714 (.A1(u0_n_31686),
    .A2(u0_n_31507),
    .B(w3[11]),
    .C(u0_n_31021),
    .Y(u0_n_30423));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62715 (.A1(u0_n_31685),
    .A2(u0_n_31500),
    .B(n_8656),
    .C(u0_n_31017),
    .Y(u0_n_30425));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62716 (.A1(n_8831),
    .A2(u0_n_31800),
    .B(u0_n_32208),
    .C(u0_n_30912),
    .Y(u0_n_30427));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62717 (.A1(\u0_w[3] [27]),
    .A2(n_8946),
    .B(u0_n_31330),
    .C(u0_n_31769),
    .Y(u0_n_30428));
 OAI221xp5_ASAP7_75t_R u0_g62718 (.A1(u0_n_31413),
    .A2(u0_n_31477),
    .B1(u0_n_31671),
    .B2(u0_n_31438),
    .C(u0_n_31911),
    .Y(u0_n_30431));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62719 (.A1(w3[11]),
    .A2(u0_n_32759),
    .B(u0_n_31324),
    .C(u0_n_31762),
    .Y(u0_n_30435));
 AOI321xp33_ASAP7_75t_L u0_g62720 (.A1(u0_n_31665),
    .A2(n_11401),
    .A3(w3[11]),
    .B1(u0_n_31395),
    .B2(u0_n_31763),
    .C(u0_n_31624),
    .Y(u0_n_30438));
 NOR4xp25_ASAP7_75t_L u0_g62721 (.A(u0_n_30913),
    .B(u0_n_31656),
    .C(u0_n_31595),
    .D(w3[18]),
    .Y(u0_n_30441));
 AOI21xp33_ASAP7_75t_L u0_g62722 (.A1(u0_n_31135),
    .A2(u0_n_33033),
    .B(u0_n_30840),
    .Y(u0_n_30443));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62723 (.A1(n_8668),
    .A2(u0_n_33138),
    .B(u0_n_31329),
    .C(u0_n_31917),
    .Y(u0_n_30445));
 OAI321xp33_ASAP7_75t_R u0_g62724 (.A1(u0_n_31654),
    .A2(u0_n_32743),
    .A3(u0_n_32751),
    .B1(u0_n_31399),
    .B2(u0_n_31769),
    .C(u0_n_31621),
    .Y(u0_n_30449));
 OA211x2_ASAP7_75t_L u0_g62725 (.A1(n_8801),
    .A2(u0_n_31151),
    .B(u0_n_31358),
    .C(u0_n_31094),
    .Y(u0_n_30450));
 OAI211xp5_ASAP7_75t_L u0_g62726 (.A1(u0_n_31945),
    .A2(u0_n_31875),
    .B(u0_n_31640),
    .C(u0_n_31108),
    .Y(u0_n_30452));
 OAI221xp5_ASAP7_75t_R u0_g62727 (.A1(u0_n_32272),
    .A2(u0_n_31617),
    .B1(u0_n_31431),
    .B2(u0_n_32385),
    .C(u0_n_31090),
    .Y(u0_n_30453));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62728 (.A1(u0_n_32763),
    .A2(u0_n_31676),
    .B(u0_n_31895),
    .C(u0_n_30775),
    .Y(u0_n_30454));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62729 (.A1(w3[14]),
    .A2(u0_n_31674),
    .B(u0_n_32353),
    .C(u0_n_30758),
    .Y(u0_n_30457));
 AOI211xp5_ASAP7_75t_SL u0_g62730 (.A1(u0_n_31874),
    .A2(w3[7]),
    .B(u0_n_31242),
    .C(u0_n_31639),
    .Y(u0_n_30459));
 NAND3xp33_ASAP7_75t_R u0_g62731 (.A(u0_n_31099),
    .B(u0_n_31657),
    .C(u0_n_31596),
    .Y(u0_n_30460));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62732 (.A1(u0_n_33033),
    .A2(u0_n_31670),
    .B(u0_n_32273),
    .C(u0_n_30755),
    .Y(u0_n_30461));
 OAI211xp5_ASAP7_75t_SL u0_g62733 (.A1(u0_n_32385),
    .A2(u0_n_31485),
    .B(u0_n_30918),
    .C(u0_n_31643),
    .Y(u0_n_30463));
 OAI31xp33_ASAP7_75t_R u0_g62734 (.A1(u0_n_31140),
    .A2(u0_n_31820),
    .A3(n_11371),
    .B(u0_n_32241),
    .Y(u0_n_30464));
 AOI32xp33_ASAP7_75t_R u0_g62735 (.A1(u0_n_31681),
    .A2(u0_n_32052),
    .A3(u0_n_31791),
    .B1(u0_n_31190),
    .B2(u0_n_32289),
    .Y(u0_n_30465));
 AOI311xp33_ASAP7_75t_L u0_g62736 (.A1(u0_n_31850),
    .A2(u0_n_31839),
    .A3(n_8625),
    .B(u0_n_30949),
    .C(u0_n_31252),
    .Y(u0_n_30467));
 OAI21xp33_ASAP7_75t_L u0_g62737 (.A1(u0_n_31988),
    .A2(u0_n_31290),
    .B(\u0_w[3] [16]),
    .Y(u0_n_30469));
 OA21x2_ASAP7_75t_R u0_g62738 (.A1(u0_n_32083),
    .A2(u0_n_31268),
    .B(w3[0]),
    .Y(u0_n_30471));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62739 (.A1(u0_n_31817),
    .A2(u0_n_31541),
    .B(u0_n_32109),
    .C(n_11401),
    .Y(u0_n_30472));
 OAI21xp33_ASAP7_75t_R u0_g62740 (.A1(u0_n_31276),
    .A2(u0_n_32774),
    .B(u0_n_32141),
    .Y(u0_n_30474));
 AOI31xp33_ASAP7_75t_SL u0_g62741 (.A1(u0_n_31814),
    .A2(u0_n_32339),
    .A3(n_11401),
    .B(u0_n_30825),
    .Y(u0_n_30476));
 AOI21xp33_ASAP7_75t_R u0_g62742 (.A1(u0_n_31151),
    .A2(u0_n_32184),
    .B(u0_n_31778),
    .Y(u0_n_30477));
 OA21x2_ASAP7_75t_R u0_g62743 (.A1(n_8820),
    .A2(u0_n_31286),
    .B(u0_n_32425),
    .Y(u0_n_30478));
 AO21x1_ASAP7_75t_R u0_g62744 (.A1(u0_n_32795),
    .A2(u0_n_31294),
    .B(u0_n_32248),
    .Y(u0_n_30480));
 AO21x1_ASAP7_75t_R u0_g62745 (.A1(u0_n_32793),
    .A2(u0_n_31275),
    .B(u0_n_32373),
    .Y(u0_n_30482));
 AOI321xp33_ASAP7_75t_L u0_g62746 (.A1(u0_n_32080),
    .A2(w3[0]),
    .A3(n_8629),
    .B1(u0_n_31443),
    .B2(u0_n_31676),
    .C(u0_n_31913),
    .Y(u0_n_30484));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62747 (.A1(u0_n_31837),
    .A2(u0_n_31547),
    .B(u0_n_32083),
    .C(u0_n_32747),
    .Y(u0_n_30486));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62748 (.A1(u0_n_31830),
    .A2(u0_n_31549),
    .B(u0_n_32053),
    .C(u0_n_32743),
    .Y(u0_n_30488));
 OAI211xp5_ASAP7_75t_L u0_g62749 (.A1(u0_n_32075),
    .A2(u0_n_31546),
    .B(u0_n_30747),
    .C(u0_n_31592),
    .Y(u0_n_30489));
 OAI211xp5_ASAP7_75t_R u0_g62750 (.A1(u0_n_32209),
    .A2(u0_n_31638),
    .B(u0_n_31261),
    .C(u0_n_31957),
    .Y(u0_n_30491));
 OAI21xp33_ASAP7_75t_L u0_g62751 (.A1(u0_n_32042),
    .A2(u0_n_31330),
    .B(u0_n_31040),
    .Y(u0_n_30492));
 O2A1O1Ixp33_ASAP7_75t_L u0_g62752 (.A1(w3[3]),
    .A2(n_8625),
    .B(u0_n_31301),
    .C(u0_n_32774),
    .Y(u0_n_30493));
 AND3x1_ASAP7_75t_R u0_g62753 (.A(u0_n_31260),
    .B(u0_n_31085),
    .C(u0_n_31520),
    .Y(u0_n_30495));
 AOI21xp33_ASAP7_75t_R u0_g62754 (.A1(u0_n_31263),
    .A2(u0_n_32113),
    .B(u0_n_30746),
    .Y(u0_n_30498));
 AOI21xp33_ASAP7_75t_R u0_g62755 (.A1(u0_n_31163),
    .A2(u0_n_31840),
    .B(u0_n_32141),
    .Y(u0_n_30501));
 OAI221xp5_ASAP7_75t_L u0_g62756 (.A1(u0_n_31607),
    .A2(u0_n_32321),
    .B1(u0_n_32053),
    .B2(u0_n_31972),
    .C(u0_n_31048),
    .Y(u0_n_30503));
 AO21x1_ASAP7_75t_R u0_g62757 (.A1(u0_n_31830),
    .A2(u0_n_31170),
    .B(u0_n_32306),
    .Y(u0_n_30504));
 NOR2xp33_ASAP7_75t_L u0_g62758 (.A(u0_n_32141),
    .B(u0_n_30749),
    .Y(u0_n_30348));
 AOI21xp33_ASAP7_75t_R u0_g62759 (.A1(u0_n_31840),
    .A2(u0_n_31187),
    .B(u0_n_32141),
    .Y(u0_n_30349));
 AOI21xp5_ASAP7_75t_L u0_g62760 (.A1(u0_n_31184),
    .A2(u0_n_31823),
    .B(u0_n_32372),
    .Y(u0_n_30350));
 AOI21xp33_ASAP7_75t_R u0_g62761 (.A1(u0_n_31819),
    .A2(u0_n_31181),
    .B(u0_n_32254),
    .Y(u0_n_30351));
 NOR2xp33_ASAP7_75t_R u0_g62763 (.A(u0_n_30725),
    .B(u0_n_30773),
    .Y(u0_n_30506));
 NAND2xp33_ASAP7_75t_SL u0_g62764 (.A(u0_n_30770),
    .B(u0_n_32308),
    .Y(u0_n_30352));
 NOR2xp33_ASAP7_75t_SL u0_g62765 (.A(u0_n_32763),
    .B(u0_n_30775),
    .Y(u0_n_30353));
 NOR2xp33_ASAP7_75t_L u0_g62766 (.A(u0_n_32254),
    .B(u0_n_30751),
    .Y(u0_n_30354));
 OR2x2_ASAP7_75t_SL u0_g62767 (.A(u0_n_32409),
    .B(u0_n_30750),
    .Y(u0_n_30355));
 NOR2xp33_ASAP7_75t_R u0_g62768 (.A(u0_n_32194),
    .B(u0_n_30753),
    .Y(u0_n_30356));
 OR2x2_ASAP7_75t_L u0_g62769 (.A(u0_n_31842),
    .B(u0_n_30761),
    .Y(u0_n_30357));
 OAI21xp33_ASAP7_75t_R u0_g62770 (.A1(u0_n_31825),
    .A2(u0_n_31182),
    .B(u0_n_32416),
    .Y(u0_n_30358));
 NAND2xp33_ASAP7_75t_R u0_g62771 (.A(u0_n_30759),
    .B(n_8801),
    .Y(u0_n_30359));
 AND2x2_ASAP7_75t_L u0_g62772 (.A(u0_n_33004),
    .B(u0_n_30754),
    .Y(u0_n_30360));
 NOR2xp33_ASAP7_75t_SL u0_g62773 (.A(u0_n_32793),
    .B(u0_n_30755),
    .Y(u0_n_30362));
 NAND2xp5_ASAP7_75t_L u0_g62774 (.A(u0_n_30759),
    .B(n_8820),
    .Y(u0_n_30364));
 NOR2xp33_ASAP7_75t_R u0_g62775 (.A(u0_n_33033),
    .B(u0_n_30755),
    .Y(u0_n_30514));
 NAND2xp33_ASAP7_75t_R u0_g62776 (.A(u0_n_32795),
    .B(u0_n_30754),
    .Y(u0_n_30366));
 NOR2xp33_ASAP7_75t_SL u0_g62777 (.A(u0_n_30767),
    .B(u0_n_30722),
    .Y(u0_n_30367));
 NAND2xp5_ASAP7_75t_L u0_g62778 (.A(u0_n_30738),
    .B(u0_n_32339),
    .Y(u0_n_30368));
 NOR2xp33_ASAP7_75t_R u0_g62779 (.A(u0_r0_rcnt[0]),
    .B(u0_n_30774),
    .Y(u0_n_30369));
 OR2x2_ASAP7_75t_SL u0_g62780 (.A(u0_n_30726),
    .B(u0_n_30768),
    .Y(u0_n_30370));
 NAND2xp5_ASAP7_75t_L u0_g62781 (.A(u0_n_32226),
    .B(u0_n_30736),
    .Y(u0_n_30372));
 AND2x2_ASAP7_75t_R u0_g62782 (.A(u0_r0_rcnt[0]),
    .B(u0_n_30773),
    .Y(u0_n_30373));
 INVx1_ASAP7_75t_SL u0_g62783 (.A(u0_n_30635),
    .Y(u0_n_30520));
 INVxp67_ASAP7_75t_L u0_g62784 (.A(u0_n_30700),
    .Y(u0_n_30521));
 AOI22xp33_ASAP7_75t_SL u0_g62785 (.A1(u0_n_31081),
    .A2(u0_n_31160),
    .B1(u0_n_31489),
    .B2(u0_n_31129),
    .Y(u0_n_30522));
 OAI221xp5_ASAP7_75t_L u0_g62786 (.A1(u0_n_31610),
    .A2(u0_n_32194),
    .B1(u0_n_31622),
    .B2(u0_n_32338),
    .C(u0_n_31055),
    .Y(u0_n_30524));
 AOI211xp5_ASAP7_75t_SL u0_g62787 (.A1(u0_n_31470),
    .A2(u0_n_32184),
    .B(u0_n_31356),
    .C(u0_n_31624),
    .Y(u0_n_30525));
 OAI21xp33_ASAP7_75t_R u0_g62788 (.A1(u0_n_31800),
    .A2(u0_n_31244),
    .B(u0_n_30987),
    .Y(u0_n_30527));
 OAI221xp5_ASAP7_75t_L u0_g62789 (.A1(u0_n_31445),
    .A2(u0_n_32242),
    .B1(u0_n_32221),
    .B2(u0_n_31919),
    .C(u0_n_30861),
    .Y(u0_n_30529));
 NOR3xp33_ASAP7_75t_R u0_g62790 (.A(u0_n_30956),
    .B(u0_n_31337),
    .C(u0_n_31789),
    .Y(u0_n_30530));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62791 (.A1(u0_n_31800),
    .A2(u0_n_31542),
    .B(u0_n_32248),
    .C(u0_n_31690),
    .Y(u0_n_30531));
 OAI211xp5_ASAP7_75t_SL u0_g62792 (.A1(u0_n_31846),
    .A2(u0_n_31266),
    .B(u0_n_31082),
    .C(u0_n_31361),
    .Y(u0_n_30532));
 OAI21xp33_ASAP7_75t_R u0_g62793 (.A1(u0_n_32017),
    .A2(u0_n_31317),
    .B(u0_n_30934),
    .Y(u0_n_30535));
 OAI221xp5_ASAP7_75t_L u0_g62794 (.A1(u0_n_31599),
    .A2(u0_n_32194),
    .B1(u0_n_32410),
    .B2(u0_n_31929),
    .C(u0_n_30902),
    .Y(u0_n_30536));
 OAI22xp33_ASAP7_75t_R u0_g62795 (.A1(u0_n_32075),
    .A2(u0_n_31202),
    .B1(u0_n_31842),
    .B2(u0_n_31314),
    .Y(u0_n_30538));
 OAI221xp5_ASAP7_75t_R u0_g62796 (.A1(u0_n_31648),
    .A2(u0_n_31842),
    .B1(u0_n_31625),
    .B2(u0_n_31886),
    .C(u0_n_31053),
    .Y(u0_n_30540));
 OAI21xp33_ASAP7_75t_L u0_g62797 (.A1(u0_n_32306),
    .A2(u0_n_31277),
    .B(u0_n_30943),
    .Y(u0_n_30541));
 OAI21xp33_ASAP7_75t_R u0_g62798 (.A1(u0_n_31830),
    .A2(u0_n_32304),
    .B(u0_n_30936),
    .Y(u0_n_30542));
 OAI21xp33_ASAP7_75t_R u0_g62799 (.A1(u0_n_32321),
    .A2(u0_n_31318),
    .B(u0_n_30817),
    .Y(u0_n_30543));
 OAI221xp5_ASAP7_75t_SL u0_g62800 (.A1(u0_n_31598),
    .A2(u0_n_32321),
    .B1(u0_n_31607),
    .B2(u0_n_32290),
    .C(u0_n_31028),
    .Y(u0_n_30544));
 OAI221xp5_ASAP7_75t_L u0_g62801 (.A1(u0_n_31276),
    .A2(u0_n_31459),
    .B1(u0_n_31531),
    .B2(u0_n_31766),
    .C(u0_n_31756),
    .Y(u0_n_30546));
 OAI211xp5_ASAP7_75t_L u0_g62802 (.A1(u0_n_32053),
    .A2(u0_n_31323),
    .B(u0_n_31112),
    .C(u0_n_31253),
    .Y(u0_n_30549));
 OAI21xp33_ASAP7_75t_R u0_g62803 (.A1(u0_n_32042),
    .A2(u0_n_31275),
    .B(u0_n_31012),
    .Y(u0_n_30550));
 OAI221xp5_ASAP7_75t_L u0_g62804 (.A1(u0_n_32338),
    .A2(u0_n_31418),
    .B1(u0_n_32185),
    .B2(u0_n_31970),
    .C(u0_n_30871),
    .Y(u0_n_30551));
 OAI21xp33_ASAP7_75t_R u0_g62805 (.A1(u0_n_32221),
    .A2(u0_n_31130),
    .B(u0_n_31026),
    .Y(u0_n_30553));
 AOI221xp5_ASAP7_75t_R u0_g62806 (.A1(u0_n_32142),
    .A2(u0_n_31499),
    .B1(u0_n_31850),
    .B2(w3[7]),
    .C(u0_n_30867),
    .Y(u0_n_30555));
 AOI221xp5_ASAP7_75t_SL u0_g62807 (.A1(u0_n_31449),
    .A2(u0_n_32386),
    .B1(u0_n_32320),
    .B2(u0_n_32717),
    .C(u0_n_30859),
    .Y(u0_n_30557));
 OAI221xp5_ASAP7_75t_SL u0_g62808 (.A1(u0_n_32410),
    .A2(u0_n_31473),
    .B1(u0_n_32194),
    .B2(u0_n_32714),
    .C(u0_n_30857),
    .Y(u0_n_30558));
 OAI22xp33_ASAP7_75t_L u0_g62809 (.A1(u0_n_31423),
    .A2(u0_n_31314),
    .B1(u0_n_31815),
    .B2(u0_n_32141),
    .Y(u0_n_30560));
 OAI222xp33_ASAP7_75t_R u0_g62810 (.A1(u0_n_31464),
    .A2(u0_n_32763),
    .B1(u0_n_31461),
    .B2(n_11457),
    .C1(u0_n_32165),
    .C2(u0_n_31963),
    .Y(u0_n_30561));
 AOI222xp33_ASAP7_75t_R u0_g62811 (.A1(u0_n_31181),
    .A2(u0_n_32241),
    .B1(u0_n_33001),
    .B2(u0_n_31627),
    .C1(u0_n_32226),
    .C2(u0_n_31965),
    .Y(u0_n_30563));
 AOI222xp33_ASAP7_75t_R u0_g62812 (.A1(u0_n_31184),
    .A2(u0_n_32386),
    .B1(u0_n_31628),
    .B2(u0_n_33033),
    .C1(u0_n_32289),
    .C2(u0_n_31959),
    .Y(u0_n_30565));
 OAI222xp33_ASAP7_75t_R u0_g62813 (.A1(u0_n_31623),
    .A2(n_8801),
    .B1(u0_n_31182),
    .B2(u0_n_32425),
    .C1(u0_n_32338),
    .C2(u0_n_31969),
    .Y(u0_n_30567));
 AOI21xp33_ASAP7_75t_R u0_g62814 (.A1(u0_n_32166),
    .A2(u0_n_31187),
    .B(u0_n_31056),
    .Y(u0_n_30569));
 AOI22xp33_ASAP7_75t_R u0_g62815 (.A1(u0_n_32737),
    .A2(u0_n_31126),
    .B1(w3[3]),
    .B2(u0_n_31127),
    .Y(u0_n_30570));
 AOI222xp33_ASAP7_75t_SL u0_g62816 (.A1(u0_n_31585),
    .A2(u0_n_32763),
    .B1(u0_n_31874),
    .B2(u0_n_31977),
    .C1(u0_n_31614),
    .C2(u0_n_32142),
    .Y(u0_n_30572));
 AOI222xp33_ASAP7_75t_R u0_g62817 (.A1(u0_n_31638),
    .A2(n_8656),
    .B1(u0_n_32241),
    .B2(u0_n_31966),
    .C1(u0_n_31545),
    .C2(w3[19]),
    .Y(u0_n_30573));
 OAI222xp33_ASAP7_75t_R u0_g62818 (.A1(u0_n_31498),
    .A2(u0_n_33033),
    .B1(u0_n_31482),
    .B2(\u0_w[3] [27]),
    .C1(u0_n_32372),
    .C2(u0_n_31959),
    .Y(u0_n_30575));
 OAI21xp33_ASAP7_75t_R u0_g62819 (.A1(u0_n_32011),
    .A2(u0_n_31130),
    .B(u0_n_31051),
    .Y(u0_n_30576));
 OAI221xp5_ASAP7_75t_R u0_g62820 (.A1(u0_n_32344),
    .A2(u0_n_31568),
    .B1(u0_n_32425),
    .B2(n_8856),
    .C(u0_n_31339),
    .Y(u0_n_30577));
 OAI221xp5_ASAP7_75t_R u0_g62821 (.A1(u0_n_31433),
    .A2(u0_n_31474),
    .B1(u0_n_31441),
    .B2(u0_n_31675),
    .C(u0_n_31915),
    .Y(u0_n_30578));
 OAI222xp33_ASAP7_75t_R u0_g62822 (.A1(u0_n_32290),
    .A2(u0_n_31659),
    .B1(u0_n_31519),
    .B2(u0_n_32321),
    .C1(u0_n_32372),
    .C2(u0_n_31781),
    .Y(u0_n_30582));
 OAI221xp5_ASAP7_75t_R u0_g62823 (.A1(u0_n_31322),
    .A2(u0_n_32409),
    .B1(u0_n_32174),
    .B2(u0_n_31928),
    .C(u0_n_31933),
    .Y(u0_n_30584));
 OAI321xp33_ASAP7_75t_L u0_g62824 (.A1(u0_n_32753),
    .A2(u0_n_31807),
    .A3(u0_n_32209),
    .B1(u0_n_31293),
    .B2(u0_n_31468),
    .C(u0_n_31760),
    .Y(u0_n_30586));
 AOI322xp5_ASAP7_75t_R u0_g62825 (.A1(u0_n_31538),
    .A2(u0_n_32193),
    .A3(u0_n_31927),
    .B1(w3[14]),
    .B2(u0_n_31169),
    .C1(u0_n_32122),
    .C2(w3[15]),
    .Y(u0_n_30589));
 AOI22xp33_ASAP7_75t_R u0_g62826 (.A1(u0_n_31325),
    .A2(u0_n_32122),
    .B1(u0_n_31322),
    .B2(u0_n_32407),
    .Y(u0_n_30591));
 AOI221xp5_ASAP7_75t_R u0_g62827 (.A1(u0_n_31573),
    .A2(u0_n_32289),
    .B1(u0_n_32320),
    .B2(u0_n_31498),
    .C(u0_n_31401),
    .Y(u0_n_30592));
 OAI221xp5_ASAP7_75t_R u0_g62828 (.A1(u0_n_31137),
    .A2(u0_n_32372),
    .B1(u0_n_31429),
    .B2(u0_n_32793),
    .C(u0_n_31396),
    .Y(u0_n_30594));
 OAI221xp5_ASAP7_75t_SL u0_g62829 (.A1(u0_n_32272),
    .A2(u0_n_31309),
    .B1(u0_n_31576),
    .B2(u0_n_32372),
    .C(u0_n_31090),
    .Y(u0_n_30595));
 AOI211xp5_ASAP7_75t_R u0_g62830 (.A1(u0_n_31265),
    .A2(u0_n_32021),
    .B(u0_n_31588),
    .C(u0_n_31402),
    .Y(u0_n_30597));
 AOI221xp5_ASAP7_75t_R u0_g62831 (.A1(u0_n_31462),
    .A2(u0_n_33001),
    .B1(u0_n_31165),
    .B2(u0_n_32248),
    .C(u0_n_31394),
    .Y(u0_n_30598));
 OAI221xp5_ASAP7_75t_R u0_g62832 (.A1(u0_n_31306),
    .A2(u0_n_32221),
    .B1(u0_n_31593),
    .B2(u0_n_31984),
    .C(u0_n_31092),
    .Y(u0_n_30599));
 OAI221xp5_ASAP7_75t_L u0_g62833 (.A1(u0_n_31886),
    .A2(u0_n_31648),
    .B1(u0_n_31461),
    .B2(u0_n_32075),
    .C(u0_n_30946),
    .Y(u0_n_30602));
 OAI322xp33_ASAP7_75t_R u0_g62834 (.A1(u0_n_31682),
    .A2(u0_n_32321),
    .A3(u0_n_31930),
    .B1(u0_n_31122),
    .B2(u0_n_32793),
    .C1(u0_n_32053),
    .C2(u0_n_32716),
    .Y(u0_n_30605));
 AOI22xp33_ASAP7_75t_L u0_g62835 (.A1(u0_n_31442),
    .A2(u0_n_31168),
    .B1(u0_n_31794),
    .B2(u0_n_31475),
    .Y(u0_n_30606));
 AOI22xp33_ASAP7_75t_R u0_g62836 (.A1(u0_n_31167),
    .A2(u0_n_31435),
    .B1(u0_n_31469),
    .B2(u0_n_31800),
    .Y(u0_n_30608));
 AOI322xp5_ASAP7_75t_L u0_g62837 (.A1(u0_n_31178),
    .A2(u0_n_31609),
    .A3(u0_n_32795),
    .B1(u0_n_31998),
    .B2(u0_n_31620),
    .C1(u0_n_32021),
    .C2(u0_n_31961),
    .Y(u0_n_30611));
 OAI322xp33_ASAP7_75t_L u0_g62838 (.A1(u0_n_31173),
    .A2(u0_n_31618),
    .A3(u0_n_33033),
    .B1(u0_n_31597),
    .B2(u0_n_32053),
    .C1(u0_n_32315),
    .C2(u0_n_31944),
    .Y(u0_n_30614));
 AOI321xp33_ASAP7_75t_R u0_g62839 (.A1(u0_n_31508),
    .A2(u0_n_31687),
    .A3(u0_n_32122),
    .B1(u0_n_32339),
    .B2(u0_n_31927),
    .C(u0_n_31636),
    .Y(u0_n_30615));
 OAI321xp33_ASAP7_75t_R u0_g62840 (.A1(u0_n_31680),
    .A2(u0_n_31492),
    .A3(u0_n_32042),
    .B1(u0_n_31930),
    .B2(u0_n_32272),
    .C(u0_n_31635),
    .Y(u0_n_30618));
 OAI321xp33_ASAP7_75t_R u0_g62841 (.A1(u0_n_31501),
    .A2(u0_n_31684),
    .A3(u0_n_31988),
    .B1(u0_n_31918),
    .B2(u0_n_32221),
    .C(u0_n_31632),
    .Y(u0_n_30623));
 OAI321xp33_ASAP7_75t_R u0_g62842 (.A1(u0_n_31688),
    .A2(u0_n_32075),
    .A3(u0_n_31503),
    .B1(u0_n_31924),
    .B2(u0_n_31875),
    .C(u0_n_31633),
    .Y(u0_n_30626));
 OAI322xp33_ASAP7_75t_R u0_g62843 (.A1(u0_n_31661),
    .A2(u0_n_31522),
    .A3(u0_n_31988),
    .B1(u0_n_31463),
    .B2(n_8656),
    .C1(u0_n_32209),
    .C2(w3[20]),
    .Y(u0_n_30629));
 OAI22xp5_ASAP7_75t_L u0_g62844 (.A1(u0_n_31649),
    .A2(u0_n_31131),
    .B1(u0_n_31614),
    .B2(u0_n_31139),
    .Y(u0_n_30632));
 OAI22xp5_ASAP7_75t_L u0_g62845 (.A1(u0_n_31164),
    .A2(u0_n_31159),
    .B1(u0_n_31820),
    .B2(u0_n_31128),
    .Y(u0_n_30635));
 OAI322xp33_ASAP7_75t_SL u0_g62846 (.A1(u0_n_31518),
    .A2(u0_n_31654),
    .A3(u0_n_32042),
    .B1(u0_n_32751),
    .B2(u0_n_31429),
    .C1(u0_n_32290),
    .C2(w3[28]),
    .Y(u0_n_30640));
 OAI322xp33_ASAP7_75t_R u0_g62847 (.A1(u0_n_32254),
    .A2(u0_n_31984),
    .A3(w3[17]),
    .B1(u0_n_31627),
    .B2(u0_n_32221),
    .C1(u0_n_31988),
    .C2(u0_n_31953),
    .Y(u0_n_30644));
 OA21x2_ASAP7_75t_SL u0_g62848 (.A1(u0_n_31650),
    .A2(u0_n_31147),
    .B(u0_n_30873),
    .Y(u0_n_30647));
 AOI211xp5_ASAP7_75t_R u0_g62849 (.A1(u0_n_31168),
    .A2(u0_n_32113),
    .B(u0_n_31084),
    .C(u0_n_31245),
    .Y(u0_n_30648));
 AOI22xp33_ASAP7_75t_R u0_g62850 (.A1(u0_n_31154),
    .A2(u0_n_31138),
    .B1(u0_n_31840),
    .B2(u0_n_31121),
    .Y(u0_n_30650));
 OAI22xp33_ASAP7_75t_R u0_g62851 (.A1(u0_n_31107),
    .A2(u0_n_32174),
    .B1(u0_n_31303),
    .B2(u0_n_32409),
    .Y(u0_n_30652));
 AOI221xp5_ASAP7_75t_R u0_g62852 (.A1(u0_n_32113),
    .A2(u0_n_32714),
    .B1(u0_n_31284),
    .B2(u0_n_32184),
    .C(u0_n_31591),
    .Y(u0_n_30653));
 OAI211xp5_ASAP7_75t_R u0_g62853 (.A1(u0_n_31875),
    .A2(u0_n_31105),
    .B(u0_n_31592),
    .C(u0_n_31942),
    .Y(u0_n_30654));
 AOI22xp33_ASAP7_75t_R u0_g62854 (.A1(u0_n_31874),
    .A2(u0_n_31146),
    .B1(u0_n_32080),
    .B2(u0_n_31570),
    .Y(u0_n_30658));
 OAI32xp33_ASAP7_75t_R u0_g62855 (.A1(u0_n_31140),
    .A2(u0_n_31542),
    .A3(u0_n_32017),
    .B1(u0_n_32242),
    .B2(u0_n_31250),
    .Y(u0_n_30659));
 AOI221xp5_ASAP7_75t_R u0_g62856 (.A1(u0_n_31113),
    .A2(u0_n_32273),
    .B1(u0_n_32308),
    .B2(u0_n_31923),
    .C(u0_n_31939),
    .Y(u0_n_30663));
 AOI322xp5_ASAP7_75t_SL u0_g62857 (.A1(u0_n_31176),
    .A2(u0_n_31604),
    .A3(n_8801),
    .B1(u0_n_32122),
    .B2(u0_n_31599),
    .C1(u0_n_32193),
    .C2(u0_n_31938),
    .Y(u0_n_30667));
 AOI221xp5_ASAP7_75t_R u0_g62858 (.A1(u0_n_31280),
    .A2(u0_n_32304),
    .B1(u0_n_32052),
    .B2(u0_n_32716),
    .C(u0_n_31584),
    .Y(u0_n_30668));
 OAI221xp5_ASAP7_75t_R u0_g62859 (.A1(u0_n_31104),
    .A2(u0_n_32221),
    .B1(u0_n_32023),
    .B2(u0_n_31935),
    .C(u0_n_31950),
    .Y(u0_n_30670));
 AOI322xp5_ASAP7_75t_L u0_g62860 (.A1(u0_n_31174),
    .A2(u0_n_31615),
    .A3(u0_n_32766),
    .B1(u0_n_32073),
    .B2(u0_n_31603),
    .C1(u0_n_31841),
    .C2(u0_n_31945),
    .Y(u0_n_30672));
 AOI321xp33_ASAP7_75t_R u0_g62861 (.A1(u0_n_31895),
    .A2(u0_n_31815),
    .A3(w3[7]),
    .B1(u0_n_31326),
    .B2(u0_n_32084),
    .C(u0_n_31780),
    .Y(u0_n_30674));
 AOI22xp33_ASAP7_75t_L u0_g62862 (.A1(u0_n_31439),
    .A2(u0_n_31122),
    .B1(u0_n_31792),
    .B2(u0_n_31478),
    .Y(u0_n_30676));
 AOI221xp5_ASAP7_75t_R u0_g62863 (.A1(u0_n_31465),
    .A2(u0_n_31986),
    .B1(u0_n_31288),
    .B2(u0_n_32226),
    .C(u0_n_31787),
    .Y(u0_n_30679));
 AOI22xp33_ASAP7_75t_L u0_g62864 (.A1(u0_n_31443),
    .A2(u0_n_31132),
    .B1(u0_n_31796),
    .B2(u0_n_31460),
    .Y(u0_n_30680));
 AOI22xp33_ASAP7_75t_R u0_g62865 (.A1(u0_n_32353),
    .A2(u0_n_31156),
    .B1(u0_n_31826),
    .B2(u0_n_32175),
    .Y(u0_n_30683));
 AOI21xp5_ASAP7_75t_R u0_g62866 (.A1(u0_n_31177),
    .A2(u0_n_32339),
    .B(u0_n_30994),
    .Y(u0_n_30685));
 AOI221xp5_ASAP7_75t_R u0_g62867 (.A1(u0_n_32073),
    .A2(u0_n_32697),
    .B1(u0_n_31126),
    .B2(u0_n_31850),
    .C(u0_n_31587),
    .Y(u0_n_30686));
 AOI22xp33_ASAP7_75t_R u0_g62868 (.A1(u0_n_31135),
    .A2(u0_n_32289),
    .B1(u0_n_31597),
    .B2(u0_n_32040),
    .Y(u0_n_30688));
 AOI22xp33_ASAP7_75t_R u0_g62869 (.A1(u0_n_32320),
    .A2(u0_n_31134),
    .B1(u0_n_31824),
    .B2(u0_n_32040),
    .Y(u0_n_30690));
 OAI221xp5_ASAP7_75t_L u0_g62870 (.A1(u0_n_31305),
    .A2(u0_n_32338),
    .B1(u0_n_31575),
    .B2(u0_n_32425),
    .C(u0_n_31118),
    .Y(u0_n_30692));
 AO22x1_ASAP7_75t_R u0_g62871 (.A1(u0_n_32175),
    .A2(u0_n_31142),
    .B1(u0_n_31825),
    .B2(u0_n_32109),
    .Y(u0_n_30695));
 AOI22xp33_ASAP7_75t_R u0_g62872 (.A1(u0_n_32084),
    .A2(u0_n_31235),
    .B1(u0_n_31874),
    .B2(u0_n_31533),
    .Y(u0_n_30697));
 OAI22xp33_ASAP7_75t_R u0_g62873 (.A1(u0_n_31842),
    .A2(u0_n_31136),
    .B1(u0_n_31840),
    .B2(u0_n_32075),
    .Y(u0_n_30698));
 AOI211xp5_ASAP7_75t_SL u0_g62874 (.A1(u0_n_31167),
    .A2(u0_n_31986),
    .B(u0_n_31248),
    .C(u0_n_31115),
    .Y(u0_n_30700));
 OAI221xp5_ASAP7_75t_R u0_g62875 (.A1(u0_n_31155),
    .A2(u0_n_32141),
    .B1(u0_n_31645),
    .B2(u0_n_32773),
    .C(u0_n_31388),
    .Y(u0_n_30702));
 AOI221xp5_ASAP7_75t_L u0_g62876 (.A1(u0_n_31630),
    .A2(n_8820),
    .B1(u0_n_31156),
    .B2(u0_n_32416),
    .C(u0_n_31398),
    .Y(u0_n_30704));
 AOI221xp5_ASAP7_75t_R u0_g62877 (.A1(u0_n_31301),
    .A2(u0_n_32073),
    .B1(u0_n_31570),
    .B2(u0_n_32773),
    .C(u0_n_31249),
    .Y(u0_n_30705));
 AOI221xp5_ASAP7_75t_SL u0_g62878 (.A1(u0_n_31307),
    .A2(u0_n_31986),
    .B1(u0_n_31391),
    .B2(u0_n_32795),
    .C(u0_n_31248),
    .Y(u0_n_30708));
 AO221x1_ASAP7_75t_L u0_g62879 (.A1(u0_n_31310),
    .A2(u0_n_32063),
    .B1(u0_n_31569),
    .B2(u0_n_32793),
    .C(u0_n_31247),
    .Y(u0_n_30711));
 AOI22xp33_ASAP7_75t_R u0_g62880 (.A1(u0_n_31986),
    .A2(u0_n_31282),
    .B1(u0_n_32260),
    .B2(u0_n_31545),
    .Y(u0_n_30715));
 INVxp67_ASAP7_75t_R u0_g62881 (.A(u0_n_30720),
    .Y(u0_n_30719));
 INVxp67_ASAP7_75t_R u0_g62882 (.A(u0_n_30724),
    .Y(u0_n_30723));
 INVxp33_ASAP7_75t_R u0_g62883 (.A(u0_n_30730),
    .Y(u0_n_30729));
 INVxp67_ASAP7_75t_R u0_g62884 (.A(u0_n_30743),
    .Y(u0_n_30742));
 INVxp33_ASAP7_75t_R u0_g62885 (.A(u0_n_30749),
    .Y(u0_n_30748));
 INVxp33_ASAP7_75t_R u0_g62886 (.A(u0_n_30753),
    .Y(u0_n_30752));
 INVxp67_ASAP7_75t_R u0_g62887 (.A(u0_n_30757),
    .Y(u0_n_30756));
 INVxp33_ASAP7_75t_R u0_g62888 (.A(u0_n_30759),
    .Y(u0_n_30758));
 INVxp33_ASAP7_75t_R u0_g62889 (.A(u0_n_30763),
    .Y(u0_n_30764));
 INVxp67_ASAP7_75t_R u0_g62890 (.A(u0_n_30767),
    .Y(u0_n_30766));
 INVxp33_ASAP7_75t_R u0_g62891 (.A(u0_n_30770),
    .Y(u0_n_30769));
 INVxp67_ASAP7_75t_L u0_g62892 (.A(u0_n_30771),
    .Y(u0_n_30772));
 INVxp33_ASAP7_75t_R u0_g62893 (.A(u0_n_30773),
    .Y(u0_n_30774));
 INVxp33_ASAP7_75t_R u0_g62894 (.A(u0_n_30775),
    .Y(u0_n_30776));
 NOR2xp33_ASAP7_75t_R u0_g62895 (.A(u0_n_31841),
    .B(u0_n_31327),
    .Y(u0_n_30777));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62896 (.A1(u0_n_32793),
    .A2(u0_n_31803),
    .B(u0_n_32272),
    .C(u0_n_31497),
    .Y(u0_n_30778));
 OAI21xp33_ASAP7_75t_L u0_g62897 (.A1(u0_n_32306),
    .A2(u0_n_31651),
    .B(u0_n_31621),
    .Y(u0_n_30779));
 AOI211xp5_ASAP7_75t_R u0_g62898 (.A1(u0_n_32273),
    .A2(u0_n_31972),
    .B(u0_n_31680),
    .C(u0_n_32743),
    .Y(u0_n_30782));
 NOR2xp33_ASAP7_75t_R u0_g62899 (.A(u0_n_31336),
    .B(u0_n_31313),
    .Y(u0_n_30784));
 NAND2xp33_ASAP7_75t_R u0_g62900 (.A(u0_n_32839),
    .B(u0_n_31333),
    .Y(u0_n_30785));
 OAI211xp5_ASAP7_75t_R u0_g62901 (.A1(u0_n_31951),
    .A2(u0_n_32338),
    .B(u0_n_31687),
    .C(n_11401),
    .Y(u0_n_30786));
 OAI211xp5_ASAP7_75t_R u0_g62902 (.A1(u0_n_31936),
    .A2(u0_n_31900),
    .B(u0_n_31689),
    .C(w3[0]),
    .Y(u0_n_30788));
 NOR2xp33_ASAP7_75t_R u0_g62903 (.A(u0_n_31093),
    .B(u0_n_31238),
    .Y(u0_n_30789));
 AOI21xp33_ASAP7_75t_R u0_g62904 (.A1(u0_n_31644),
    .A2(n_11457),
    .B(u0_n_31495),
    .Y(u0_n_30791));
 AO21x1_ASAP7_75t_R u0_g62905 (.A1(u0_n_31525),
    .A2(u0_n_31473),
    .B(u0_n_32121),
    .Y(u0_n_30793));
 A2O1A1Ixp33_ASAP7_75t_R u0_g62906 (.A1(u0_n_33001),
    .A2(u0_n_31808),
    .B(u0_n_32208),
    .C(u0_n_31489),
    .Y(u0_n_30796));
 AOI21xp33_ASAP7_75t_R u0_g62907 (.A1(u0_n_32339),
    .A2(u0_n_31487),
    .B(u0_n_31956),
    .Y(u0_n_30798));
 NOR2xp33_ASAP7_75t_R u0_g62908 (.A(u0_n_31477),
    .B(u0_n_31236),
    .Y(u0_n_30799));
 NAND2xp5_ASAP7_75t_L u0_g62909 (.A(w3[19]),
    .B(u0_n_31264),
    .Y(u0_n_30802));
 NAND2xp5_ASAP7_75t_L u0_g62910 (.A(\u0_w[3] [27]),
    .B(u0_n_31281),
    .Y(u0_n_30804));
 NOR2xp33_ASAP7_75t_L u0_g62911 (.A(n_11435),
    .B(u0_n_31285),
    .Y(u0_n_30806));
 NAND2xp33_ASAP7_75t_R u0_g62912 (.A(u0_n_31258),
    .B(u0_n_31138),
    .Y(u0_n_30808));
 AO21x1_ASAP7_75t_R u0_g62913 (.A1(u0_n_31874),
    .A2(u0_n_31461),
    .B(u0_n_31968),
    .Y(u0_n_30810));
 AND2x2_ASAP7_75t_L u0_g62914 (.A(u0_n_31646),
    .B(u0_n_31297),
    .Y(u0_n_30811));
 AO21x1_ASAP7_75t_R u0_g62915 (.A1(u0_n_32289),
    .A2(u0_n_31482),
    .B(u0_n_31974),
    .Y(u0_n_30814));
 OAI21xp33_ASAP7_75t_R u0_g62916 (.A1(u0_n_31518),
    .A2(u0_n_31449),
    .B(u0_n_32040),
    .Y(u0_n_30817));
 A2O1A1Ixp33_ASAP7_75t_L u0_g62917 (.A1(u0_n_32763),
    .A2(u0_n_31810),
    .B(u0_n_31895),
    .C(u0_n_31464),
    .Y(u0_n_30820));
 O2A1O1Ixp33_ASAP7_75t_R u0_g62918 (.A1(u0_n_32716),
    .A2(\u0_w[3] [27]),
    .B(u0_n_31536),
    .C(u0_n_31769),
    .Y(u0_n_30822));
 AND2x2_ASAP7_75t_L u0_g62919 (.A(u0_n_32040),
    .B(u0_n_31122),
    .Y(u0_n_30824));
 O2A1O1Ixp33_ASAP7_75t_SL u0_g62920 (.A1(w3[11]),
    .A2(u0_n_32714),
    .B(u0_n_31529),
    .C(u0_n_31762),
    .Y(u0_n_30825));
 AOI21xp33_ASAP7_75t_R u0_g62921 (.A1(u0_n_31543),
    .A2(u0_n_31916),
    .B(u0_n_31917),
    .Y(u0_n_30826));
 OAI31xp33_ASAP7_75t_R u0_g62922 (.A1(u0_n_32290),
    .A2(u0_n_31803),
    .A3(u0_n_32743),
    .B(u0_n_31751),
    .Y(u0_n_30828));
 OAI211xp5_ASAP7_75t_L u0_g62923 (.A1(w3[27]),
    .A2(n_8942),
    .B(u0_n_31088),
    .C(w3[30]),
    .Y(u0_n_30831));
 AOI21xp33_ASAP7_75t_R u0_g62924 (.A1(u0_n_31767),
    .A2(u0_n_31397),
    .B(u0_n_31755),
    .Y(u0_n_30833));
 OAI211xp5_ASAP7_75t_L u0_g62925 (.A1(u0_n_31935),
    .A2(u0_n_32242),
    .B(u0_n_31099),
    .C(u0_n_31393),
    .Y(u0_n_30835));
 OAI211xp5_ASAP7_75t_R u0_g62926 (.A1(u0_n_31920),
    .A2(u0_n_32141),
    .B(u0_n_31388),
    .C(u0_n_31108),
    .Y(u0_n_30837));
 OAI211xp5_ASAP7_75t_R u0_g62927 (.A1(u0_n_31922),
    .A2(u0_n_32387),
    .B(u0_n_31112),
    .C(u0_n_31396),
    .Y(u0_n_30840));
 OAI211xp5_ASAP7_75t_L u0_g62928 (.A1(w3[11]),
    .A2(\u0_w[3] [12]),
    .B(u0_n_31091),
    .C(n_8820),
    .Y(u0_n_30843));
 OAI31xp33_ASAP7_75t_L u0_g62929 (.A1(u0_n_31966),
    .A2(u0_n_31917),
    .A3(n_8831),
    .B(u0_n_31760),
    .Y(u0_n_30845));
 NOR2xp33_ASAP7_75t_R u0_g62930 (.A(u0_n_32385),
    .B(u0_n_31239),
    .Y(u0_n_30847));
 NAND2xp33_ASAP7_75t_R u0_g62931 (.A(u0_n_31986),
    .B(u0_n_31237),
    .Y(u0_n_30849));
 NAND2xp33_ASAP7_75t_R u0_g62932 (.A(u0_n_32122),
    .B(u0_n_31233),
    .Y(u0_n_30851));
 NOR2xp33_ASAP7_75t_L u0_g62933 (.A(u0_n_31534),
    .B(u0_n_31179),
    .Y(u0_n_30853));
 OR2x2_ASAP7_75t_SL u0_g62934 (.A(u0_n_31114),
    .B(u0_n_31249),
    .Y(u0_n_30854));
 NAND2xp33_ASAP7_75t_R u0_g62935 (.A(u0_n_32353),
    .B(u0_n_31142),
    .Y(u0_n_30857));
 NAND2xp33_ASAP7_75t_R u0_g62936 (.A(u0_n_32373),
    .B(u0_n_31141),
    .Y(u0_n_30858));
 NOR2xp33_ASAP7_75t_L u0_g62937 (.A(u0_n_31133),
    .B(u0_n_32290),
    .Y(u0_n_30859));
 AND2x2_ASAP7_75t_R u0_g62938 (.A(u0_n_31657),
    .B(u0_n_31261),
    .Y(u0_n_30861));
 NOR2xp33_ASAP7_75t_R u0_g62939 (.A(u0_n_31838),
    .B(u0_n_31291),
    .Y(u0_n_30864));
 NOR2xp33_ASAP7_75t_R u0_g62940 (.A(u0_n_31875),
    .B(u0_n_31136),
    .Y(u0_n_30867));
 NAND2xp33_ASAP7_75t_R u0_g62941 (.A(u0_n_32248),
    .B(u0_n_31329),
    .Y(u0_n_30868));
 AND2x2_ASAP7_75t_L u0_g62942 (.A(u0_n_31821),
    .B(u0_n_31308),
    .Y(u0_n_30869));
 NAND2xp33_ASAP7_75t_R u0_g62943 (.A(u0_n_32122),
    .B(u0_n_31286),
    .Y(u0_n_30871));
 OR2x2_ASAP7_75t_L u0_g62944 (.A(u0_n_32194),
    .B(u0_n_31162),
    .Y(u0_n_30872));
 NAND2xp5_ASAP7_75t_L u0_g62945 (.A(u0_n_31600),
    .B(u0_n_31158),
    .Y(u0_n_30873));
 NOR2xp33_ASAP7_75t_L u0_g62946 (.A(u0_n_32193),
    .B(u0_n_31324),
    .Y(u0_n_30875));
 NAND2xp33_ASAP7_75t_R u0_g62947 (.A(u0_n_32175),
    .B(u0_n_31166),
    .Y(u0_n_30876));
 NOR2xp33_ASAP7_75t_R u0_g62950 (.A(u0_n_32344),
    .B(u0_n_31120),
    .Y(u0_n_30717));
 NOR2xp33_ASAP7_75t_L u0_g62951 (.A(u0_n_32108),
    .B(u0_n_31116),
    .Y(u0_n_30718));
 NOR2xp33_ASAP7_75t_L u0_g62952 (.A(u0_n_31900),
    .B(u0_n_31161),
    .Y(u0_n_30720));
 NAND2xp5_ASAP7_75t_L u0_g62953 (.A(u0_n_32052),
    .B(u0_n_31117),
    .Y(u0_n_30721));
 NOR2xp33_ASAP7_75t_SL u0_g62954 (.A(u0_n_31900),
    .B(u0_n_31187),
    .Y(u0_n_30722));
 NAND2xp5_ASAP7_75t_L u0_g62955 (.A(u0_n_32208),
    .B(u0_n_31153),
    .Y(u0_n_30724));
 NAND2xp33_ASAP7_75t_R u0_g62956 (.A(n_11520),
    .B(u0_n_31332),
    .Y(u0_n_30725));
 NOR2xp33_ASAP7_75t_SL u0_g62957 (.A(u0_n_32290),
    .B(u0_n_31184),
    .Y(u0_n_30726));
 NOR2xp33_ASAP7_75t_R u0_g62958 (.A(u0_n_32083),
    .B(u0_n_31109),
    .Y(u0_n_30727));
 NOR2xp33_ASAP7_75t_L u0_g62959 (.A(u0_n_31524),
    .B(u0_n_31182),
    .Y(u0_n_30728));
 NAND2xp5_ASAP7_75t_L u0_g62960 (.A(u0_n_32273),
    .B(u0_n_31148),
    .Y(u0_n_30730));
 NOR2xp33_ASAP7_75t_R u0_g62961 (.A(n_11520),
    .B(u0_n_31332),
    .Y(u0_n_30731));
 NOR2xp33_ASAP7_75t_R u0_g62962 (.A(u0_n_31526),
    .B(u0_n_31186),
    .Y(u0_n_30732));
 NOR2xp33_ASAP7_75t_R u0_g62963 (.A(n_11520),
    .B(u0_n_31333),
    .Y(u0_n_30733));
 NOR2xp33_ASAP7_75t_R u0_g62964 (.A(u0_n_31664),
    .B(u0_n_31332),
    .Y(u0_n_30734));
 NAND2xp5_ASAP7_75t_R u0_g62965 (.A(u0_n_31184),
    .B(u0_n_31519),
    .Y(u0_n_30735));
 NAND2xp5_ASAP7_75t_L u0_g62966 (.A(u0_n_31181),
    .B(u0_n_31178),
    .Y(u0_n_30736));
 NAND2xp5_ASAP7_75t_L u0_g62967 (.A(u0_n_31319),
    .B(u0_n_32273),
    .Y(u0_n_30737));
 NAND2xp5_ASAP7_75t_L u0_g62968 (.A(u0_n_31183),
    .B(u0_n_31176),
    .Y(u0_n_30738));
 NOR2xp33_ASAP7_75t_R u0_g62969 (.A(u0_n_31522),
    .B(u0_n_31180),
    .Y(u0_n_30739));
 NOR2xp33_ASAP7_75t_SL u0_g62970 (.A(u0_n_32372),
    .B(u0_n_31111),
    .Y(u0_n_30740));
 NAND2xp33_ASAP7_75t_L u0_g62971 (.A(u0_n_31111),
    .B(u0_n_32304),
    .Y(u0_n_30741));
 NOR2xp67_ASAP7_75t_L u0_g62972 (.A(u0_n_32209),
    .B(u0_n_31317),
    .Y(u0_n_30743));
 NOR2xp33_ASAP7_75t_L u0_g62973 (.A(u0_n_32344),
    .B(u0_n_31313),
    .Y(u0_n_30744));
 NAND2xp5_ASAP7_75t_L u0_g62974 (.A(u0_n_32407),
    .B(u0_n_31101),
    .Y(u0_n_30745));
 NOR2xp33_ASAP7_75t_SL u0_g62975 (.A(u0_n_32194),
    .B(u0_n_31101),
    .Y(u0_n_30746));
 NOR2xp33_ASAP7_75t_R u0_g62976 (.A(u0_n_31846),
    .B(u0_n_31100),
    .Y(u0_n_30890));
 NAND2xp33_ASAP7_75t_R u0_g62977 (.A(u0_n_31100),
    .B(u0_n_32142),
    .Y(u0_n_30747));
 NAND2xp5_ASAP7_75t_L u0_g62978 (.A(u0_n_31837),
    .B(u0_n_31163),
    .Y(u0_n_30749));
 OR2x2_ASAP7_75t_L u0_g62979 (.A(u0_n_31817),
    .B(u0_n_31125),
    .Y(u0_n_30750));
 OR2x2_ASAP7_75t_L u0_g62980 (.A(u0_n_31822),
    .B(u0_n_31140),
    .Y(u0_n_30751));
 NAND2xp5_ASAP7_75t_R u0_g62981 (.A(u0_n_31687),
    .B(u0_n_31176),
    .Y(u0_n_30753));
 NOR2xp67_ASAP7_75t_R u0_g62982 (.A(n_8656),
    .B(u0_n_31282),
    .Y(u0_n_30754));
 NAND2xp5_ASAP7_75t_SL u0_g62983 (.A(u0_n_31273),
    .B(w3[27]),
    .Y(u0_n_30755));
 NOR2xp33_ASAP7_75t_L u0_g62984 (.A(u0_n_31776),
    .B(u0_n_31182),
    .Y(u0_n_30757));
 NOR2xp33_ASAP7_75t_L u0_g62985 (.A(u0_n_32749),
    .B(u0_n_31263),
    .Y(u0_n_30759));
 NOR2xp33_ASAP7_75t_R u0_g62986 (.A(u0_n_31772),
    .B(u0_n_31186),
    .Y(u0_n_30760));
 NAND2xp5_ASAP7_75t_SL u0_g62987 (.A(u0_n_31689),
    .B(u0_n_31174),
    .Y(u0_n_30761));
 NOR2xp33_ASAP7_75t_SL u0_g62988 (.A(u0_n_31316),
    .B(u0_n_31875),
    .Y(u0_n_30762));
 NOR2xp33_ASAP7_75t_R u0_g62989 (.A(u0_n_31786),
    .B(u0_n_31180),
    .Y(u0_n_30763));
 NAND2xp5_ASAP7_75t_R u0_g62990 (.A(u0_n_31184),
    .B(u0_n_31781),
    .Y(u0_n_30765));
 NOR2xp33_ASAP7_75t_SL u0_g62991 (.A(u0_n_31875),
    .B(u0_n_31174),
    .Y(u0_n_30767));
 NOR2xp33_ASAP7_75t_R u0_g62992 (.A(u0_n_31172),
    .B(u0_n_32272),
    .Y(u0_n_30768));
 NOR2xp33_ASAP7_75t_SL u0_g62993 (.A(u0_n_31680),
    .B(u0_n_31173),
    .Y(u0_n_30770));
 NAND2xp5_ASAP7_75t_L u0_g62994 (.A(u0_n_31178),
    .B(u0_n_31685),
    .Y(u0_n_30771));
 AOI21xp33_ASAP7_75t_R u0_g62995 (.A1(u0_n_31448),
    .A2(u0_r0_rcnt[3]),
    .B(u0_n_31110),
    .Y(u0_n_30773));
 NAND2xp5_ASAP7_75t_SL u0_g62996 (.A(w3[3]),
    .B(u0_n_31259),
    .Y(u0_n_30775));
 INVxp67_ASAP7_75t_SL u0_g62997 (.A(u0_n_30960),
    .Y(u0_n_30899));
 INVxp33_ASAP7_75t_R u0_g62998 (.A(u0_n_30977),
    .Y(u0_n_30900));
 INVxp67_ASAP7_75t_R u0_g62999 (.A(u0_n_30990),
    .Y(u0_n_30901));
 INVxp33_ASAP7_75t_R u0_g63000 (.A(u0_n_31033),
    .Y(u0_n_30902));
 INVxp33_ASAP7_75t_R u0_g63001 (.A(u0_n_30912),
    .Y(u0_n_30911));
 OAI221xp5_ASAP7_75t_SL u0_g63002 (.A1(u0_n_31631),
    .A2(u0_n_32749),
    .B1(u0_n_32344),
    .B2(\u0_w[3] [12]),
    .C(u0_n_31479),
    .Y(u0_n_30914));
 A2O1A1Ixp33_ASAP7_75t_R u0_g63003 (.A1(w3[14]),
    .A2(u0_n_31814),
    .B(u0_n_32339),
    .C(u0_n_31502),
    .Y(u0_n_30915));
 AOI211xp5_ASAP7_75t_SL u0_g63004 (.A1(u0_n_32289),
    .A2(u0_n_31930),
    .B(u0_n_31295),
    .C(u0_n_31406),
    .Y(u0_n_30918));
 AOI211xp5_ASAP7_75t_SL u0_g63005 (.A1(u0_n_32241),
    .A2(u0_n_31962),
    .B(u0_n_31086),
    .C(\u0_w[3] [16]),
    .Y(u0_n_30921));
 AO21x1_ASAP7_75t_R u0_g63006 (.A1(u0_n_31819),
    .A2(u0_n_31588),
    .B(u0_n_31086),
    .Y(u0_n_30922));
 AO21x1_ASAP7_75t_R u0_g63007 (.A1(u0_n_32260),
    .A2(u0_n_31465),
    .B(u0_n_31513),
    .Y(u0_n_30926));
 OR3x1_ASAP7_75t_R u0_g63008 (.A(u0_n_31417),
    .B(u0_n_31534),
    .C(u0_n_31918),
    .Y(u0_n_30928));
 AOI21xp33_ASAP7_75t_R u0_g63009 (.A1(u0_n_31840),
    .A2(u0_n_31977),
    .B(u0_n_31131),
    .Y(u0_n_30931));
 AO21x1_ASAP7_75t_L u0_g63010 (.A1(u0_n_32122),
    .A2(u0_n_31568),
    .B(u0_n_31817),
    .Y(u0_n_30932));
 OAI21xp33_ASAP7_75t_R u0_g63011 (.A1(u0_n_31522),
    .A2(u0_n_31493),
    .B(u0_n_31986),
    .Y(u0_n_30934));
 O2A1O1Ixp33_ASAP7_75t_L u0_g63012 (.A1(u0_n_31946),
    .A2(u0_n_31816),
    .B(u0_n_31895),
    .C(w3[2]),
    .Y(u0_n_30935));
 OAI21xp33_ASAP7_75t_R u0_g63013 (.A1(u0_n_32042),
    .A2(u0_n_31573),
    .B(u0_n_31830),
    .Y(u0_n_30936));
 OAI211xp5_ASAP7_75t_L u0_g63014 (.A1(u0_n_31938),
    .A2(u0_n_32410),
    .B(u0_n_31083),
    .C(u0_n_32745),
    .Y(u0_n_30938));
 OAI21xp33_ASAP7_75t_R u0_g63015 (.A1(u0_n_32011),
    .A2(u0_n_31601),
    .B(u0_n_31390),
    .Y(u0_n_30941));
 AOI211xp5_ASAP7_75t_L u0_g63016 (.A1(u0_n_32373),
    .A2(u0_n_31944),
    .B(u0_n_31087),
    .C(w3[24]),
    .Y(u0_n_30943));
 AOI22xp33_ASAP7_75t_R u0_g63017 (.A1(u0_n_31841),
    .A2(u0_n_31602),
    .B1(u0_n_31920),
    .B2(u0_n_32142),
    .Y(u0_n_30946));
 O2A1O1Ixp33_ASAP7_75t_R u0_g63018 (.A1(u0_n_32766),
    .A2(u0_n_31937),
    .B(u0_n_32075),
    .C(u0_n_31920),
    .Y(u0_n_30949));
 OAI22xp33_ASAP7_75t_R u0_g63019 (.A1(u0_n_31498),
    .A2(u0_n_32315),
    .B1(u0_n_31617),
    .B2(u0_n_32385),
    .Y(u0_n_30950));
 A2O1A1Ixp33_ASAP7_75t_R u0_g63020 (.A1(w3[30]),
    .A2(u0_n_31971),
    .B(u0_n_32052),
    .C(u0_n_31923),
    .Y(u0_n_30952));
 A2O1A1Ixp33_ASAP7_75t_R u0_g63021 (.A1(n_8820),
    .A2(u0_n_31951),
    .B(u0_n_32109),
    .C(u0_n_31929),
    .Y(u0_n_30953));
 OAI22xp33_ASAP7_75t_R u0_g63022 (.A1(u0_n_31464),
    .A2(u0_n_31846),
    .B1(u0_n_31615),
    .B2(u0_n_32165),
    .Y(u0_n_30956));
 AOI21xp33_ASAP7_75t_R u0_g63023 (.A1(u0_n_31679),
    .A2(u0_n_33004),
    .B(u0_n_32208),
    .Y(u0_n_30958));
 AOI221xp5_ASAP7_75t_L u0_g63024 (.A1(u0_n_32407),
    .A2(u0_n_31814),
    .B1(u0_n_32339),
    .B2(u0_n_32714),
    .C(u0_n_31647),
    .Y(u0_n_30959));
 A2O1A1Ixp33_ASAP7_75t_L u0_g63025 (.A1(u0_n_32793),
    .A2(u0_n_31959),
    .B(u0_n_32373),
    .C(u0_n_31269),
    .Y(u0_n_30960));
 OAI221xp5_ASAP7_75t_R u0_g63026 (.A1(u0_n_32254),
    .A2(u0_n_31807),
    .B1(u0_n_32221),
    .B2(n_8831),
    .C(u0_n_31657),
    .Y(u0_n_30961));
 O2A1O1Ixp33_ASAP7_75t_R u0_g63027 (.A1(u0_n_33001),
    .A2(u0_n_31966),
    .B(u0_n_32254),
    .C(u0_n_31271),
    .Y(u0_n_30963));
 AOI221xp5_ASAP7_75t_R u0_g63028 (.A1(u0_n_32166),
    .A2(u0_n_31810),
    .B1(u0_n_31874),
    .B2(u0_n_32697),
    .C(u0_n_31639),
    .Y(u0_n_30964));
 NAND3xp33_ASAP7_75t_L u0_g63029 (.A(u0_n_31244),
    .B(u0_n_31657),
    .C(u0_n_31404),
    .Y(u0_n_30967));
 O2A1O1Ixp33_ASAP7_75t_R u0_g63030 (.A1(u0_n_32763),
    .A2(u0_n_31964),
    .B(u0_n_32165),
    .C(u0_n_31124),
    .Y(u0_n_30969));
 OAI21xp33_ASAP7_75t_R u0_g63031 (.A1(u0_n_31792),
    .A2(u0_n_31537),
    .B(u0_n_32373),
    .Y(u0_n_30971));
 AOI21xp5_ASAP7_75t_R u0_g63032 (.A1(u0_n_31793),
    .A2(u0_n_31529),
    .B(u0_n_32410),
    .Y(u0_n_30972));
 AOI21xp33_ASAP7_75t_R u0_g63033 (.A1(u0_n_31531),
    .A2(u0_n_31795),
    .B(u0_n_32141),
    .Y(u0_n_30975));
 AO21x1_ASAP7_75t_R u0_g63034 (.A1(u0_n_31970),
    .A2(u0_n_31665),
    .B(u0_n_32344),
    .Y(u0_n_30976));
 A2O1A1Ixp33_ASAP7_75t_R u0_g63035 (.A1(u0_n_31976),
    .A2(u0_n_31823),
    .B(u0_n_32053),
    .C(u0_n_31621),
    .Y(u0_n_30977));
 OAI21xp33_ASAP7_75t_R u0_g63036 (.A1(u0_n_31792),
    .A2(u0_n_31682),
    .B(u0_n_32308),
    .Y(u0_n_30978));
 OAI21xp33_ASAP7_75t_R u0_g63037 (.A1(u0_n_31462),
    .A2(u0_n_31493),
    .B(u0_n_32241),
    .Y(u0_n_30980));
 NAND4xp25_ASAP7_75t_R u0_g63038 (.A(u0_n_31494),
    .B(u0_n_31463),
    .C(u0_n_31754),
    .D(u0_n_33001),
    .Y(u0_n_30983));
 OAI21xp33_ASAP7_75t_R u0_g63039 (.A1(u0_n_31796),
    .A2(u0_n_31533),
    .B(u0_n_31850),
    .Y(u0_n_30985));
 OAI21xp33_ASAP7_75t_R u0_g63040 (.A1(u0_n_31794),
    .A2(u0_n_31539),
    .B(u0_n_32193),
    .Y(u0_n_30986));
 OAI21xp33_ASAP7_75t_R u0_g63041 (.A1(u0_n_31800),
    .A2(u0_n_31534),
    .B(u0_n_32012),
    .Y(u0_n_30987));
 OAI211xp5_ASAP7_75t_L u0_g63042 (.A1(u0_n_32717),
    .A2(u0_n_32290),
    .B(u0_n_31643),
    .C(u0_n_31360),
    .Y(u0_n_30988));
 OAI22xp5_ASAP7_75t_L u0_g63043 (.A1(u0_n_32174),
    .A2(u0_n_31502),
    .B1(u0_n_31604),
    .B2(u0_n_32409),
    .Y(u0_n_30990));
 NAND3xp33_ASAP7_75t_R u0_g63044 (.A(u0_n_31279),
    .B(u0_n_31643),
    .C(u0_n_31427),
    .Y(u0_n_30992));
 OAI21xp5_ASAP7_75t_R u0_g63045 (.A1(n_8820),
    .A2(u0_n_31392),
    .B(u0_n_31246),
    .Y(u0_n_30994));
 A2O1A1Ixp33_ASAP7_75t_R u0_g63046 (.A1(u0_n_31821),
    .A2(u0_n_31799),
    .B(u0_n_32221),
    .C(u0_n_32254),
    .Y(u0_n_30996));
 OAI21xp33_ASAP7_75t_R u0_g63047 (.A1(u0_n_31674),
    .A2(u0_n_31686),
    .B(u0_n_32407),
    .Y(u0_n_30997));
 OA211x2_ASAP7_75t_R u0_g63048 (.A1(u0_n_31801),
    .A2(u0_n_31425),
    .B(u0_n_31777),
    .C(u0_n_32685),
    .Y(u0_n_30998));
 AOI22xp33_ASAP7_75t_R u0_g63049 (.A1(u0_n_32749),
    .A2(u0_n_31488),
    .B1(u0_n_31969),
    .B2(u0_n_32407),
    .Y(u0_n_31000));
 AO22x1_ASAP7_75t_L u0_g63050 (.A1(u0_n_31998),
    .A2(u0_n_31638),
    .B1(u0_n_31935),
    .B2(u0_n_32260),
    .Y(u0_n_31001));
 OAI211xp5_ASAP7_75t_R u0_g63051 (.A1(u0_n_31811),
    .A2(u0_n_31404),
    .B(u0_n_31759),
    .C(u0_n_31770),
    .Y(u0_n_31002));
 AOI221xp5_ASAP7_75t_R u0_g63052 (.A1(u0_n_31753),
    .A2(u0_n_31820),
    .B1(u0_n_31465),
    .B2(w3[19]),
    .C(u0_n_33001),
    .Y(u0_n_31004));
 OAI211xp5_ASAP7_75t_R u0_g63053 (.A1(u0_n_31954),
    .A2(u0_n_32221),
    .B(u0_n_31685),
    .C(\u0_w[3] [16]),
    .Y(u0_n_31005));
 AO22x1_ASAP7_75t_L u0_g63054 (.A1(u0_n_31465),
    .A2(u0_n_31469),
    .B1(u0_n_31679),
    .B2(u0_n_31435),
    .Y(u0_n_31006));
 OAI221xp5_ASAP7_75t_L u0_g63055 (.A1(u0_n_32372),
    .A2(u0_n_31971),
    .B1(u0_n_31972),
    .B2(\u0_w[3] [27]),
    .C(u0_n_31342),
    .Y(u0_n_31009));
 AOI22xp33_ASAP7_75t_R u0_g63056 (.A1(u0_n_32208),
    .A2(u0_n_31608),
    .B1(u0_n_32241),
    .B2(u0_n_31480),
    .Y(u0_n_31011));
 AOI22xp33_ASAP7_75t_R u0_g63057 (.A1(u0_n_32273),
    .A2(u0_n_31431),
    .B1(u0_n_31960),
    .B2(u0_n_32304),
    .Y(u0_n_31012));
 AOI22xp33_ASAP7_75t_L u0_g63058 (.A1(u0_n_32353),
    .A2(u0_n_31605),
    .B1(u0_n_32407),
    .B2(u0_n_31418),
    .Y(u0_n_31014));
 AOI22xp33_ASAP7_75t_L u0_g63059 (.A1(u0_n_31874),
    .A2(u0_n_31616),
    .B1(u0_n_32142),
    .B2(u0_n_31424),
    .Y(u0_n_31016));
 AOI221xp5_ASAP7_75t_R u0_g63060 (.A1(u0_n_31627),
    .A2(u0_n_32021),
    .B1(u0_n_32241),
    .B2(u0_n_31953),
    .C(u0_n_31552),
    .Y(u0_n_31017));
 OAI221xp5_ASAP7_75t_R u0_g63061 (.A1(u0_n_32053),
    .A2(n_8942),
    .B1(u0_n_31805),
    .B2(u0_n_32793),
    .C(w3[26]),
    .Y(u0_n_31019));
 OAI222xp33_ASAP7_75t_R u0_g63062 (.A1(u0_n_32410),
    .A2(u0_n_31951),
    .B1(u0_n_31623),
    .B2(u0_n_32185),
    .C1(u0_n_31952),
    .C2(w3[11]),
    .Y(u0_n_31021));
 OAI22xp33_ASAP7_75t_R u0_g63063 (.A1(u0_n_31424),
    .A2(u0_n_31900),
    .B1(u0_n_31963),
    .B2(u0_n_31842),
    .Y(u0_n_31023));
 AOI22xp33_ASAP7_75t_R u0_g63064 (.A1(u0_n_32241),
    .A2(u0_n_31493),
    .B1(n_8831),
    .B2(u0_n_32012),
    .Y(u0_n_31026));
 AOI22xp33_ASAP7_75t_R u0_g63065 (.A1(u0_n_31481),
    .A2(u0_n_32226),
    .B1(u0_n_32012),
    .B2(u0_n_31966),
    .Y(u0_n_31027));
 AOI22xp5_ASAP7_75t_L u0_g63066 (.A1(u0_n_32040),
    .A2(u0_n_31483),
    .B1(u0_n_31922),
    .B2(u0_n_32373),
    .Y(u0_n_31028));
 OAI221xp5_ASAP7_75t_SL u0_g63067 (.A1(u0_n_32165),
    .A2(u0_n_31936),
    .B1(u0_n_31937),
    .B2(w3[3]),
    .C(u0_n_31340),
    .Y(u0_n_31030));
 OAI22xp33_ASAP7_75t_R u0_g63068 (.A1(u0_n_32344),
    .A2(u0_n_31610),
    .B1(u0_n_32108),
    .B2(u0_n_31487),
    .Y(u0_n_31033));
 AO22x1_ASAP7_75t_R u0_g63069 (.A1(u0_n_32304),
    .A2(u0_n_31576),
    .B1(u0_n_31803),
    .B2(u0_n_32289),
    .Y(u0_n_31036));
 AOI221xp5_ASAP7_75t_R u0_g63070 (.A1(u0_n_32339),
    .A2(u0_n_31926),
    .B1(u0_n_31471),
    .B2(u0_n_32407),
    .C(u0_n_31411),
    .Y(u0_n_31038));
 AOI211xp5_ASAP7_75t_R u0_g63071 (.A1(u0_n_31428),
    .A2(u0_n_31805),
    .B(u0_n_31768),
    .C(w3[26]),
    .Y(u0_n_31040));
 AO22x1_ASAP7_75t_R u0_g63072 (.A1(u0_n_31823),
    .A2(u0_n_31584),
    .B1(u0_n_32320),
    .B2(u0_n_31606),
    .Y(u0_n_31041));
 AOI22xp33_ASAP7_75t_R u0_g63073 (.A1(u0_n_31587),
    .A2(u0_n_31840),
    .B1(u0_n_31613),
    .B2(u0_n_31850),
    .Y(u0_n_31043));
 AOI22xp33_ASAP7_75t_R u0_g63074 (.A1(u0_n_31826),
    .A2(u0_n_31591),
    .B1(u0_n_32184),
    .B2(u0_n_31611),
    .Y(u0_n_31045));
 AOI22xp33_ASAP7_75t_R u0_g63075 (.A1(u0_n_32273),
    .A2(u0_n_31629),
    .B1(u0_n_31976),
    .B2(u0_n_31401),
    .Y(u0_n_31048));
 AOI22xp33_ASAP7_75t_R u0_g63076 (.A1(w3[3]),
    .A2(u0_n_31586),
    .B1(u0_n_32737),
    .B2(u0_n_31531),
    .Y(u0_n_31050));
 AOI22xp33_ASAP7_75t_R u0_g63077 (.A1(u0_n_31594),
    .A2(u0_n_31678),
    .B1(u0_n_31820),
    .B2(u0_n_31998),
    .Y(u0_n_31051));
 AOI32xp33_ASAP7_75t_R u0_g63078 (.A1(u0_n_32142),
    .A2(u0_n_31977),
    .A3(n_8747),
    .B1(u0_n_32084),
    .B2(u0_n_31936),
    .Y(u0_n_31053));
 AOI22xp33_ASAP7_75t_R u0_g63079 (.A1(w3[27]),
    .A2(u0_n_31580),
    .B1(u0_n_32751),
    .B2(u0_n_31536),
    .Y(u0_n_31054));
 AOI32xp33_ASAP7_75t_R u0_g63080 (.A1(u0_n_32407),
    .A2(u0_n_31983),
    .A3(n_8851),
    .B1(u0_n_32109),
    .B2(u0_n_31951),
    .Y(u0_n_31055));
 OAI22xp33_ASAP7_75t_R u0_g63081 (.A1(u0_n_32773),
    .A2(u0_n_31626),
    .B1(u0_n_31964),
    .B2(u0_n_31875),
    .Y(u0_n_31056));
 OAI221xp5_ASAP7_75t_L u0_g63082 (.A1(u0_n_31669),
    .A2(n_8820),
    .B1(u0_n_32410),
    .B2(u0_n_32759),
    .C(u0_n_31955),
    .Y(u0_n_31057));
 AOI22xp33_ASAP7_75t_R u0_g63083 (.A1(u0_n_31590),
    .A2(w3[19]),
    .B1(u0_n_31543),
    .B2(n_8656),
    .Y(u0_n_31059));
 OAI22xp33_ASAP7_75t_R u0_g63084 (.A1(n_8801),
    .A2(u0_n_31582),
    .B1(u0_n_31982),
    .B2(u0_n_32338),
    .Y(u0_n_31061));
 AOI22xp33_ASAP7_75t_R u0_g63085 (.A1(u0_n_33033),
    .A2(u0_n_31579),
    .B1(u0_n_31976),
    .B2(u0_n_32273),
    .Y(u0_n_31063));
 OAI22xp33_ASAP7_75t_R u0_g63086 (.A1(u0_n_31875),
    .A2(u0_n_31672),
    .B1(u0_n_31773),
    .B2(u0_n_32141),
    .Y(u0_n_31064));
 OAI22xp33_ASAP7_75t_R u0_g63087 (.A1(u0_n_32344),
    .A2(u0_n_31668),
    .B1(u0_n_31775),
    .B2(u0_n_32410),
    .Y(u0_n_31065));
 OAI221xp5_ASAP7_75t_R u0_g63088 (.A1(u0_n_32763),
    .A2(u0_n_31673),
    .B1(u0_n_32160),
    .B2(n_8625),
    .C(u0_n_31967),
    .Y(u0_n_31066));
 AOI22xp33_ASAP7_75t_R u0_g63089 (.A1(u0_n_31589),
    .A2(u0_n_33001),
    .B1(u0_n_31985),
    .B2(u0_n_32208),
    .Y(u0_n_31068));
 OAI221xp5_ASAP7_75t_R u0_g63090 (.A1(u0_n_31666),
    .A2(u0_n_33001),
    .B1(u0_n_32254),
    .B2(u0_n_33138),
    .C(u0_n_31957),
    .Y(u0_n_31069));
 AOI22xp33_ASAP7_75t_R u0_g63091 (.A1(u0_n_32175),
    .A2(u0_n_31575),
    .B1(u0_n_32353),
    .B2(u0_n_31813),
    .Y(u0_n_31070));
 OAI22xp33_ASAP7_75t_R u0_g63092 (.A1(u0_n_32209),
    .A2(u0_n_31667),
    .B1(u0_n_32254),
    .B2(u0_n_31785),
    .Y(u0_n_31072));
 AOI221xp5_ASAP7_75t_R u0_g63093 (.A1(u0_n_31659),
    .A2(u0_n_32793),
    .B1(u0_n_32386),
    .B2(n_8942),
    .C(u0_n_31974),
    .Y(u0_n_31073));
 AOI22xp33_ASAP7_75t_R u0_g63094 (.A1(u0_n_31486),
    .A2(\u0_w[3] [27]),
    .B1(u0_n_32751),
    .B2(u0_n_31518),
    .Y(u0_n_30903));
 XNOR2xp5_ASAP7_75t_R u0_g63095 (.A(u0_n_31714),
    .B(u0_n_32675),
    .Y(u0_n_30904));
 AOI22xp33_ASAP7_75t_R u0_g63096 (.A1(n_11457),
    .A2(u0_n_31466),
    .B1(u0_n_32737),
    .B2(u0_n_31526),
    .Y(u0_n_30905));
 XNOR2xp5_ASAP7_75t_R u0_g63097 (.A(u0_n_31733),
    .B(w1[30]),
    .Y(u0_n_31076));
 XOR2xp5_ASAP7_75t_R u0_g63098 (.A(u0_n_31712),
    .B(w1[10]),
    .Y(u0_n_30906));
 OAI22xp33_ASAP7_75t_R u0_g63099 (.A1(n_11435),
    .A2(u0_n_31524),
    .B1(u0_n_32749),
    .B2(u0_n_31471),
    .Y(u0_n_30907));
 AO21x1_ASAP7_75t_R u0_g63100 (.A1(u0_n_31812),
    .A2(u0_n_31678),
    .B(u0_n_31988),
    .Y(u0_n_30908));
 AND3x1_ASAP7_75t_R u0_g63101 (.A(u0_n_31170),
    .B(u0_n_32386),
    .C(u0_n_31830),
    .Y(u0_n_30909));
 AOI22xp33_ASAP7_75t_L u0_g63102 (.A1(u0_n_31446),
    .A2(w3[19]),
    .B1(u0_n_31522),
    .B2(n_8656),
    .Y(u0_n_30910));
 NOR3xp33_ASAP7_75t_SL u0_g63103 (.A(u0_n_31542),
    .B(u0_n_31450),
    .C(u0_n_32254),
    .Y(u0_n_30912));
 AO21x1_ASAP7_75t_L u0_g63104 (.A1(u0_n_32021),
    .A2(u0_n_31542),
    .B(u0_n_31089),
    .Y(u0_n_30913));
 INVxp33_ASAP7_75t_R u0_g63105 (.A(u0_n_31085),
    .Y(u0_n_31084));
 INVxp33_ASAP7_75t_R u0_g63106 (.A(u0_n_31094),
    .Y(u0_n_31093));
 INVxp67_ASAP7_75t_R u0_g63107 (.A(u0_n_31104),
    .Y(u0_n_31103));
 INVxp67_ASAP7_75t_R u0_g63108 (.A(u0_n_31107),
    .Y(u0_n_31106));
 INVxp67_ASAP7_75t_R u0_g63109 (.A(u0_n_31124),
    .Y(u0_n_31123));
 INVxp67_ASAP7_75t_L u0_g63110 (.A(u0_n_31126),
    .Y(u0_n_31127));
 INVx1_ASAP7_75t_L u0_g63111 (.A(u0_n_31129),
    .Y(u0_n_31128));
 INVxp67_ASAP7_75t_R u0_g63112 (.A(u0_n_31134),
    .Y(u0_n_31133));
 INVxp67_ASAP7_75t_R u0_g63113 (.A(u0_n_31146),
    .Y(u0_n_31145));
 INVx1_ASAP7_75t_L u0_g63114 (.A(u0_n_31150),
    .Y(u0_n_31149));
 INVxp33_ASAP7_75t_R u0_g63115 (.A(u0_n_31153),
    .Y(u0_n_31152));
 INVxp67_ASAP7_75t_R u0_g63116 (.A(u0_n_31155),
    .Y(u0_n_31154));
 INVxp33_ASAP7_75t_L u0_g63117 (.A(u0_n_31158),
    .Y(u0_n_31157));
 INVxp67_ASAP7_75t_R u0_g63118 (.A(u0_n_31160),
    .Y(u0_n_31159));
 INVxp67_ASAP7_75t_R u0_g63119 (.A(u0_n_31165),
    .Y(u0_n_31164));
 INVxp67_ASAP7_75t_R u0_g63120 (.A(u0_n_31169),
    .Y(u0_n_31168));
 INVx1_ASAP7_75t_SL u0_g63121 (.A(u0_n_31172),
    .Y(u0_n_31173));
 INVxp33_ASAP7_75t_R u0_g63122 (.A(u0_n_31174),
    .Y(u0_n_31175));
 INVx1_ASAP7_75t_R u0_g63123 (.A(u0_n_31176),
    .Y(u0_n_31177));
 INVxp67_ASAP7_75t_R u0_g63124 (.A(u0_n_31178),
    .Y(u0_n_31179));
 INVx1_ASAP7_75t_SL u0_g63125 (.A(u0_n_31180),
    .Y(u0_n_31181));
 INVxp67_ASAP7_75t_R u0_g63126 (.A(u0_n_31182),
    .Y(u0_n_31183));
 INVxp33_ASAP7_75t_R u0_g63127 (.A(u0_n_31184),
    .Y(u0_n_31185));
 INVx1_ASAP7_75t_L u0_g63128 (.A(u0_n_31186),
    .Y(u0_n_31187));
 AND2x2_ASAP7_75t_R u0_g63129 (.A(u0_n_32877),
    .B(u0_n_31448),
    .Y(u0_n_31188));
 NAND2xp33_ASAP7_75t_R u0_g63130 (.A(u0_n_31959),
    .B(u0_n_31655),
    .Y(u0_n_31190));
 NAND2xp33_ASAP7_75t_R u0_g63131 (.A(n_11516),
    .B(u0_n_31963),
    .Y(u0_n_31191));
 NAND2xp33_ASAP7_75t_R u0_g63132 (.A(u0_n_31929),
    .B(u0_n_31444),
    .Y(u0_n_31192));
 NOR2xp33_ASAP7_75t_R u0_g63133 (.A(n_11435),
    .B(u0_n_31528),
    .Y(u0_n_31193));
 NOR2xp33_ASAP7_75t_R u0_g63134 (.A(u0_n_31499),
    .B(u0_n_31644),
    .Y(u0_n_31195));
 NOR2xp33_ASAP7_75t_R u0_g63135 (.A(u0_n_31450),
    .B(u0_n_31632),
    .Y(u0_n_31196));
 NAND2xp33_ASAP7_75t_R u0_g63136 (.A(u0_n_31577),
    .B(u0_n_31427),
    .Y(u0_n_31198));
 NAND2xp33_ASAP7_75t_R u0_g63137 (.A(u0_n_32835),
    .B(u0_n_31664),
    .Y(u0_n_31200));
 NOR2xp33_ASAP7_75t_R u0_g63138 (.A(u0_n_31526),
    .B(u0_n_31499),
    .Y(u0_n_31202));
 NAND2xp33_ASAP7_75t_R u0_g63139 (.A(u0_n_31400),
    .B(u0_n_31821),
    .Y(u0_n_31081));
 NAND2xp33_ASAP7_75t_R u0_g63140 (.A(u0_n_32080),
    .B(u0_n_31397),
    .Y(u0_n_31082));
 NAND2xp5_ASAP7_75t_L u0_g63141 (.A(u0_n_32113),
    .B(u0_n_31395),
    .Y(u0_n_31083));
 NAND2xp5_ASAP7_75t_R u0_g63142 (.A(u0_n_32353),
    .B(u0_n_31473),
    .Y(u0_n_31085));
 AND2x2_ASAP7_75t_L u0_g63143 (.A(u0_n_31965),
    .B(u0_n_31402),
    .Y(u0_n_31086));
 NOR2xp33_ASAP7_75t_L u0_g63144 (.A(u0_n_31399),
    .B(u0_n_32042),
    .Y(u0_n_31087));
 NOR2xp33_ASAP7_75t_SL u0_g63145 (.A(u0_n_31430),
    .B(u0_n_31449),
    .Y(u0_n_31088));
 AND2x2_ASAP7_75t_SL u0_g63146 (.A(u0_n_32012),
    .B(u0_n_31450),
    .Y(u0_n_31089));
 NAND2xp33_ASAP7_75t_R u0_g63147 (.A(u0_n_32040),
    .B(u0_n_31485),
    .Y(u0_n_31090));
 AND2x2_ASAP7_75t_L u0_g63148 (.A(u0_n_31473),
    .B(u0_n_31631),
    .Y(u0_n_31091));
 NAND2xp33_ASAP7_75t_R u0_g63149 (.A(u0_n_31986),
    .B(u0_n_31445),
    .Y(u0_n_31092));
 NAND2xp33_ASAP7_75t_R u0_g63150 (.A(u0_n_32175),
    .B(u0_n_31418),
    .Y(u0_n_31094));
 NAND2xp33_ASAP7_75t_R u0_g63151 (.A(u0_n_31546),
    .B(n_8629),
    .Y(u0_n_31095));
 NAND2xp33_ASAP7_75t_L u0_g63152 (.A(u0_n_32080),
    .B(u0_n_31467),
    .Y(u0_n_31096));
 NOR2xp33_ASAP7_75t_R u0_g63153 (.A(u0_n_32759),
    .B(u0_n_31540),
    .Y(u0_n_31097));
 NAND2xp33_ASAP7_75t_R u0_g63154 (.A(w3[20]),
    .B(u0_n_31544),
    .Y(u0_n_31098));
 NAND2xp33_ASAP7_75t_R u0_g63155 (.A(u0_n_32012),
    .B(u0_n_31480),
    .Y(u0_n_31099));
 NOR2xp33_ASAP7_75t_SL u0_g63156 (.A(u0_n_31530),
    .B(u0_n_31484),
    .Y(u0_n_31100));
 NOR2xp33_ASAP7_75t_L u0_g63157 (.A(u0_n_31528),
    .B(u0_n_31470),
    .Y(u0_n_31101));
 NAND2xp33_ASAP7_75t_R u0_g63158 (.A(u0_n_31548),
    .B(w3[28]),
    .Y(u0_n_31102));
 NOR2xp33_ASAP7_75t_R u0_g63159 (.A(u0_n_31534),
    .B(u0_n_31450),
    .Y(u0_n_31104));
 NOR2xp33_ASAP7_75t_L u0_g63160 (.A(u0_n_31533),
    .B(u0_n_31484),
    .Y(u0_n_31105));
 NOR2xp33_ASAP7_75t_R u0_g63161 (.A(u0_n_31470),
    .B(u0_n_31539),
    .Y(u0_n_31107));
 NAND2xp5_ASAP7_75t_R u0_g63162 (.A(u0_n_31850),
    .B(u0_n_31424),
    .Y(u0_n_31108));
 NOR2xp33_ASAP7_75t_R u0_g63163 (.A(u0_n_31816),
    .B(u0_n_31676),
    .Y(u0_n_31109));
 NOR2xp33_ASAP7_75t_R u0_g63164 (.A(u0_r0_rcnt[3]),
    .B(u0_n_31448),
    .Y(u0_n_31110));
 NAND2xp5_ASAP7_75t_L u0_g63165 (.A(u0_n_31536),
    .B(u0_n_31651),
    .Y(u0_n_31111));
 OR2x2_ASAP7_75t_R u0_g63166 (.A(u0_n_32315),
    .B(u0_n_31431),
    .Y(u0_n_31112));
 NAND2xp33_ASAP7_75t_R u0_g63167 (.A(u0_n_31651),
    .B(u0_n_31683),
    .Y(u0_n_31113));
 NOR2xp33_ASAP7_75t_L u0_g63168 (.A(u0_n_31499),
    .B(u0_n_31875),
    .Y(u0_n_31114));
 NOR2xp33_ASAP7_75t_SL u0_g63169 (.A(u0_n_32209),
    .B(u0_n_31493),
    .Y(u0_n_31115));
 NOR2xp33_ASAP7_75t_L u0_g63170 (.A(u0_n_31801),
    .B(u0_n_31674),
    .Y(u0_n_31116));
 NAND2xp5_ASAP7_75t_L u0_g63171 (.A(u0_n_31671),
    .B(u0_n_31805),
    .Y(u0_n_31117));
 OR2x2_ASAP7_75t_R u0_g63172 (.A(u0_n_32108),
    .B(u0_n_31471),
    .Y(u0_n_31118));
 NOR2xp33_ASAP7_75t_R u0_g63173 (.A(u0_n_32290),
    .B(u0_n_31449),
    .Y(u0_n_31119));
 NOR2x1_ASAP7_75t_L u0_g63174 (.A(u0_n_31814),
    .B(u0_n_31686),
    .Y(u0_n_31120));
 NOR2xp33_ASAP7_75t_R u0_g63175 (.A(u0_n_31846),
    .B(u0_n_31495),
    .Y(u0_n_31121));
 NOR2xp33_ASAP7_75t_L u0_g63176 (.A(u0_n_31416),
    .B(u0_n_31485),
    .Y(u0_n_31122));
 NAND2xp5_ASAP7_75t_L u0_g63177 (.A(u0_n_31457),
    .B(u0_n_31689),
    .Y(u0_n_31124));
 NOR2xp67_ASAP7_75t_SL u0_g63178 (.A(\u0_w[3] [12]),
    .B(u0_n_31541),
    .Y(u0_n_31125));
 NOR2xp33_ASAP7_75t_SL u0_g63179 (.A(u0_n_31838),
    .B(u0_n_31456),
    .Y(u0_n_31126));
 NOR2xp33_ASAP7_75t_L u0_g63180 (.A(u0_n_32017),
    .B(u0_n_31510),
    .Y(u0_n_31129));
 NOR2xp33_ASAP7_75t_R u0_g63181 (.A(u0_n_31820),
    .B(u0_n_31522),
    .Y(u0_n_31130));
 NAND2xp5_ASAP7_75t_L u0_g63182 (.A(u0_n_32080),
    .B(u0_n_31496),
    .Y(u0_n_31131));
 NOR2xp33_ASAP7_75t_L u0_g63183 (.A(u0_n_31456),
    .B(u0_n_31467),
    .Y(u0_n_31132));
 NAND2xp5_ASAP7_75t_L u0_g63184 (.A(u0_n_31823),
    .B(u0_n_31519),
    .Y(u0_n_31134));
 NOR2xp33_ASAP7_75t_L u0_g63185 (.A(u0_n_31492),
    .B(u0_n_31682),
    .Y(u0_n_31135));
 NOR2xp33_ASAP7_75t_R u0_g63186 (.A(u0_n_31839),
    .B(u0_n_31526),
    .Y(u0_n_31136));
 NAND2xp5_ASAP7_75t_L u0_g63187 (.A(u0_n_31415),
    .B(u0_n_31805),
    .Y(u0_n_31137));
 NOR2xp33_ASAP7_75t_R u0_g63188 (.A(u0_n_31875),
    .B(u0_n_31495),
    .Y(u0_n_31138));
 NAND2xp5_ASAP7_75t_L u0_g63189 (.A(u0_n_32142),
    .B(u0_n_31496),
    .Y(u0_n_31139));
 NOR2xp33_ASAP7_75t_SL u0_g63190 (.A(w3[20]),
    .B(u0_n_31544),
    .Y(u0_n_31140));
 NAND2xp5_ASAP7_75t_R u0_g63191 (.A(u0_n_31803),
    .B(u0_n_31536),
    .Y(u0_n_31141));
 NAND2xp5_ASAP7_75t_R u0_g63192 (.A(u0_n_31826),
    .B(u0_n_31525),
    .Y(u0_n_31142));
 NOR2xp33_ASAP7_75t_L u0_g63193 (.A(u0_n_31534),
    .B(u0_n_31501),
    .Y(u0_n_31143));
 NOR2xp33_ASAP7_75t_R u0_g63194 (.A(u0_n_31503),
    .B(u0_n_31533),
    .Y(u0_n_31144));
 NAND2xp5_ASAP7_75t_L u0_g63195 (.A(u0_n_31809),
    .B(u0_n_31531),
    .Y(u0_n_31146));
 NAND2xp5_ASAP7_75t_L u0_g63196 (.A(u0_n_31986),
    .B(u0_n_31509),
    .Y(u0_n_31147));
 NAND2xp5_ASAP7_75t_SL u0_g63197 (.A(u0_n_31681),
    .B(u0_n_31803),
    .Y(u0_n_31148));
 NAND2xp5_ASAP7_75t_L u0_g63198 (.A(u0_n_31807),
    .B(u0_n_31543),
    .Y(u0_n_31150));
 NAND2xp33_ASAP7_75t_R u0_g63199 (.A(u0_n_31538),
    .B(u0_n_31508),
    .Y(u0_n_31151));
 NAND2xp5_ASAP7_75t_L u0_g63200 (.A(u0_n_31807),
    .B(u0_n_31685),
    .Y(u0_n_31153));
 NAND2xp5_ASAP7_75t_R u0_g63201 (.A(u0_n_31457),
    .B(u0_n_31815),
    .Y(u0_n_31155));
 NOR2xp33_ASAP7_75t_R u0_g63202 (.A(u0_n_31801),
    .B(u0_n_31437),
    .Y(u0_n_31156));
 NOR2xp33_ASAP7_75t_L u0_g63203 (.A(u0_n_32254),
    .B(u0_n_31510),
    .Y(u0_n_31158));
 NOR2xp33_ASAP7_75t_SL u0_g63204 (.A(u0_n_32221),
    .B(u0_n_31510),
    .Y(u0_n_31160));
 NOR2xp33_ASAP7_75t_L u0_g63205 (.A(u0_n_31810),
    .B(u0_n_31688),
    .Y(u0_n_31161));
 NOR2xp33_ASAP7_75t_L u0_g63206 (.A(u0_n_31814),
    .B(u0_n_31528),
    .Y(u0_n_31162));
 NAND2xp5_ASAP7_75t_L u0_g63207 (.A(n_8625),
    .B(u0_n_31547),
    .Y(u0_n_31163));
 NOR2xp33_ASAP7_75t_L u0_g63208 (.A(u0_n_31811),
    .B(u0_n_31421),
    .Y(u0_n_31165));
 NOR2xp33_ASAP7_75t_SL u0_g63209 (.A(u0_n_31686),
    .B(u0_n_31437),
    .Y(u0_n_31166));
 NAND2xp5_ASAP7_75t_R u0_g63210 (.A(u0_n_31400),
    .B(u0_n_31481),
    .Y(u0_n_31167));
 NAND2xp33_ASAP7_75t_R u0_g63211 (.A(u0_n_31436),
    .B(u0_n_31471),
    .Y(u0_n_31169));
 NAND2xp5_ASAP7_75t_R u0_g63212 (.A(n_8964),
    .B(u0_n_31549),
    .Y(u0_n_31170));
 NAND2xp5_ASAP7_75t_SL u0_g63213 (.A(n_8946),
    .B(u0_n_31548),
    .Y(u0_n_31172));
 NAND2xp5_ASAP7_75t_SL u0_g63214 (.A(u0_n_31840),
    .B(u0_n_31526),
    .Y(u0_n_31174));
 NAND2xp5_ASAP7_75t_SL u0_g63215 (.A(u0_n_31826),
    .B(u0_n_31524),
    .Y(u0_n_31176));
 NAND2xp5_ASAP7_75t_SL u0_g63216 (.A(u0_n_33138),
    .B(u0_n_31544),
    .Y(u0_n_31178));
 NOR2xp67_ASAP7_75t_L u0_g63217 (.A(u0_n_32761),
    .B(u0_n_31544),
    .Y(u0_n_31180));
 AND2x2_ASAP7_75t_L u0_g63218 (.A(\u0_w[3] [12]),
    .B(u0_n_31540),
    .Y(u0_n_31182));
 NAND2x1_ASAP7_75t_L u0_g63219 (.A(n_8963),
    .B(u0_n_31549),
    .Y(u0_n_31184));
 NOR2x1_ASAP7_75t_SL u0_g63220 (.A(n_8625),
    .B(u0_n_31546),
    .Y(u0_n_31186));
 INVxp67_ASAP7_75t_R u0_g63221 (.A(u0_n_31232),
    .Y(u0_n_31231));
 INVxp33_ASAP7_75t_R u0_g63222 (.A(u0_n_31235),
    .Y(u0_n_31234));
 INVxp33_ASAP7_75t_R u0_g63223 (.A(u0_n_31242),
    .Y(u0_n_31241));
 INVxp33_ASAP7_75t_R u0_g63224 (.A(u0_n_31246),
    .Y(u0_n_31245));
 INVxp33_ASAP7_75t_R u0_g63225 (.A(u0_n_31254),
    .Y(u0_n_31253));
 INVxp67_ASAP7_75t_L u0_g63226 (.A(u0_n_31265),
    .Y(u0_n_31264));
 INVxp67_ASAP7_75t_R u0_g63227 (.A(u0_n_31267),
    .Y(u0_n_31266));
 INVxp33_ASAP7_75t_R u0_g63228 (.A(u0_n_31272),
    .Y(u0_n_31271));
 INVxp33_ASAP7_75t_R u0_g63229 (.A(u0_n_31273),
    .Y(u0_n_31274));
 INVxp67_ASAP7_75t_R u0_g63230 (.A(u0_n_31279),
    .Y(u0_n_31278));
 INVxp33_ASAP7_75t_R u0_g63231 (.A(u0_n_31281),
    .Y(u0_n_31280));
 INVxp33_ASAP7_75t_R u0_g63232 (.A(u0_n_31282),
    .Y(u0_n_31283));
 INVxp33_ASAP7_75t_R u0_g63233 (.A(u0_n_31285),
    .Y(u0_n_31284));
 INVxp67_ASAP7_75t_R u0_g63234 (.A(u0_n_31288),
    .Y(u0_n_31287));
 INVxp33_ASAP7_75t_R u0_g63235 (.A(u0_n_31290),
    .Y(u0_n_31289));
 INVxp33_ASAP7_75t_R u0_g63236 (.A(u0_n_31291),
    .Y(u0_n_31292));
 INVxp67_ASAP7_75t_R u0_g63237 (.A(u0_n_31294),
    .Y(u0_n_31293));
 INVxp67_ASAP7_75t_SL u0_g63238 (.A(u0_n_31296),
    .Y(u0_n_31295));
 INVxp67_ASAP7_75t_L u0_g63239 (.A(u0_n_31297),
    .Y(u0_n_31298));
 INVxp33_ASAP7_75t_R u0_g63240 (.A(u0_n_31300),
    .Y(u0_n_31299));
 INVxp33_ASAP7_75t_R u0_g63241 (.A(u0_n_31301),
    .Y(u0_n_31302));
 INVxp67_ASAP7_75t_R u0_g63242 (.A(u0_n_31305),
    .Y(u0_n_31304));
 INVxp67_ASAP7_75t_R u0_g63243 (.A(u0_n_31306),
    .Y(u0_n_31307));
 INVxp67_ASAP7_75t_R u0_g63244 (.A(u0_n_31310),
    .Y(u0_n_31309));
 HB1xp67_ASAP7_75t_L u0_g63246 (.A(u0_n_31316),
    .Y(u0_n_31314));
 INVxp33_ASAP7_75t_R u0_g63247 (.A(u0_n_31319),
    .Y(u0_n_31318));
 INVxp67_ASAP7_75t_L u0_g63248 (.A(u0_n_31325),
    .Y(u0_n_31324));
 INVxp33_ASAP7_75t_R u0_g63249 (.A(u0_n_31327),
    .Y(u0_n_31326));
 INVxp33_ASAP7_75t_R u0_g63250 (.A(u0_n_31329),
    .Y(u0_n_31328));
 INVxp67_ASAP7_75t_R u0_g63251 (.A(u0_n_31330),
    .Y(u0_n_31331));
 INVxp33_ASAP7_75t_R u0_g63252 (.A(u0_n_31332),
    .Y(u0_n_31333));
 OAI22xp33_ASAP7_75t_R u0_g63253 (.A1(u0_n_32108),
    .A2(\u0_w[3] [12]),
    .B1(u0_n_31802),
    .B2(n_8801),
    .Y(u0_n_31334));
 OAI221xp5_ASAP7_75t_R u0_g63254 (.A1(u0_n_31830),
    .A2(u0_n_32751),
    .B1(\u0_w[3] [27]),
    .B2(u0_n_32717),
    .C(u0_n_33033),
    .Y(u0_n_31335));
 OAI221xp5_ASAP7_75t_R u0_g63255 (.A1(u0_n_31818),
    .A2(u0_n_32749),
    .B1(w3[11]),
    .B2(w3[15]),
    .C(w3[14]),
    .Y(u0_n_31336));
 NOR2xp33_ASAP7_75t_R u0_g63256 (.A(u0_n_32075),
    .B(u0_n_31434),
    .Y(u0_n_31337));
 NAND2xp33_ASAP7_75t_R u0_g63257 (.A(u0_n_32175),
    .B(u0_n_31502),
    .Y(u0_n_31339));
 NAND2xp33_ASAP7_75t_R u0_g63258 (.A(u0_n_31850),
    .B(u0_n_31625),
    .Y(u0_n_31340));
 NAND2xp33_ASAP7_75t_R u0_g63259 (.A(u0_n_32304),
    .B(u0_n_31628),
    .Y(u0_n_31342));
 NAND2xp33_ASAP7_75t_L u0_g63260 (.A(u0_n_31965),
    .B(u0_n_31662),
    .Y(u0_n_31344));
 NOR2xp33_ASAP7_75t_R u0_g63261 (.A(u0_n_32165),
    .B(u0_n_31546),
    .Y(u0_n_31346));
 OAI21xp33_ASAP7_75t_R u0_g63262 (.A1(u0_n_31954),
    .A2(u0_n_31998),
    .B(u0_n_31934),
    .Y(u0_n_31347));
 AOI21xp33_ASAP7_75t_R u0_g63263 (.A1(u0_n_31795),
    .A2(u0_n_31837),
    .B(u0_n_31875),
    .Y(u0_n_31349));
 AOI21xp33_ASAP7_75t_R u0_g63264 (.A1(u0_n_31826),
    .A2(u0_n_31983),
    .B(u0_n_32108),
    .Y(u0_n_31350));
 AOI21xp33_ASAP7_75t_R u0_g63265 (.A1(u0_n_31895),
    .A2(u0_n_31924),
    .B(u0_n_31639),
    .Y(u0_n_31352));
 OAI21xp33_ASAP7_75t_R u0_g63266 (.A1(n_11346),
    .A2(u0_n_31796),
    .B(u0_n_31895),
    .Y(u0_n_31353));
 OA21x2_ASAP7_75t_R u0_g63267 (.A1(n_8656),
    .A2(u0_n_31822),
    .B(u0_n_31916),
    .Y(u0_n_31354));
 NAND3xp33_ASAP7_75t_R u0_g63268 (.A(u0_n_32175),
    .B(u0_n_31825),
    .C(u0_n_32759),
    .Y(u0_n_31355));
 OAI21xp33_ASAP7_75t_L u0_g63269 (.A1(u0_n_31794),
    .A2(u0_n_32409),
    .B(u0_n_31581),
    .Y(u0_n_31356));
 AOI21xp33_ASAP7_75t_R u0_g63270 (.A1(u0_n_32407),
    .A2(u0_n_31929),
    .B(u0_n_31398),
    .Y(u0_n_31358));
 AOI21xp5_ASAP7_75t_R u0_g63271 (.A1(u0_n_31804),
    .A2(u0_n_32373),
    .B(u0_n_32743),
    .Y(u0_n_31360));
 AOI21xp33_ASAP7_75t_R u0_g63272 (.A1(u0_n_32166),
    .A2(u0_n_31946),
    .B(w3[0]),
    .Y(u0_n_31361));
 NAND2xp5_ASAP7_75t_SL u0_g63273 (.A(u0_n_32084),
    .B(u0_n_31648),
    .Y(u0_n_31232));
 NOR2xp33_ASAP7_75t_R u0_g63274 (.A(u0_n_31817),
    .B(u0_n_31541),
    .Y(u0_n_31363));
 NAND2xp5_ASAP7_75t_L u0_g63275 (.A(u0_n_31983),
    .B(u0_n_31541),
    .Y(u0_n_31233));
 NAND2xp33_ASAP7_75t_R u0_g63276 (.A(u0_n_31546),
    .B(u0_n_31977),
    .Y(u0_n_31235));
 NAND2xp33_ASAP7_75t_R u0_g63277 (.A(u0_n_31548),
    .B(u0_n_31976),
    .Y(u0_n_31236));
 NAND2xp33_ASAP7_75t_R u0_g63278 (.A(u0_n_31985),
    .B(u0_n_31544),
    .Y(u0_n_31237));
 OAI21xp33_ASAP7_75t_R u0_g63279 (.A1(u0_n_31938),
    .A2(u0_n_32344),
    .B(u0_n_31646),
    .Y(u0_n_31238));
 NOR2xp33_ASAP7_75t_R u0_g63280 (.A(u0_n_31680),
    .B(u0_n_31670),
    .Y(u0_n_31239));
 NAND2xp33_ASAP7_75t_R u0_g63281 (.A(u0_n_31685),
    .B(u0_n_31678),
    .Y(u0_n_31240));
 NOR2xp33_ASAP7_75t_L u0_g63282 (.A(u0_n_32083),
    .B(u0_n_31530),
    .Y(u0_n_31242));
 NAND2xp5_ASAP7_75t_R u0_g63283 (.A(u0_n_32122),
    .B(u0_n_31529),
    .Y(u0_n_31243));
 NAND2xp5_ASAP7_75t_L u0_g63284 (.A(u0_n_31986),
    .B(u0_n_31543),
    .Y(u0_n_31244));
 OAI21xp33_ASAP7_75t_R u0_g63285 (.A1(u0_n_31801),
    .A2(u0_n_31814),
    .B(u0_n_32175),
    .Y(u0_n_31246));
 AOI21xp33_ASAP7_75t_R u0_g63286 (.A1(u0_n_31803),
    .A2(u0_n_31805),
    .B(u0_n_32321),
    .Y(u0_n_31247));
 AOI21xp33_ASAP7_75t_R u0_g63287 (.A1(u0_n_31812),
    .A2(u0_n_31807),
    .B(u0_n_32017),
    .Y(u0_n_31248));
 AOI21xp33_ASAP7_75t_R u0_g63288 (.A1(u0_n_31815),
    .A2(u0_n_31809),
    .B(u0_n_31846),
    .Y(u0_n_31249));
 NOR2xp33_ASAP7_75t_R u0_g63289 (.A(u0_n_31661),
    .B(u0_n_31667),
    .Y(u0_n_31250));
 NAND2xp5_ASAP7_75t_R u0_g63290 (.A(u0_n_31669),
    .B(u0_n_31665),
    .Y(u0_n_31251));
 NOR2xp33_ASAP7_75t_R u0_g63291 (.A(u0_n_32165),
    .B(u0_n_31434),
    .Y(u0_n_31252));
 OAI21xp33_ASAP7_75t_R u0_g63292 (.A1(u0_n_31943),
    .A2(u0_n_32272),
    .B(u0_n_31643),
    .Y(u0_n_31254));
 NAND2xp33_ASAP7_75t_R u0_g63293 (.A(n_11516),
    .B(u0_n_31673),
    .Y(u0_n_31255));
 NOR2xp33_ASAP7_75t_SL u0_g63294 (.A(u0_n_31654),
    .B(u0_n_31659),
    .Y(u0_n_31256));
 NAND2xp33_ASAP7_75t_R u0_g63295 (.A(u0_n_31545),
    .B(u0_n_31821),
    .Y(u0_n_31257));
 AO21x1_ASAP7_75t_R u0_g63296 (.A1(n_8625),
    .A2(u0_n_31924),
    .B(u0_n_31838),
    .Y(u0_n_31258));
 NAND2xp5_ASAP7_75t_L u0_g63297 (.A(u0_n_31673),
    .B(u0_n_31837),
    .Y(u0_n_31259));
 OR2x2_ASAP7_75t_L u0_g63298 (.A(u0_n_32409),
    .B(u0_n_31433),
    .Y(u0_n_31260));
 OR2x2_ASAP7_75t_SL u0_g63299 (.A(u0_n_31988),
    .B(u0_n_31650),
    .Y(u0_n_31261));
 NOR2xp33_ASAP7_75t_R u0_g63300 (.A(u0_n_32385),
    .B(u0_n_31413),
    .Y(u0_n_31370));
 NOR2xp33_ASAP7_75t_R u0_g63301 (.A(u0_n_31824),
    .B(u0_n_31537),
    .Y(u0_n_31262));
 NOR2x1_ASAP7_75t_L u0_g63302 (.A(u0_n_31817),
    .B(u0_n_31668),
    .Y(u0_n_31263));
 NOR2xp67_ASAP7_75t_SL u0_g63303 (.A(u0_n_31421),
    .B(u0_n_31822),
    .Y(u0_n_31265));
 NAND2xp33_ASAP7_75t_L u0_g63304 (.A(u0_n_31977),
    .B(u0_n_31532),
    .Y(u0_n_31267));
 NAND2xp5_ASAP7_75t_R u0_g63305 (.A(u0_n_31840),
    .B(u0_n_31531),
    .Y(u0_n_31268));
 NOR2xp67_ASAP7_75t_L u0_g63306 (.A(u0_n_31416),
    .B(u0_n_31680),
    .Y(u0_n_31269));
 NAND2xp5_ASAP7_75t_L u0_g63307 (.A(u0_n_31529),
    .B(u0_n_31826),
    .Y(u0_n_31270));
 NOR2xp33_ASAP7_75t_SL u0_g63308 (.A(u0_n_31421),
    .B(u0_n_31684),
    .Y(u0_n_31272));
 NAND2xp5_ASAP7_75t_L u0_g63309 (.A(u0_n_31827),
    .B(u0_n_31660),
    .Y(u0_n_31273));
 NOR2xp33_ASAP7_75t_L u0_g63310 (.A(u0_n_31944),
    .B(u0_n_31654),
    .Y(u0_n_31275));
 NAND2xp5_ASAP7_75t_R u0_g63311 (.A(n_11516),
    .B(u0_n_31945),
    .Y(u0_n_31276));
 NOR2xp33_ASAP7_75t_R u0_g63312 (.A(u0_n_31975),
    .B(u0_n_31682),
    .Y(u0_n_31277));
 NAND2xp33_ASAP7_75t_R u0_g63313 (.A(u0_n_32040),
    .B(u0_n_31536),
    .Y(u0_n_31279));
 AND2x2_ASAP7_75t_SL u0_g63314 (.A(u0_n_31972),
    .B(u0_n_31497),
    .Y(u0_n_31281));
 AND2x2_ASAP7_75t_SL u0_g63315 (.A(u0_n_31821),
    .B(u0_n_31666),
    .Y(u0_n_31282));
 NOR2xp33_ASAP7_75t_L u0_g63316 (.A(u0_n_31951),
    .B(u0_n_31502),
    .Y(u0_n_31285));
 NAND2xp5_ASAP7_75t_L u0_g63317 (.A(u0_n_31665),
    .B(u0_n_31938),
    .Y(u0_n_31286));
 NAND2xp5_ASAP7_75t_R u0_g63318 (.A(u0_n_31535),
    .B(u0_n_31985),
    .Y(u0_n_31288));
 NAND2xp5_ASAP7_75t_R u0_g63319 (.A(u0_n_31543),
    .B(u0_n_31819),
    .Y(u0_n_31290));
 NAND2xp33_ASAP7_75t_R u0_g63320 (.A(u0_n_31546),
    .B(u0_n_31841),
    .Y(u0_n_31291));
 NOR2xp33_ASAP7_75t_SL u0_g63321 (.A(u0_n_31962),
    .B(u0_n_31661),
    .Y(u0_n_31294));
 NAND2xp5_ASAP7_75t_SL u0_g63322 (.A(u0_n_31607),
    .B(u0_n_32040),
    .Y(u0_n_31296));
 NAND2xp5_ASAP7_75t_SL u0_g63323 (.A(u0_n_31610),
    .B(u0_n_32113),
    .Y(u0_n_31297));
 NOR2xp33_ASAP7_75t_L u0_g63324 (.A(u0_n_32174),
    .B(u0_n_31540),
    .Y(u0_n_31300));
 NOR2xp33_ASAP7_75t_L u0_g63325 (.A(u0_n_31676),
    .B(u0_n_31533),
    .Y(u0_n_31301));
 NAND2xp5_ASAP7_75t_R u0_g63326 (.A(u0_n_31538),
    .B(u0_n_31983),
    .Y(u0_n_31303));
 NAND2xp5_ASAP7_75t_SL u0_g63327 (.A(u0_n_31675),
    .B(u0_n_31538),
    .Y(u0_n_31305));
 NAND2xp5_ASAP7_75t_SL u0_g63328 (.A(u0_n_31535),
    .B(u0_n_31678),
    .Y(u0_n_31306));
 NOR2xp33_ASAP7_75t_SL u0_g63329 (.A(u0_n_31545),
    .B(u0_n_32011),
    .Y(u0_n_31308));
 NOR2xp33_ASAP7_75t_SL u0_g63330 (.A(u0_n_31670),
    .B(u0_n_31682),
    .Y(u0_n_31310));
 NOR2xp33_ASAP7_75t_R u0_g63331 (.A(u0_n_32306),
    .B(u0_n_31549),
    .Y(u0_n_31311));
 AOI21xp5_ASAP7_75t_L u0_g63332 (.A1(u0_n_31821),
    .A2(u0_n_32735),
    .B(u0_n_31684),
    .Y(u0_n_31312));
 AOI21xp5_ASAP7_75t_L u0_g63333 (.A1(u0_n_31983),
    .A2(n_8856),
    .B(u0_n_31507),
    .Y(u0_n_31313));
 AOI21xp5_ASAP7_75t_SL u0_g63334 (.A1(u0_n_31977),
    .A2(w3[1]),
    .B(u0_n_31503),
    .Y(u0_n_31316));
 OA21x2_ASAP7_75t_SL u0_g63335 (.A1(u0_n_32735),
    .A2(u0_n_31984),
    .B(u0_n_31500),
    .Y(u0_n_31317));
 OAI21xp33_ASAP7_75t_L u0_g63336 (.A1(u0_n_32706),
    .A2(u0_n_31975),
    .B(u0_n_31491),
    .Y(u0_n_31319));
 OAI21xp5_ASAP7_75t_L u0_g63337 (.A1(n_8747),
    .A2(u0_n_31838),
    .B(u0_n_31461),
    .Y(u0_n_31320));
 AOI21xp5_ASAP7_75t_SL u0_g63338 (.A1(u0_n_31818),
    .A2(n_8856),
    .B(u0_n_31488),
    .Y(u0_n_31322));
 AOI21xp33_ASAP7_75t_SL u0_g63339 (.A1(u0_n_31827),
    .A2(u0_n_32704),
    .B(u0_n_31483),
    .Y(u0_n_31323));
 NAND2xp5_ASAP7_75t_R u0_g63340 (.A(u0_n_31669),
    .B(u0_n_31529),
    .Y(u0_n_31325));
 NOR2xp33_ASAP7_75t_SL u0_g63341 (.A(u0_n_31530),
    .B(u0_n_31672),
    .Y(u0_n_31327));
 NOR2xp33_ASAP7_75t_L u0_g63342 (.A(u0_n_31667),
    .B(u0_n_31542),
    .Y(u0_n_31329));
 NOR2xp67_ASAP7_75t_L u0_g63343 (.A(u0_n_31659),
    .B(u0_n_31537),
    .Y(u0_n_31330));
 OAI21xp33_ASAP7_75t_R u0_g63344 (.A1(u0_r0_rcnt[2]),
    .A2(u0_n_31749),
    .B(u0_n_31448),
    .Y(u0_n_31332));
 INVxp33_ASAP7_75t_R u0_g63345 (.A(u0_n_31394),
    .Y(u0_n_31393));
 INVxp33_ASAP7_75t_R u0_g63346 (.A(u0_n_31408),
    .Y(u0_n_31407));
 INVxp33_ASAP7_75t_R u0_g63347 (.A(u0_n_31411),
    .Y(u0_n_31412));
 INVxp33_ASAP7_75t_R u0_g63348 (.A(u0_n_31414),
    .Y(u0_n_31413));
 INVxp67_ASAP7_75t_R u0_g63349 (.A(u0_n_31416),
    .Y(u0_n_31415));
 INVxp33_ASAP7_75t_R u0_g63350 (.A(u0_n_31419),
    .Y(u0_n_31420));
 INVxp67_ASAP7_75t_R u0_g63351 (.A(u0_n_31422),
    .Y(u0_n_31423));
 INVxp33_ASAP7_75t_R u0_g63352 (.A(u0_n_31427),
    .Y(u0_n_31428));
 INVxp33_ASAP7_75t_R u0_g63353 (.A(u0_n_31430),
    .Y(u0_n_31429));
 INVxp67_ASAP7_75t_R u0_g63354 (.A(u0_n_31437),
    .Y(u0_n_31436));
 INVxp33_ASAP7_75t_R u0_g63355 (.A(u0_n_31439),
    .Y(u0_n_31438));
 INVxp67_ASAP7_75t_R u0_g63356 (.A(u0_n_31442),
    .Y(u0_n_31441));
 INVxp33_ASAP7_75t_R u0_g63357 (.A(u0_n_31445),
    .Y(u0_n_31446));
 INVxp33_ASAP7_75t_R u0_g63358 (.A(u0_n_31451),
    .Y(u0_n_31452));
 INVxp33_ASAP7_75t_R u0_g63359 (.A(u0_n_31454),
    .Y(u0_n_31455));
 INVxp67_ASAP7_75t_R u0_g63360 (.A(u0_n_31456),
    .Y(u0_n_31457));
 INVxp67_ASAP7_75t_R u0_g63361 (.A(u0_n_31459),
    .Y(u0_n_31460));
 INVxp33_ASAP7_75t_R u0_g63362 (.A(u0_n_31463),
    .Y(u0_n_31462));
 INVxp33_ASAP7_75t_R u0_g63363 (.A(u0_n_31467),
    .Y(u0_n_31466));
 INVxp67_ASAP7_75t_R u0_g63364 (.A(u0_n_31468),
    .Y(u0_n_31469));
 INVxp67_ASAP7_75t_R u0_g63365 (.A(u0_n_31474),
    .Y(u0_n_31475));
 INVxp67_ASAP7_75t_R u0_g63366 (.A(u0_n_31477),
    .Y(u0_n_31478));
 INVxp67_ASAP7_75t_R u0_g63367 (.A(u0_n_31481),
    .Y(u0_n_31480));
 INVxp67_ASAP7_75t_R u0_g63368 (.A(u0_n_31483),
    .Y(u0_n_31482));
 INVxp33_ASAP7_75t_R u0_g63369 (.A(u0_n_31485),
    .Y(u0_n_31486));
 INVxp33_ASAP7_75t_R u0_g63370 (.A(u0_n_31488),
    .Y(u0_n_31487));
 INVxp67_ASAP7_75t_R u0_g63371 (.A(u0_n_31491),
    .Y(u0_n_31492));
 INVx1_ASAP7_75t_R u0_g63372 (.A(u0_n_31494),
    .Y(u0_n_31493));
 INVx1_ASAP7_75t_L u0_g63373 (.A(u0_n_31495),
    .Y(u0_n_31496));
 INVxp33_ASAP7_75t_R u0_g63374 (.A(u0_n_31497),
    .Y(u0_n_31498));
 INVxp67_ASAP7_75t_R u0_g63375 (.A(u0_n_31500),
    .Y(u0_n_31501));
 INVxp33_ASAP7_75t_R u0_g63377 (.A(u0_n_31503),
    .Y(u0_n_31504));
 INVxp67_ASAP7_75t_R u0_g63379 (.A(u0_n_31507),
    .Y(u0_n_31508));
 INVxp67_ASAP7_75t_R u0_g63380 (.A(u0_n_31510),
    .Y(u0_n_31509));
 INVxp33_ASAP7_75t_R u0_g63381 (.A(u0_n_31512),
    .Y(u0_n_31513));
 INVxp33_ASAP7_75t_R u0_g63382 (.A(u0_n_31514),
    .Y(u0_n_31515));
 INVxp33_ASAP7_75t_R u0_g63383 (.A(u0_n_31516),
    .Y(u0_n_31517));
 INVx1_ASAP7_75t_SL u0_g63384 (.A(u0_n_31518),
    .Y(u0_n_31519));
 INVx1_ASAP7_75t_R u0_g63385 (.A(u0_n_31520),
    .Y(u0_n_31521));
 INVxp33_ASAP7_75t_R u0_g63386 (.A(u0_n_31522),
    .Y(u0_n_31523));
 INVxp67_ASAP7_75t_L u0_g63387 (.A(u0_n_31524),
    .Y(u0_n_31525));
 INVxp33_ASAP7_75t_R u0_g63388 (.A(u0_n_31526),
    .Y(u0_n_31527));
 INVx1_ASAP7_75t_SL u0_g63389 (.A(u0_n_31528),
    .Y(u0_n_31529));
 INVx1_ASAP7_75t_SL u0_g63390 (.A(u0_n_31530),
    .Y(u0_n_31531));
 INVx1_ASAP7_75t_L u0_g63391 (.A(u0_n_31532),
    .Y(u0_n_31533));
 INVx1_ASAP7_75t_SL u0_g63392 (.A(u0_n_31534),
    .Y(u0_n_31535));
 INVx1_ASAP7_75t_R u0_g63393 (.A(u0_n_31536),
    .Y(u0_n_31537));
 INVx1_ASAP7_75t_SL u0_g63394 (.A(u0_n_31538),
    .Y(u0_n_31539));
 INVx1_ASAP7_75t_SL u0_g63395 (.A(u0_n_31540),
    .Y(u0_n_31541));
 INVx1_ASAP7_75t_R u0_g63396 (.A(u0_n_31542),
    .Y(u0_n_31543));
 INVx1_ASAP7_75t_R u0_g63397 (.A(u0_n_31544),
    .Y(u0_n_31545));
 INVx1_ASAP7_75t_SL u0_g63398 (.A(u0_n_31546),
    .Y(u0_n_31547));
 INVx2_ASAP7_75t_L u0_g63399 (.A(u0_n_31548),
    .Y(u0_n_31549));
 NAND2xp33_ASAP7_75t_R u0_g63400 (.A(u0_n_32763),
    .B(u0_n_31748),
    .Y(u0_n_31550));
 NOR2xp33_ASAP7_75t_R u0_g63401 (.A(u0_n_31747),
    .B(u0_n_31816),
    .Y(u0_n_31551));
 NOR2xp33_ASAP7_75t_R u0_g63402 (.A(w3[19]),
    .B(u0_n_31953),
    .Y(u0_n_31552));
 NOR2xp33_ASAP7_75t_R u0_g63403 (.A(u0_n_31753),
    .B(u0_n_31811),
    .Y(u0_n_31553));
 NAND2xp33_ASAP7_75t_R u0_g63404 (.A(n_8748),
    .B(u0_n_31895),
    .Y(u0_n_31388));
 NAND2xp33_ASAP7_75t_R u0_g63405 (.A(w3[21]),
    .B(u0_n_31957),
    .Y(u0_n_31389));
 NOR2xp33_ASAP7_75t_R u0_g63406 (.A(w3[21]),
    .B(u0_n_31949),
    .Y(u0_n_31390));
 NAND2xp33_ASAP7_75t_R u0_g63407 (.A(u0_n_31819),
    .B(u0_n_31821),
    .Y(u0_n_31391));
 NOR2xp33_ASAP7_75t_R u0_g63408 (.A(u0_n_31825),
    .B(u0_n_31817),
    .Y(u0_n_31392));
 NOR2xp33_ASAP7_75t_R u0_g63409 (.A(u0_n_32735),
    .B(u0_n_32209),
    .Y(u0_n_31394));
 NOR2xp33_ASAP7_75t_L u0_g63410 (.A(w3[15]),
    .B(u0_n_31969),
    .Y(u0_n_31395));
 NAND2xp33_ASAP7_75t_R u0_g63411 (.A(u0_n_32704),
    .B(u0_n_32273),
    .Y(u0_n_31396));
 NOR2xp33_ASAP7_75t_SL u0_g63412 (.A(n_11346),
    .B(u0_n_31964),
    .Y(u0_n_31397));
 NOR2xp33_ASAP7_75t_R u0_g63413 (.A(n_8851),
    .B(u0_n_32338),
    .Y(u0_n_31398));
 NAND2xp5_ASAP7_75t_L u0_g63414 (.A(u0_n_32716),
    .B(u0_n_31959),
    .Y(u0_n_31399));
 NAND2xp5_ASAP7_75t_L u0_g63415 (.A(w3[17]),
    .B(u0_n_31808),
    .Y(u0_n_31400));
 NOR2xp33_ASAP7_75t_SL u0_g63416 (.A(u0_n_32704),
    .B(u0_n_32372),
    .Y(u0_n_31401));
 NOR2xp33_ASAP7_75t_SL u0_g63417 (.A(n_8831),
    .B(u0_n_31988),
    .Y(u0_n_31402));
 NAND2xp33_ASAP7_75t_R u0_g63418 (.A(n_11507),
    .B(u0_n_31967),
    .Y(u0_n_31403));
 NAND2xp5_ASAP7_75t_R u0_g63419 (.A(n_8831),
    .B(u0_n_32208),
    .Y(u0_n_31404));
 NAND2xp33_ASAP7_75t_R u0_g63420 (.A(w3[5]),
    .B(u0_n_31790),
    .Y(u0_n_31405));
 NAND2xp5_ASAP7_75t_R u0_g63421 (.A(w3[29]),
    .B(u0_n_31973),
    .Y(u0_n_31406));
 NAND2xp33_ASAP7_75t_R u0_g63422 (.A(w3[29]),
    .B(u0_n_31798),
    .Y(u0_n_31408));
 NAND2xp5_ASAP7_75t_R u0_g63423 (.A(u0_n_32012),
    .B(u0_n_32753),
    .Y(u0_n_31409));
 NAND2xp33_ASAP7_75t_R u0_g63424 (.A(w3[2]),
    .B(u0_n_31841),
    .Y(u0_n_31410));
 NAND2xp33_ASAP7_75t_R u0_g63425 (.A(w3[13]),
    .B(u0_n_31955),
    .Y(u0_n_31411));
 NAND2xp33_ASAP7_75t_R u0_g63426 (.A(u0_n_31781),
    .B(u0_n_31805),
    .Y(u0_n_31414));
 NOR2xp33_ASAP7_75t_L u0_g63427 (.A(n_8963),
    .B(u0_n_31781),
    .Y(u0_n_31416));
 NAND2xp5_ASAP7_75t_L u0_g63428 (.A(u0_n_32012),
    .B(w3[18]),
    .Y(u0_n_31417));
 NOR2xp33_ASAP7_75t_L u0_g63429 (.A(u0_n_31814),
    .B(n_8856),
    .Y(u0_n_31418));
 NOR2xp33_ASAP7_75t_R u0_g63430 (.A(w3[5]),
    .B(u0_n_31941),
    .Y(u0_n_31419));
 NOR2xp67_ASAP7_75t_L u0_g63431 (.A(w3[20]),
    .B(u0_n_31785),
    .Y(u0_n_31421));
 NOR2xp33_ASAP7_75t_L u0_g63432 (.A(u0_n_32697),
    .B(u0_n_32083),
    .Y(u0_n_31422));
 NOR2xp33_ASAP7_75t_SL u0_g63433 (.A(u0_n_31810),
    .B(w3[1]),
    .Y(u0_n_31424));
 NAND2xp33_ASAP7_75t_R u0_g63434 (.A(w3[15]),
    .B(u0_n_32339),
    .Y(u0_n_31425));
 NAND2xp33_ASAP7_75t_R u0_g63435 (.A(w3[2]),
    .B(u0_n_32142),
    .Y(u0_n_31426));
 NAND2xp5_ASAP7_75t_R u0_g63436 (.A(u0_n_32717),
    .B(u0_n_32273),
    .Y(u0_n_31427));
 NOR2xp33_ASAP7_75t_L u0_g63437 (.A(u0_n_32706),
    .B(u0_n_31971),
    .Y(u0_n_31430));
 NAND2xp5_ASAP7_75t_R u0_g63438 (.A(u0_n_32706),
    .B(u0_n_31803),
    .Y(u0_n_31431));
 NAND2xp33_ASAP7_75t_R u0_g63439 (.A(w3[21]),
    .B(u0_n_31788),
    .Y(u0_n_31432));
 NOR2xp33_ASAP7_75t_R u0_g63440 (.A(u0_n_31776),
    .B(u0_n_31801),
    .Y(u0_n_31433));
 NOR2xp33_ASAP7_75t_L u0_g63441 (.A(u0_n_31772),
    .B(u0_n_31816),
    .Y(u0_n_31434));
 NOR2xp33_ASAP7_75t_R u0_g63442 (.A(u0_n_32753),
    .B(u0_n_32254),
    .Y(u0_n_31435));
 NOR2xp33_ASAP7_75t_SL u0_g63443 (.A(w3[9]),
    .B(u0_n_31813),
    .Y(u0_n_31437));
 NOR2xp33_ASAP7_75t_R u0_g63444 (.A(u0_n_32743),
    .B(u0_n_32372),
    .Y(u0_n_31439));
 NOR2xp33_ASAP7_75t_R u0_g63445 (.A(w3[24]),
    .B(u0_n_32306),
    .Y(u0_n_31440));
 NOR2xp33_ASAP7_75t_L u0_g63446 (.A(u0_n_32745),
    .B(u0_n_32410),
    .Y(u0_n_31442));
 NOR2xp33_ASAP7_75t_R u0_g63447 (.A(u0_n_32747),
    .B(u0_n_32160),
    .Y(u0_n_31443));
 NOR2xp33_ASAP7_75t_R u0_g63448 (.A(n_11401),
    .B(u0_n_32174),
    .Y(u0_n_31444));
 NAND2xp5_ASAP7_75t_R u0_g63449 (.A(u0_n_31812),
    .B(u0_n_31819),
    .Y(u0_n_31445));
 NOR2xp33_ASAP7_75t_R u0_g63450 (.A(u0_n_31783),
    .B(u0_n_32685),
    .Y(u0_n_31447));
 NAND2xp33_ASAP7_75t_R u0_g63451 (.A(u0_r0_rcnt[2]),
    .B(u0_n_31749),
    .Y(u0_n_31448));
 AND2x2_ASAP7_75t_L u0_g63452 (.A(u0_n_32698),
    .B(u0_n_31971),
    .Y(u0_n_31449));
 NOR2xp33_ASAP7_75t_SL u0_g63453 (.A(w3[20]),
    .B(u0_n_31918),
    .Y(u0_n_31450));
 NAND2xp5_ASAP7_75t_R u0_g63454 (.A(n_11401),
    .B(u0_n_31764),
    .Y(u0_n_31451));
 NAND2xp5_ASAP7_75t_R u0_g63455 (.A(u0_n_32689),
    .B(u0_n_31973),
    .Y(u0_n_31454));
 NOR2xp33_ASAP7_75t_SL u0_g63456 (.A(w3[1]),
    .B(u0_n_31809),
    .Y(u0_n_31456));
 NAND2xp5_ASAP7_75t_R u0_g63457 (.A(w3[24]),
    .B(u0_n_31751),
    .Y(u0_n_31458));
 NAND2xp5_ASAP7_75t_R u0_g63458 (.A(w3[0]),
    .B(u0_n_31841),
    .Y(u0_n_31459));
 NAND2xp5_ASAP7_75t_L u0_g63459 (.A(n_8747),
    .B(u0_n_31838),
    .Y(u0_n_31461));
 NAND2xp5_ASAP7_75t_L u0_g63460 (.A(w3[17]),
    .B(u0_n_31953),
    .Y(u0_n_31463));
 NOR2xp67_ASAP7_75t_L u0_g63461 (.A(u0_n_31838),
    .B(u0_n_31772),
    .Y(u0_n_31464));
 NAND2xp5_ASAP7_75t_R u0_g63462 (.A(u0_n_31785),
    .B(u0_n_31812),
    .Y(u0_n_31465));
 NAND2xp5_ASAP7_75t_L u0_g63463 (.A(u0_n_31815),
    .B(u0_n_31840),
    .Y(u0_n_31467));
 NAND2xp5_ASAP7_75t_L u0_g63464 (.A(\u0_w[3] [16]),
    .B(u0_n_32012),
    .Y(u0_n_31468));
 NOR2xp33_ASAP7_75t_SL u0_g63465 (.A(u0_n_31926),
    .B(w3[12]),
    .Y(u0_n_31470));
 NAND2xp5_ASAP7_75t_R u0_g63466 (.A(w3[9]),
    .B(u0_n_31813),
    .Y(u0_n_31471));
 NAND2xp5_ASAP7_75t_L u0_g63467 (.A(n_8851),
    .B(u0_n_31951),
    .Y(u0_n_31473));
 NAND2xp5_ASAP7_75t_R u0_g63468 (.A(n_11401),
    .B(u0_n_32193),
    .Y(u0_n_31474));
 NAND2xp5_ASAP7_75t_L u0_g63469 (.A(w3[24]),
    .B(u0_n_32308),
    .Y(u0_n_31477));
 AND2x2_ASAP7_75t_L u0_g63470 (.A(u0_n_32685),
    .B(u0_n_31955),
    .Y(u0_n_31479));
 NAND2xp5_ASAP7_75t_L u0_g63471 (.A(u0_n_32735),
    .B(u0_n_31807),
    .Y(u0_n_31481));
 NOR2xp33_ASAP7_75t_SL u0_g63472 (.A(w3[25]),
    .B(u0_n_31827),
    .Y(u0_n_31483));
 NOR2x1_ASAP7_75t_SL u0_g63473 (.A(w3[4]),
    .B(u0_n_31924),
    .Y(u0_n_31484));
 NAND2xp5_ASAP7_75t_SL u0_g63474 (.A(u0_n_31823),
    .B(u0_n_31805),
    .Y(u0_n_31485));
 NOR2xp33_ASAP7_75t_SL u0_g63475 (.A(n_8856),
    .B(u0_n_31818),
    .Y(u0_n_31488));
 NOR2xp33_ASAP7_75t_L u0_g63476 (.A(u0_n_31822),
    .B(u0_n_31786),
    .Y(u0_n_31489));
 NAND2xp5_ASAP7_75t_L u0_g63477 (.A(u0_n_32698),
    .B(u0_n_31975),
    .Y(u0_n_31491));
 NAND2xp5_ASAP7_75t_SL u0_g63478 (.A(u0_n_32735),
    .B(u0_n_31954),
    .Y(u0_n_31494));
 NAND2xp5_ASAP7_75t_SL u0_g63479 (.A(u0_n_32691),
    .B(u0_n_31967),
    .Y(u0_n_31495));
 NAND2xp5_ASAP7_75t_SL u0_g63480 (.A(u0_n_31827),
    .B(u0_n_31781),
    .Y(u0_n_31497));
 NOR2xp67_ASAP7_75t_L u0_g63481 (.A(u0_n_31937),
    .B(w3[1]),
    .Y(u0_n_31499));
 NAND2x1_ASAP7_75t_SL u0_g63482 (.A(u0_n_32735),
    .B(u0_n_31984),
    .Y(u0_n_31500));
 AND2x2_ASAP7_75t_L u0_g63483 (.A(u0_n_31818),
    .B(u0_n_31775),
    .Y(u0_n_31502));
 NOR2xp67_ASAP7_75t_L u0_g63484 (.A(w3[1]),
    .B(u0_n_31981),
    .Y(u0_n_31503));
 AND2x2_ASAP7_75t_SL u0_g63485 (.A(n_8851),
    .B(u0_n_31982),
    .Y(u0_n_31507));
 NAND2x1_ASAP7_75t_L u0_g63486 (.A(u0_n_32731),
    .B(u0_n_31957),
    .Y(u0_n_31510));
 NOR2xp33_ASAP7_75t_SL u0_g63487 (.A(u0_n_31787),
    .B(w3[21]),
    .Y(u0_n_31512));
 NOR2xp33_ASAP7_75t_SL u0_g63488 (.A(w3[5]),
    .B(u0_n_31789),
    .Y(u0_n_31514));
 NOR2xp67_ASAP7_75t_R u0_g63490 (.A(w3[29]),
    .B(u0_n_31797),
    .Y(u0_n_31516));
 NOR2xp33_ASAP7_75t_SL u0_g63491 (.A(u0_n_31782),
    .B(n_8942),
    .Y(u0_n_31518));
 NOR2xp33_ASAP7_75t_SL u0_g63492 (.A(w3[13]),
    .B(u0_n_31783),
    .Y(u0_n_31520));
 AND2x2_ASAP7_75t_L u0_g63493 (.A(u0_n_33138),
    .B(u0_n_31785),
    .Y(u0_n_31522));
 AND2x2_ASAP7_75t_SL u0_g63494 (.A(u0_n_32759),
    .B(u0_n_31775),
    .Y(u0_n_31524));
 AND2x2_ASAP7_75t_SL u0_g63495 (.A(n_8625),
    .B(u0_n_31773),
    .Y(u0_n_31526));
 NOR2x1_ASAP7_75t_SL u0_g63496 (.A(u0_n_32759),
    .B(u0_n_31776),
    .Y(u0_n_31528));
 NOR2x1_ASAP7_75t_SL u0_g63497 (.A(n_8623),
    .B(u0_n_31772),
    .Y(u0_n_31530));
 NAND2xp5_ASAP7_75t_L u0_g63498 (.A(w3[4]),
    .B(u0_n_31945),
    .Y(u0_n_31532));
 NOR2x1_ASAP7_75t_SL u0_g63499 (.A(u0_n_32761),
    .B(u0_n_31962),
    .Y(u0_n_31534));
 OR2x2_ASAP7_75t_SL u0_g63500 (.A(n_8964),
    .B(u0_n_31782),
    .Y(u0_n_31536));
 NAND2xp5_ASAP7_75t_SL u0_g63501 (.A(\u0_w[3] [12]),
    .B(u0_n_31938),
    .Y(u0_n_31538));
 NAND2x1_ASAP7_75t_SL u0_g63502 (.A(u0_n_31775),
    .B(u0_n_31826),
    .Y(u0_n_31540));
 AND2x2_ASAP7_75t_SL u0_g63503 (.A(w3[20]),
    .B(u0_n_31785),
    .Y(u0_n_31542));
 AND2x4_ASAP7_75t_SL u0_g63504 (.A(u0_n_31819),
    .B(u0_n_31785),
    .Y(u0_n_31544));
 NOR2x1_ASAP7_75t_SL u0_g63505 (.A(u0_n_31772),
    .B(u0_n_31839),
    .Y(u0_n_31546));
 AND2x4_ASAP7_75t_SL u0_g63506 (.A(u0_n_31823),
    .B(u0_n_31781),
    .Y(u0_n_31548));
 INVxp33_ASAP7_75t_R u0_g63507 (.A(u0_n_31572),
    .Y(u0_n_31571));
 INVxp33_ASAP7_75t_R u0_g63508 (.A(u0_n_31578),
    .Y(u0_n_31577));
 INVxp33_ASAP7_75t_R u0_g63509 (.A(u0_n_31580),
    .Y(u0_n_31579));
 INVxp33_ASAP7_75t_R u0_g63510 (.A(u0_n_31586),
    .Y(u0_n_31585));
 INVxp33_ASAP7_75t_R u0_g63511 (.A(u0_n_31590),
    .Y(u0_n_31589));
 INVxp33_ASAP7_75t_R u0_g63512 (.A(u0_n_31594),
    .Y(u0_n_31593));
 INVxp33_ASAP7_75t_R u0_g63513 (.A(u0_n_31596),
    .Y(u0_n_31595));
 INVxp67_ASAP7_75t_R u0_g63514 (.A(u0_n_31598),
    .Y(u0_n_31597));
 INVxp33_ASAP7_75t_R u0_g63515 (.A(u0_n_31600),
    .Y(u0_n_31601));
 INVxp33_ASAP7_75t_R u0_g63516 (.A(u0_n_31602),
    .Y(u0_n_31603));
 INVxp33_ASAP7_75t_R u0_g63517 (.A(u0_n_31605),
    .Y(u0_n_31604));
 INVxp33_ASAP7_75t_R u0_g63518 (.A(u0_n_31609),
    .Y(u0_n_31608));
 INVxp33_ASAP7_75t_R u0_g63519 (.A(u0_n_31612),
    .Y(u0_n_31611));
 INVxp33_ASAP7_75t_R u0_g63520 (.A(u0_n_31614),
    .Y(u0_n_31613));
 INVxp33_ASAP7_75t_R u0_g63521 (.A(u0_n_31616),
    .Y(u0_n_31615));
 INVx1_ASAP7_75t_L u0_g63522 (.A(u0_n_31618),
    .Y(u0_n_31617));
 INVxp33_ASAP7_75t_R u0_g63523 (.A(u0_n_31620),
    .Y(u0_n_31619));
 INVxp33_ASAP7_75t_R u0_g63524 (.A(u0_n_31623),
    .Y(u0_n_31622));
 INVxp33_ASAP7_75t_R u0_g63525 (.A(u0_n_31625),
    .Y(u0_n_31626));
 INVxp67_ASAP7_75t_R u0_g63526 (.A(u0_n_31629),
    .Y(u0_n_31628));
 INVxp33_ASAP7_75t_R u0_g63527 (.A(u0_n_31631),
    .Y(u0_n_31630));
 INVxp33_ASAP7_75t_R u0_g63528 (.A(u0_n_31635),
    .Y(u0_n_31634));
 INVxp33_ASAP7_75t_R u0_g63529 (.A(u0_n_31637),
    .Y(u0_n_31636));
 INVxp33_ASAP7_75t_R u0_g63530 (.A(u0_n_31639),
    .Y(u0_n_31640));
 INVxp33_ASAP7_75t_R u0_g63532 (.A(u0_n_31644),
    .Y(u0_n_31645));
 INVxp67_ASAP7_75t_R u0_g63533 (.A(u0_n_31646),
    .Y(u0_n_31647));
 INVxp67_ASAP7_75t_R u0_g63534 (.A(u0_n_31648),
    .Y(u0_n_31649));
 INVxp33_ASAP7_75t_R u0_g63535 (.A(n_11516),
    .Y(u0_n_31653));
 INVxp33_ASAP7_75t_R u0_g63536 (.A(u0_n_31654),
    .Y(u0_n_31655));
 INVxp33_ASAP7_75t_R u0_g63537 (.A(u0_n_31657),
    .Y(u0_n_31656));
 INVx1_ASAP7_75t_L u0_g63538 (.A(u0_n_31660),
    .Y(u0_n_31659));
 INVxp67_ASAP7_75t_L u0_g63539 (.A(u0_n_31661),
    .Y(u0_n_31662));
 INVxp33_ASAP7_75t_R u0_g63540 (.A(n_11520),
    .Y(u0_n_31664));
 INVxp67_ASAP7_75t_R u0_g63541 (.A(u0_n_31666),
    .Y(u0_n_31667));
 INVxp67_ASAP7_75t_SL u0_g63542 (.A(u0_n_31668),
    .Y(u0_n_31669));
 INVxp67_ASAP7_75t_L u0_g63543 (.A(u0_n_31670),
    .Y(u0_n_31671));
 INVx1_ASAP7_75t_L u0_g63544 (.A(u0_n_31672),
    .Y(u0_n_31673));
 INVxp67_ASAP7_75t_SL u0_g63545 (.A(u0_n_31674),
    .Y(u0_n_31675));
 INVxp33_ASAP7_75t_R u0_g63546 (.A(u0_n_31676),
    .Y(u0_n_31677));
 INVxp33_ASAP7_75t_R u0_g63547 (.A(u0_n_31678),
    .Y(u0_n_31679));
 INVxp67_ASAP7_75t_SL u0_g63548 (.A(u0_n_31680),
    .Y(u0_n_31681));
 INVx1_ASAP7_75t_R u0_g63549 (.A(u0_n_31682),
    .Y(u0_n_31683));
 INVx1_ASAP7_75t_SL u0_g63550 (.A(u0_n_31684),
    .Y(u0_n_31685));
 INVxp67_ASAP7_75t_R u0_g63551 (.A(u0_n_31686),
    .Y(u0_n_31687));
 INVx1_ASAP7_75t_L u0_g63552 (.A(u0_n_31688),
    .Y(u0_n_31689));
 NOR2xp33_ASAP7_75t_R u0_g63553 (.A(u0_n_31800),
    .B(u0_n_32209),
    .Y(u0_n_31690));
 NOR2xp33_ASAP7_75t_R u0_g63554 (.A(u0_n_31811),
    .B(u0_n_31984),
    .Y(u0_n_31691));
 NOR2xp33_ASAP7_75t_R u0_g63555 (.A(u0_n_31820),
    .B(u0_n_31984),
    .Y(u0_n_31692));
 XOR2xp5_ASAP7_75t_R u0_g63556 (.A(w1[11]),
    .B(w2[11]),
    .Y(u0_n_31693));
 XOR2xp5_ASAP7_75t_R u0_g63557 (.A(w1[9]),
    .B(w0[9]),
    .Y(u0_n_31694));
 XOR2xp5_ASAP7_75t_R u0_g63558 (.A(w1[12]),
    .B(w0[12]),
    .Y(u0_n_31696));
 NAND2xp33_ASAP7_75t_R u0_g63559 (.A(u0_n_32759),
    .B(u0_n_31926),
    .Y(u0_n_31568));
 XNOR2xp5_ASAP7_75t_R u0_g63560 (.A(w1[19]),
    .B(w2[19]),
    .Y(u0_n_31698));
 XNOR2xp5_ASAP7_75t_R u0_g63561 (.A(w1[6]),
    .B(w2[6]),
    .Y(u0_n_31700));
 XOR2xp5_ASAP7_75t_R u0_g63562 (.A(w2[7]),
    .B(w1[7]),
    .Y(u0_n_31702));
 XOR2xp5_ASAP7_75t_R u0_g63563 (.A(w2[22]),
    .B(w1[22]),
    .Y(u0_n_31704));
 XOR2xp5_ASAP7_75t_R u0_g63564 (.A(w1[10]),
    .B(w0[10]),
    .Y(u0_n_31706));
 XOR2xp5_ASAP7_75t_R u0_g63565 (.A(w1[1]),
    .B(w0[1]),
    .Y(u0_n_31707));
 XNOR2xp5_ASAP7_75t_R u0_g63566 (.A(w1[30]),
    .B(w2[30]),
    .Y(u0_n_31709));
 NAND2xp33_ASAP7_75t_R u0_g63567 (.A(u0_n_31827),
    .B(u0_n_31823),
    .Y(u0_n_31569));
 NAND2xp33_ASAP7_75t_R u0_g63568 (.A(u0_n_31840),
    .B(u0_n_31837),
    .Y(u0_n_31570));
 XOR2xp5_ASAP7_75t_R u0_g63569 (.A(w2[26]),
    .B(w1[26]),
    .Y(u0_n_31572));
 NOR2xp33_ASAP7_75t_R u0_g63570 (.A(n_8942),
    .B(u0_n_31931),
    .Y(u0_n_31573));
 XNOR2xp5_ASAP7_75t_R u0_g63571 (.A(w2[10]),
    .B(u0_n_32683),
    .Y(u0_n_31712));
 XNOR2xp5_ASAP7_75t_R u0_g63572 (.A(w2[29]),
    .B(w3[29]),
    .Y(u0_n_31574));
 XOR2xp5_ASAP7_75t_R u0_g63573 (.A(w2[26]),
    .B(w3[26]),
    .Y(u0_n_31714));
 XNOR2xp5_ASAP7_75t_R u0_g63574 (.A(w2[15]),
    .B(u0_n_32714),
    .Y(u0_n_31715));
 XNOR2xp5_ASAP7_75t_R u0_g63575 (.A(w2[31]),
    .B(u0_n_32717),
    .Y(u0_n_31717));
 XOR2xp5_ASAP7_75t_R u0_g63576 (.A(w1[17]),
    .B(w0[17]),
    .Y(u0_n_31718));
 XNOR2xp5_ASAP7_75t_R u0_g63577 (.A(w2[2]),
    .B(u0_n_32695),
    .Y(u0_n_31720));
 XNOR2xp5_ASAP7_75t_R u0_g63578 (.A(w2[18]),
    .B(w3[18]),
    .Y(u0_n_31721));
 XNOR2xp5_ASAP7_75t_R u0_g63579 (.A(w2[24]),
    .B(w3[24]),
    .Y(u0_n_31722));
 XNOR2xp5_ASAP7_75t_R u0_g63580 (.A(w2[27]),
    .B(\u0_w[3] [27]),
    .Y(u0_n_31723));
 XNOR2xp5_ASAP7_75t_R u0_g63581 (.A(w2[4]),
    .B(n_8629),
    .Y(u0_n_31724));
 NAND2xp33_ASAP7_75t_L u0_g63582 (.A(u0_n_31983),
    .B(u0_n_31802),
    .Y(u0_n_31575));
 XNOR2xp5_ASAP7_75t_R u0_g63583 (.A(w2[20]),
    .B(u0_n_33138),
    .Y(u0_n_31726));
 NAND2xp33_ASAP7_75t_R u0_g63584 (.A(u0_n_31805),
    .B(u0_n_31976),
    .Y(u0_n_31576));
 AOI22xp33_ASAP7_75t_R u0_g63585 (.A1(n_8946),
    .A2(w2[28]),
    .B1(n_8942),
    .B2(u0_n_32571),
    .Y(u0_n_31727));
 XOR2xp5_ASAP7_75t_R u0_g63586 (.A(w0[14]),
    .B(w3[14]),
    .Y(u0_n_31729));
 NOR2xp33_ASAP7_75t_L u0_g63587 (.A(u0_n_32290),
    .B(u0_n_31791),
    .Y(u0_n_31578));
 NAND2xp33_ASAP7_75t_R u0_g63588 (.A(u0_n_31823),
    .B(u0_n_31791),
    .Y(u0_n_31580));
 XNOR2xp5_ASAP7_75t_R u0_g63589 (.A(w0[25]),
    .B(w1[25]),
    .Y(u0_n_31730));
 NAND2xp5_ASAP7_75t_L u0_g63590 (.A(u0_n_31794),
    .B(u0_n_32353),
    .Y(u0_n_31581));
 NAND2xp33_ASAP7_75t_R u0_g63591 (.A(u0_n_31826),
    .B(u0_n_31793),
    .Y(u0_n_31582));
 NAND2xp33_ASAP7_75t_R u0_g63592 (.A(u0_n_31815),
    .B(u0_n_31977),
    .Y(u0_n_31583));
 NOR2xp33_ASAP7_75t_L u0_g63593 (.A(u0_n_32385),
    .B(u0_n_31804),
    .Y(u0_n_31584));
 NAND2xp5_ASAP7_75t_R u0_g63594 (.A(u0_n_31840),
    .B(u0_n_31795),
    .Y(u0_n_31586));
 NOR2xp33_ASAP7_75t_L u0_g63595 (.A(u0_n_31810),
    .B(u0_n_32141),
    .Y(u0_n_31587));
 NOR2xp33_ASAP7_75t_R u0_g63596 (.A(u0_n_31808),
    .B(u0_n_32254),
    .Y(u0_n_31588));
 XOR2xp5_ASAP7_75t_R u0_g63597 (.A(w2[30]),
    .B(u0_n_33033),
    .Y(u0_n_31733));
 NAND2xp5_ASAP7_75t_R u0_g63598 (.A(u0_n_31819),
    .B(u0_n_31799),
    .Y(u0_n_31590));
 XNOR2xp5_ASAP7_75t_R u0_g63599 (.A(w2[3]),
    .B(w1[3]),
    .Y(u0_n_31734));
 XOR2xp5_ASAP7_75t_R u0_g63600 (.A(w2[23]),
    .B(w1[23]),
    .Y(u0_n_31736));
 XOR2xp5_ASAP7_75t_R u0_g63601 (.A(w2[5]),
    .B(w1[5]),
    .Y(u0_n_31738));
 XNOR2xp5_ASAP7_75t_R u0_g63602 (.A(w1[15]),
    .B(w2[15]),
    .Y(u0_n_31740));
 NOR2xp33_ASAP7_75t_R u0_g63603 (.A(u0_n_31814),
    .B(u0_n_32410),
    .Y(u0_n_31591));
 NAND2xp33_ASAP7_75t_R u0_g63604 (.A(u0_n_31841),
    .B(u0_n_31921),
    .Y(u0_n_31592));
 NOR2xp33_ASAP7_75t_R u0_g63605 (.A(u0_n_32254),
    .B(u0_n_31811),
    .Y(u0_n_31594));
 NAND2xp33_ASAP7_75t_R u0_g63606 (.A(u0_n_31962),
    .B(u0_n_32208),
    .Y(u0_n_31596));
 NAND2xp5_ASAP7_75t_L u0_g63607 (.A(u0_n_31959),
    .B(u0_n_31827),
    .Y(u0_n_31598));
 NAND2xp5_ASAP7_75t_R u0_g63608 (.A(u0_n_31818),
    .B(u0_n_31970),
    .Y(u0_n_31599));
 NAND2xp33_ASAP7_75t_R u0_g63609 (.A(u0_n_31934),
    .B(u0_n_31819),
    .Y(u0_n_31600));
 NOR2xp33_ASAP7_75t_SL u0_g63610 (.A(u0_n_31838),
    .B(u0_n_31964),
    .Y(u0_n_31602));
 NAND2xp33_ASAP7_75t_L u0_g63611 (.A(u0_n_31938),
    .B(u0_n_31818),
    .Y(u0_n_31605));
 NAND2xp33_ASAP7_75t_R u0_g63612 (.A(u0_n_31923),
    .B(u0_n_31823),
    .Y(u0_n_31606));
 NOR2x1_ASAP7_75t_SL u0_g63613 (.A(u0_n_31824),
    .B(u0_n_31971),
    .Y(u0_n_31607));
 NOR2xp33_ASAP7_75t_SL u0_g63614 (.A(u0_n_31822),
    .B(u0_n_31962),
    .Y(u0_n_31609));
 NOR2xp33_ASAP7_75t_SL u0_g63615 (.A(u0_n_31951),
    .B(u0_n_31825),
    .Y(u0_n_31610));
 NOR2xp33_ASAP7_75t_R u0_g63616 (.A(u0_n_31825),
    .B(u0_n_31928),
    .Y(u0_n_31612));
 NOR2xp33_ASAP7_75t_L u0_g63617 (.A(u0_n_31839),
    .B(u0_n_31920),
    .Y(u0_n_31614));
 NAND2xp5_ASAP7_75t_R u0_g63618 (.A(u0_n_31945),
    .B(u0_n_31837),
    .Y(u0_n_31616));
 NAND2xp5_ASAP7_75t_R u0_g63619 (.A(u0_n_31830),
    .B(u0_n_31943),
    .Y(u0_n_31618));
 NAND2xp5_ASAP7_75t_L u0_g63620 (.A(u0_n_31965),
    .B(u0_n_31821),
    .Y(u0_n_31620));
 NAND2xp5_ASAP7_75t_L u0_g63621 (.A(u0_n_31835),
    .B(u0_n_32273),
    .Y(u0_n_31621));
 NAND2xp33_ASAP7_75t_R u0_g63622 (.A(u0_n_31818),
    .B(u0_n_31813),
    .Y(u0_n_31623));
 NOR2xp33_ASAP7_75t_SL u0_g63623 (.A(u0_n_32344),
    .B(u0_n_31818),
    .Y(u0_n_31624));
 NOR2xp33_ASAP7_75t_L u0_g63624 (.A(u0_n_31810),
    .B(u0_n_31838),
    .Y(u0_n_31625));
 NOR2xp33_ASAP7_75t_SL u0_g63625 (.A(u0_n_31808),
    .B(u0_n_31822),
    .Y(u0_n_31627));
 NAND2xp5_ASAP7_75t_L u0_g63626 (.A(u0_n_31827),
    .B(u0_n_31803),
    .Y(u0_n_31629));
 NOR2xp33_ASAP7_75t_SL u0_g63627 (.A(u0_n_31825),
    .B(u0_n_31969),
    .Y(u0_n_31631));
 NAND2xp5_ASAP7_75t_R u0_g63628 (.A(u0_n_32012),
    .B(u0_n_31812),
    .Y(u0_n_31632));
 NAND2xp33_ASAP7_75t_R u0_g63629 (.A(u0_n_31815),
    .B(u0_n_31841),
    .Y(u0_n_31633));
 NAND2xp33_ASAP7_75t_L u0_g63630 (.A(u0_n_32308),
    .B(u0_n_31805),
    .Y(u0_n_31635));
 NAND2xp5_ASAP7_75t_R u0_g63631 (.A(u0_n_31802),
    .B(u0_n_32175),
    .Y(u0_n_31637));
 NOR2xp33_ASAP7_75t_R u0_g63632 (.A(u0_n_32761),
    .B(u0_n_31961),
    .Y(u0_n_31638));
 NOR2xp33_ASAP7_75t_L u0_g63633 (.A(u0_n_31815),
    .B(u0_n_31905),
    .Y(u0_n_31639));
 XNOR2xp5_ASAP7_75t_R u0_g63634 (.A(w1[14]),
    .B(w2[14]),
    .Y(u0_n_31642));
 NAND2xp5_ASAP7_75t_R u0_g63635 (.A(u0_n_31806),
    .B(u0_n_32273),
    .Y(u0_n_31643));
 NAND2xp5_ASAP7_75t_L u0_g63636 (.A(u0_n_31840),
    .B(u0_n_31963),
    .Y(u0_n_31644));
 NAND2xp5_ASAP7_75t_R u0_g63637 (.A(u0_n_32339),
    .B(u0_n_31801),
    .Y(u0_n_31646));
 NOR2xp67_ASAP7_75t_R u0_g63638 (.A(u0_n_31839),
    .B(u0_n_31936),
    .Y(u0_n_31648));
 NAND2xp5_ASAP7_75t_SL u0_g63639 (.A(u0_n_31819),
    .B(u0_n_31953),
    .Y(u0_n_31650));
 NAND2xp5_ASAP7_75t_SL u0_g63640 (.A(n_8946),
    .B(u0_n_31931),
    .Y(u0_n_31651));
 NOR2x1_ASAP7_75t_R u0_g63642 (.A(n_8964),
    .B(u0_n_31930),
    .Y(u0_n_31654));
 NAND2xp5_ASAP7_75t_L u0_g63643 (.A(u0_n_32208),
    .B(u0_n_31811),
    .Y(u0_n_31657));
 NAND2xp5_ASAP7_75t_SL u0_g63644 (.A(n_8964),
    .B(u0_n_31943),
    .Y(u0_n_31660));
 NOR2xp33_ASAP7_75t_SL u0_g63645 (.A(u0_n_32761),
    .B(u0_n_31918),
    .Y(u0_n_31661));
 NAND2x1_ASAP7_75t_SL u0_g63647 (.A(u0_n_31927),
    .B(\u0_w[3] [12]),
    .Y(u0_n_31665));
 NAND2xp5_ASAP7_75t_SL u0_g63648 (.A(u0_n_31961),
    .B(u0_n_32761),
    .Y(u0_n_31666));
 AND2x2_ASAP7_75t_SL u0_g63649 (.A(u0_n_32759),
    .B(u0_n_31938),
    .Y(u0_n_31668));
 NOR2xp67_ASAP7_75t_R u0_g63650 (.A(u0_n_31824),
    .B(n_8963),
    .Y(u0_n_31670));
 AND2x2_ASAP7_75t_SL u0_g63651 (.A(n_8623),
    .B(u0_n_31945),
    .Y(u0_n_31672));
 NOR2xp33_ASAP7_75t_SL u0_g63652 (.A(w3[12]),
    .B(u0_n_31825),
    .Y(u0_n_31674));
 NOR2xp67_ASAP7_75t_R u0_g63653 (.A(w3[4]),
    .B(u0_n_31839),
    .Y(u0_n_31676));
 NAND2xp5_ASAP7_75t_L u0_g63654 (.A(u0_n_32761),
    .B(u0_n_31819),
    .Y(u0_n_31678));
 AND2x2_ASAP7_75t_SL u0_g63655 (.A(w3[28]),
    .B(u0_n_31824),
    .Y(u0_n_31680));
 AND2x2_ASAP7_75t_L u0_g63656 (.A(n_8963),
    .B(u0_n_31943),
    .Y(u0_n_31682));
 NOR2xp67_ASAP7_75t_L u0_g63657 (.A(u0_n_32761),
    .B(u0_n_31819),
    .Y(u0_n_31684));
 AND2x2_ASAP7_75t_SL u0_g63658 (.A(\u0_w[3] [12]),
    .B(u0_n_31825),
    .Y(u0_n_31686));
 AND2x2_ASAP7_75t_L u0_g63659 (.A(w3[4]),
    .B(u0_n_31839),
    .Y(u0_n_31688));
 INVxp33_ASAP7_75t_R u0_g63660 (.A(u0_n_31748),
    .Y(u0_n_31747));
 INVxp67_ASAP7_75t_L u0_g63661 (.A(n_11521),
    .Y(u0_n_31749));
 INVxp33_ASAP7_75t_R u0_g63662 (.A(u0_n_31754),
    .Y(u0_n_31753));
 INVxp67_ASAP7_75t_R u0_g63663 (.A(u0_n_31755),
    .Y(u0_n_31756));
 INVxp33_ASAP7_75t_R u0_g63664 (.A(u0_n_31762),
    .Y(u0_n_31763));
 INVxp33_ASAP7_75t_R u0_g63665 (.A(u0_n_31764),
    .Y(u0_n_31765));
 INVxp33_ASAP7_75t_R u0_g63666 (.A(u0_n_31766),
    .Y(u0_n_31767));
 INVxp67_ASAP7_75t_R u0_g63667 (.A(u0_n_31770),
    .Y(u0_n_31771));
 INVx1_ASAP7_75t_L u0_g63668 (.A(u0_n_31772),
    .Y(u0_n_31773));
 INVx2_ASAP7_75t_SL u0_g63669 (.A(u0_n_31775),
    .Y(u0_n_31776));
 INVxp33_ASAP7_75t_R u0_g63670 (.A(u0_n_31777),
    .Y(u0_n_31778));
 INVxp33_ASAP7_75t_R u0_g63671 (.A(u0_n_31779),
    .Y(u0_n_31780));
 INVxp67_ASAP7_75t_SL u0_g63672 (.A(u0_n_31781),
    .Y(u0_n_31782));
 INVxp33_ASAP7_75t_R u0_g63673 (.A(u0_n_31783),
    .Y(u0_n_31784));
 INVxp33_ASAP7_75t_R u0_g63674 (.A(u0_n_31785),
    .Y(u0_n_31786));
 INVxp67_ASAP7_75t_R u0_g63675 (.A(u0_n_31787),
    .Y(u0_n_31788));
 INVxp67_ASAP7_75t_R u0_g63676 (.A(u0_n_31789),
    .Y(u0_n_31790));
 INVxp33_ASAP7_75t_R u0_g63677 (.A(u0_n_31791),
    .Y(u0_n_31792));
 INVxp67_ASAP7_75t_R u0_g63678 (.A(u0_n_31793),
    .Y(u0_n_31794));
 INVxp67_ASAP7_75t_R u0_g63679 (.A(u0_n_31795),
    .Y(u0_n_31796));
 INVxp67_ASAP7_75t_R u0_g63680 (.A(u0_n_31797),
    .Y(u0_n_31798));
 INVx1_ASAP7_75t_L u0_g63681 (.A(u0_n_31799),
    .Y(u0_n_31800));
 INVxp33_ASAP7_75t_R u0_g63682 (.A(u0_n_31801),
    .Y(u0_n_31802));
 INVxp67_ASAP7_75t_R u0_g63683 (.A(u0_n_31803),
    .Y(u0_n_31804));
 INVxp67_ASAP7_75t_L u0_g63684 (.A(u0_n_31805),
    .Y(u0_n_31806));
 INVx1_ASAP7_75t_SL u0_g63685 (.A(u0_n_31807),
    .Y(u0_n_31808));
 INVx1_ASAP7_75t_L u0_g63686 (.A(u0_n_31809),
    .Y(u0_n_31810));
 INVx1_ASAP7_75t_L u0_g63687 (.A(u0_n_31811),
    .Y(u0_n_31812));
 INVx1_ASAP7_75t_SL u0_g63688 (.A(u0_n_31813),
    .Y(u0_n_31814));
 INVx1_ASAP7_75t_R u0_g63689 (.A(u0_n_31815),
    .Y(u0_n_31816));
 INVx2_ASAP7_75t_SL u0_g63690 (.A(u0_n_31817),
    .Y(u0_n_31818));
 INVx1_ASAP7_75t_R u0_g63691 (.A(u0_n_31819),
    .Y(u0_n_31820));
 INVx2_ASAP7_75t_SL u0_g63692 (.A(u0_n_31821),
    .Y(u0_n_31822));
 INVx2_ASAP7_75t_SL u0_g63693 (.A(u0_n_31823),
    .Y(u0_n_31824));
 INVx2_ASAP7_75t_SL u0_g63694 (.A(u0_n_31825),
    .Y(u0_n_31826));
 INVx2_ASAP7_75t_L u0_g63698 (.A(u0_n_31835),
    .Y(u0_n_31830));
 INVxp67_ASAP7_75t_SL u0_g63699 (.A(u0_n_31827),
    .Y(u0_n_31835));
 INVx2_ASAP7_75t_R u0_g63700 (.A(u0_n_31837),
    .Y(u0_n_31838));
 INVx2_ASAP7_75t_SL u0_g63701 (.A(u0_n_31839),
    .Y(u0_n_31840));
 INVx3_ASAP7_75t_SL u0_g63702 (.A(u0_n_31846),
    .Y(u0_n_31841));
 INVx3_ASAP7_75t_L u0_g63710 (.A(u0_n_31841),
    .Y(u0_n_31842));
 INVx2_ASAP7_75t_L u0_g63715 (.A(u0_n_31842),
    .Y(u0_n_31850));
 INVx2_ASAP7_75t_L u0_g63737 (.A(u0_n_31875),
    .Y(u0_n_31874));
 INVx1_ASAP7_75t_SL u0_g63741 (.A(u0_n_31874),
    .Y(u0_n_31886));
 BUFx3_ASAP7_75t_SL u0_g63745 (.A(u0_n_31905),
    .Y(u0_n_31875));
 INVx1_ASAP7_75t_L u0_g63751 (.A(u0_n_31895),
    .Y(u0_n_31900));
 INVx2_ASAP7_75t_R u0_g63752 (.A(u0_n_31875),
    .Y(u0_n_31895));
 NAND2xp33_ASAP7_75t_R u0_g63755 (.A(u0_n_32839),
    .B(u0_n_32673),
    .Y(u0_n_31906));
 NAND2xp33_ASAP7_75t_R u0_g63756 (.A(u0_n_32737),
    .B(n_8625),
    .Y(u0_n_31748));
 NOR2xp33_ASAP7_75t_L u0_g63758 (.A(w3[26]),
    .B(w3[29]),
    .Y(u0_n_31751));
 NAND2xp33_ASAP7_75t_R u0_g63759 (.A(u0_n_33001),
    .B(n_11371),
    .Y(u0_n_31752));
 NAND2xp5_ASAP7_75t_L u0_g63760 (.A(n_8656),
    .B(u0_n_33138),
    .Y(u0_n_31754));
 NAND2xp5_ASAP7_75t_R u0_g63761 (.A(u0_n_32695),
    .B(u0_n_32691),
    .Y(u0_n_31755));
 NOR2xp33_ASAP7_75t_L u0_g63762 (.A(n_11401),
    .B(w3[13]),
    .Y(u0_n_31757));
 NAND2xp33_ASAP7_75t_R u0_g63763 (.A(u0_n_32763),
    .B(w3[2]),
    .Y(u0_n_31758));
 NOR2xp33_ASAP7_75t_R u0_g63764 (.A(w3[16]),
    .B(w3[21]),
    .Y(u0_n_31759));
 NOR2xp33_ASAP7_75t_L u0_g63765 (.A(w3[21]),
    .B(n_11371),
    .Y(u0_n_31760));
 NOR2xp33_ASAP7_75t_R u0_g63766 (.A(n_11482),
    .B(n_11507),
    .Y(u0_n_31761));
 NAND2xp33_ASAP7_75t_R u0_g63767 (.A(w3[14]),
    .B(w3[8]),
    .Y(u0_n_31762));
 NOR2xp33_ASAP7_75t_R u0_g63768 (.A(w3[10]),
    .B(w3[13]),
    .Y(u0_n_31764));
 NAND2xp5_ASAP7_75t_R u0_g63769 (.A(u0_n_32763),
    .B(w3[0]),
    .Y(u0_n_31766));
 NAND2xp5_ASAP7_75t_L u0_g63770 (.A(u0_n_32743),
    .B(u0_n_32689),
    .Y(u0_n_31768));
 NAND2xp5_ASAP7_75t_R u0_g63771 (.A(w3[30]),
    .B(w3[24]),
    .Y(u0_n_31769));
 NOR2xp67_ASAP7_75t_L u0_g63772 (.A(w3[18]),
    .B(w3[16]),
    .Y(u0_n_31770));
 NOR2x1p5_ASAP7_75t_SL u0_g63773 (.A(w3[7]),
    .B(w3[1]),
    .Y(u0_n_31772));
 AND2x2_ASAP7_75t_R u0_g63774 (.A(u0_n_32687),
    .B(u0_n_32743),
    .Y(u0_n_31774));
 OR2x2_ASAP7_75t_SL u0_g63775 (.A(w3[15]),
    .B(w3[9]),
    .Y(u0_n_31775));
 NOR2xp33_ASAP7_75t_L u0_g63776 (.A(w3[10]),
    .B(w3[8]),
    .Y(u0_n_31777));
 NOR2xp33_ASAP7_75t_L u0_g63777 (.A(w3[2]),
    .B(w3[0]),
    .Y(u0_n_31779));
 OR2x2_ASAP7_75t_SL u0_g63778 (.A(w3[31]),
    .B(w3[25]),
    .Y(u0_n_31781));
 NAND2xp5_ASAP7_75t_L u0_g63779 (.A(w3[8]),
    .B(w3[10]),
    .Y(u0_n_31783));
 NAND2x1p5_ASAP7_75t_SL u0_g63780 (.A(n_8833),
    .B(u0_n_32735),
    .Y(u0_n_31785));
 NAND2xp5_ASAP7_75t_L u0_g63781 (.A(\u0_w[3] [16]),
    .B(w3[18]),
    .Y(u0_n_31787));
 OR2x2_ASAP7_75t_SL u0_g63782 (.A(u0_n_32747),
    .B(u0_n_32695),
    .Y(u0_n_31789));
 NAND2xp5_ASAP7_75t_SL u0_g63783 (.A(n_8946),
    .B(u0_n_32698),
    .Y(u0_n_31791));
 NAND2xp5_ASAP7_75t_L u0_g63784 (.A(n_8851),
    .B(u0_n_32759),
    .Y(u0_n_31793));
 NAND2xp5_ASAP7_75t_L u0_g63785 (.A(n_8623),
    .B(n_8742),
    .Y(u0_n_31795));
 OR2x2_ASAP7_75t_L u0_g63786 (.A(u0_n_32743),
    .B(u0_n_32687),
    .Y(u0_n_31797));
 NAND2xp5_ASAP7_75t_SL u0_g63787 (.A(u0_n_33138),
    .B(u0_n_32735),
    .Y(u0_n_31799));
 AND2x2_ASAP7_75t_SL u0_g63788 (.A(w3[9]),
    .B(\u0_w[3] [12]),
    .Y(u0_n_31801));
 NAND2xp5_ASAP7_75t_SL u0_g63789 (.A(u0_n_32716),
    .B(n_8946),
    .Y(u0_n_31803));
 OR2x2_ASAP7_75t_SL u0_g63790 (.A(u0_n_32698),
    .B(n_8946),
    .Y(u0_n_31805));
 NAND2xp5_ASAP7_75t_SL u0_g63791 (.A(u0_n_32761),
    .B(n_8833),
    .Y(u0_n_31807));
 OR2x2_ASAP7_75t_SL u0_g63792 (.A(w3[7]),
    .B(w3[4]),
    .Y(u0_n_31809));
 AND2x2_ASAP7_75t_SL u0_g63793 (.A(w3[17]),
    .B(w3[20]),
    .Y(u0_n_31811));
 OR2x2_ASAP7_75t_SL u0_g63794 (.A(w3[15]),
    .B(\u0_w[3] [12]),
    .Y(u0_n_31813));
 OR2x2_ASAP7_75t_SL u0_g63795 (.A(n_8742),
    .B(n_8623),
    .Y(u0_n_31815));
 AND2x4_ASAP7_75t_SL u0_g63796 (.A(w3[15]),
    .B(\u0_w[3] [12]),
    .Y(u0_n_31817));
 NAND2x1p5_ASAP7_75t_SL u0_g63797 (.A(w3[23]),
    .B(w3[17]),
    .Y(u0_n_31819));
 OR2x2_ASAP7_75t_SL u0_g63798 (.A(n_8833),
    .B(u0_n_32761),
    .Y(u0_n_31821));
 OR2x6_ASAP7_75t_SL u0_g63799 (.A(u0_n_32698),
    .B(u0_n_32715),
    .Y(u0_n_31823));
 AND2x4_ASAP7_75t_SL u0_g63800 (.A(w3[9]),
    .B(w3[15]),
    .Y(u0_n_31825));
 NAND2xp5_ASAP7_75t_SL u0_g63801 (.A(w3[31]),
    .B(w3[28]),
    .Y(u0_n_31827));
 NAND2x1p5_ASAP7_75t_SL u0_g63802 (.A(w3[4]),
    .B(w3[7]),
    .Y(u0_n_31837));
 AND2x4_ASAP7_75t_SL u0_g63803 (.A(w3[1]),
    .B(w3[7]),
    .Y(u0_n_31839));
 NAND2x1p5_ASAP7_75t_SL u0_g63804 (.A(u0_n_32737),
    .B(u0_n_32766),
    .Y(u0_n_31846));
 NAND2xp5_ASAP7_75t_L u0_g63805 (.A(w3[6]),
    .B(w3[3]),
    .Y(u0_n_31905));
 INVxp33_ASAP7_75t_R u0_g63806 (.A(u0_n_31911),
    .Y(u0_n_31910));
 INVxp33_ASAP7_75t_R u0_g63807 (.A(u0_n_31913),
    .Y(u0_n_31912));
 INVxp33_ASAP7_75t_R u0_g63808 (.A(u0_n_31915),
    .Y(u0_n_31914));
 INVxp33_ASAP7_75t_R u0_g63809 (.A(u0_n_31918),
    .Y(u0_n_31919));
 INVxp67_ASAP7_75t_R u0_g63810 (.A(u0_n_31920),
    .Y(u0_n_31921));
 INVx1_ASAP7_75t_L u0_g63811 (.A(u0_n_31922),
    .Y(u0_n_31923));
 INVx1_ASAP7_75t_L u0_g63813 (.A(u0_n_31926),
    .Y(u0_n_31927));
 INVxp67_ASAP7_75t_R u0_g63814 (.A(u0_n_31928),
    .Y(u0_n_31929));
 INVxp67_ASAP7_75t_SL u0_g63815 (.A(u0_n_31930),
    .Y(u0_n_31931));
 INVxp67_ASAP7_75t_R u0_g63816 (.A(u0_n_31933),
    .Y(u0_n_31932));
 INVxp67_ASAP7_75t_R u0_g63817 (.A(u0_n_31934),
    .Y(u0_n_31935));
 INVx1_ASAP7_75t_SL u0_g63818 (.A(u0_n_31936),
    .Y(u0_n_31937));
 INVxp67_ASAP7_75t_R u0_g63819 (.A(u0_n_31939),
    .Y(u0_n_31940));
 INVxp33_ASAP7_75t_R u0_g63820 (.A(u0_n_31941),
    .Y(u0_n_31942));
 INVxp67_ASAP7_75t_R u0_g63821 (.A(u0_n_31943),
    .Y(u0_n_31944));
 INVxp33_ASAP7_75t_R u0_g63823 (.A(u0_n_31945),
    .Y(u0_n_31946));
 INVxp67_ASAP7_75t_R u0_g63825 (.A(u0_n_31949),
    .Y(u0_n_31950));
 INVxp33_ASAP7_75t_R u0_g63826 (.A(u0_n_31951),
    .Y(u0_n_31952));
 INVxp67_ASAP7_75t_SL u0_g63827 (.A(u0_n_31953),
    .Y(u0_n_31954));
 INVxp33_ASAP7_75t_R u0_g63828 (.A(u0_n_31955),
    .Y(u0_n_31956));
 INVxp33_ASAP7_75t_R u0_g63829 (.A(u0_n_31957),
    .Y(u0_n_31958));
 INVxp33_ASAP7_75t_R u0_g63830 (.A(u0_n_31959),
    .Y(u0_n_31960));
 INVx1_ASAP7_75t_SL u0_g63831 (.A(u0_n_31961),
    .Y(u0_n_31962));
 INVx1_ASAP7_75t_SL u0_g63832 (.A(u0_n_31963),
    .Y(u0_n_31964));
 INVx1_ASAP7_75t_L u0_g63833 (.A(u0_n_31965),
    .Y(u0_n_31966));
 INVxp67_ASAP7_75t_R u0_g63834 (.A(u0_n_31967),
    .Y(u0_n_31968));
 INVxp67_ASAP7_75t_R u0_g63835 (.A(u0_n_31969),
    .Y(u0_n_31970));
 INVx1_ASAP7_75t_SL u0_g63836 (.A(u0_n_31971),
    .Y(u0_n_31972));
 INVxp67_ASAP7_75t_R u0_g63837 (.A(u0_n_31973),
    .Y(u0_n_31974));
 INVxp67_ASAP7_75t_L u0_g63838 (.A(u0_n_31975),
    .Y(u0_n_31976));
 BUFx2_ASAP7_75t_L u0_g63842 (.A(u0_n_31981),
    .Y(u0_n_31977));
 INVx1_ASAP7_75t_L u0_g63843 (.A(u0_n_31982),
    .Y(u0_n_31983));
 INVxp67_ASAP7_75t_R u0_g63844 (.A(u0_n_31984),
    .Y(u0_n_31985));
 INVx2_ASAP7_75t_SL u0_g63852 (.A(u0_n_31988),
    .Y(u0_n_31986));
 INVx3_ASAP7_75t_SL u0_g63863 (.A(u0_n_31998),
    .Y(u0_n_31988));
 INVxp67_ASAP7_75t_L u0_g63875 (.A(u0_n_32021),
    .Y(u0_n_32023));
 BUFx2_ASAP7_75t_SL u0_g63877 (.A(u0_n_32012),
    .Y(u0_n_32021));
 INVx2_ASAP7_75t_SL u0_g63883 (.A(u0_n_32012),
    .Y(u0_n_32017));
 INVx2_ASAP7_75t_SL u0_g63884 (.A(u0_n_32011),
    .Y(u0_n_32012));
 INVx1_ASAP7_75t_L u0_g63898 (.A(u0_n_32053),
    .Y(u0_n_32052));
 BUFx2_ASAP7_75t_SL u0_g63900 (.A(u0_n_32042),
    .Y(u0_n_32053));
 INVxp67_ASAP7_75t_R u0_g63902 (.A(u0_n_32042),
    .Y(u0_n_32063));
 INVx3_ASAP7_75t_SL u0_g63907 (.A(u0_n_32040),
    .Y(u0_n_32042));
 INVx1_ASAP7_75t_L u0_g63912 (.A(u0_n_32075),
    .Y(u0_n_32073));
 INVx1_ASAP7_75t_SL u0_g63923 (.A(u0_n_32080),
    .Y(u0_n_32083));
 INVx1_ASAP7_75t_L u0_g63931 (.A(u0_n_32080),
    .Y(u0_n_32075));
 INVx1_ASAP7_75t_SL u0_g63936 (.A(u0_n_32083),
    .Y(u0_n_32084));
 INVx2_ASAP7_75t_L u0_g63946 (.A(u0_n_32113),
    .Y(u0_n_32108));
 BUFx2_ASAP7_75t_SL u0_g63952 (.A(u0_n_32113),
    .Y(u0_n_32122));
 INVx1_ASAP7_75t_L u0_g63956 (.A(u0_n_32108),
    .Y(u0_n_32109));
 INVx1_ASAP7_75t_L u0_g63959 (.A(u0_n_32122),
    .Y(u0_n_32121));
 INVx2_ASAP7_75t_L u0_g63967 (.A(u0_n_32142),
    .Y(u0_n_32141));
 INVx2_ASAP7_75t_L u0_g63968 (.A(u0_n_32160),
    .Y(u0_n_32142));
 INVx1_ASAP7_75t_SL u0_g63985 (.A(u0_n_32166),
    .Y(u0_n_32165));
 INVx1_ASAP7_75t_SL u0_g63986 (.A(u0_n_32160),
    .Y(u0_n_32166));
 INVx1_ASAP7_75t_L u0_g63995 (.A(u0_n_32184),
    .Y(u0_n_32185));
 BUFx2_ASAP7_75t_SL u0_g63999 (.A(u0_n_32175),
    .Y(u0_n_32184));
 INVx2_ASAP7_75t_SL u0_g64000 (.A(u0_n_32174),
    .Y(u0_n_32175));
 INVx2_ASAP7_75t_SL u0_g64005 (.A(u0_n_32174),
    .Y(u0_n_32193));
 INVx2_ASAP7_75t_L u0_g64011 (.A(u0_n_32193),
    .Y(u0_n_32194));
 INVx1_ASAP7_75t_L u0_g64031 (.A(u0_n_32221),
    .Y(u0_n_32226));
 INVx2_ASAP7_75t_SL u0_g64032 (.A(u0_n_32208),
    .Y(u0_n_32221));
 INVx2_ASAP7_75t_L u0_g64039 (.A(u0_n_32208),
    .Y(u0_n_32209));
 INVx1_ASAP7_75t_L u0_g64046 (.A(u0_n_32241),
    .Y(u0_n_32242));
 INVxp67_ASAP7_75t_R u0_g64049 (.A(u0_n_32248),
    .Y(u0_n_32249));
 BUFx2_ASAP7_75t_L u0_g64050 (.A(u0_n_32241),
    .Y(u0_n_32248));
 INVx2_ASAP7_75t_SL u0_g64052 (.A(u0_n_32254),
    .Y(u0_n_32241));
 INVx1_ASAP7_75t_R u0_g64060 (.A(u0_n_32254),
    .Y(u0_n_32260));
 INVx1_ASAP7_75t_L u0_g64073 (.A(u0_n_32273),
    .Y(u0_n_32272));
 INVx1_ASAP7_75t_SL u0_g64080 (.A(u0_n_32290),
    .Y(u0_n_32289));
 INVx2_ASAP7_75t_SL u0_g64088 (.A(u0_n_32273),
    .Y(u0_n_32290));
 INVx1_ASAP7_75t_R u0_g64095 (.A(u0_n_32306),
    .Y(u0_n_32308));
 INVxp67_ASAP7_75t_L u0_g64097 (.A(u0_n_32304),
    .Y(u0_n_32315));
 INVxp67_ASAP7_75t_SL u0_g64099 (.A(u0_n_32306),
    .Y(u0_n_32304));
 INVx1_ASAP7_75t_SL u0_g64102 (.A(u0_n_32321),
    .Y(u0_n_32320));
 BUFx2_ASAP7_75t_R u0_g64110 (.A(u0_n_32306),
    .Y(u0_n_32321));
 INVx2_ASAP7_75t_R u0_g64119 (.A(u0_n_32339),
    .Y(u0_n_32344));
 INVx2_ASAP7_75t_R u0_g64133 (.A(u0_n_32338),
    .Y(u0_n_32353));
 INVx2_ASAP7_75t_SL u0_g64134 (.A(u0_n_32339),
    .Y(u0_n_32338));
 INVx1_ASAP7_75t_SL u0_g64149 (.A(u0_n_32372),
    .Y(u0_n_32373));
 INVx1_ASAP7_75t_SL u0_g64153 (.A(u0_n_32386),
    .Y(u0_n_32387));
 INVx2_ASAP7_75t_R u0_g64155 (.A(u0_n_32385),
    .Y(u0_n_32386));
 BUFx3_ASAP7_75t_SL u0_g64164 (.A(u0_n_32372),
    .Y(u0_n_32385));
 INVx1_ASAP7_75t_L u0_g64182 (.A(u0_n_32416),
    .Y(u0_n_32425));
 INVx2_ASAP7_75t_L u0_g64183 (.A(u0_n_32410),
    .Y(u0_n_32416));
 INVx2_ASAP7_75t_SL u0_g64187 (.A(u0_n_32407),
    .Y(u0_n_32409));
 INVx3_ASAP7_75t_SL u0_g64189 (.A(u0_n_32410),
    .Y(u0_n_32407));
 NOR2xp33_ASAP7_75t_R u0_g64190 (.A(n_11371),
    .B(u0_n_32731),
    .Y(u0_n_31909));
 NOR2xp33_ASAP7_75t_R u0_g64191 (.A(w3[26]),
    .B(u0_n_32689),
    .Y(u0_n_31911));
 NAND2xp33_ASAP7_75t_R u0_g64192 (.A(n_11507),
    .B(u0_n_32695),
    .Y(u0_n_31913));
 NOR2xp33_ASAP7_75t_R u0_g64193 (.A(w3[10]),
    .B(u0_n_32685),
    .Y(u0_n_31915));
 NAND2xp5_ASAP7_75t_R u0_g64194 (.A(n_8831),
    .B(n_8656),
    .Y(u0_n_31916));
 NAND2xp33_ASAP7_75t_R u0_g64195 (.A(w3[22]),
    .B(\u0_w[3] [16]),
    .Y(u0_n_31917));
 AND2x2_ASAP7_75t_SL u0_g64196 (.A(w3[17]),
    .B(n_8833),
    .Y(u0_n_31918));
 NOR2xp33_ASAP7_75t_L u0_g64197 (.A(w3[1]),
    .B(n_8623),
    .Y(u0_n_31920));
 NOR2xp33_ASAP7_75t_SL u0_g64198 (.A(n_8946),
    .B(w3[25]),
    .Y(u0_n_31922));
 NOR2x1_ASAP7_75t_SL u0_g64199 (.A(w3[7]),
    .B(n_8742),
    .Y(u0_n_31924));
 NOR2x1_ASAP7_75t_SL u0_g64200 (.A(w3[15]),
    .B(n_8851),
    .Y(u0_n_31926));
 NOR2xp33_ASAP7_75t_R u0_g64201 (.A(w3[9]),
    .B(u0_n_32759),
    .Y(u0_n_31928));
 AND2x2_ASAP7_75t_SL u0_g64202 (.A(w3[25]),
    .B(u0_n_32716),
    .Y(u0_n_31930));
 NOR2xp33_ASAP7_75t_R u0_g64203 (.A(w3[10]),
    .B(u0_n_32745),
    .Y(u0_n_31933));
 NAND2xp5_ASAP7_75t_R u0_g64204 (.A(u0_n_32735),
    .B(w3[20]),
    .Y(u0_n_31934));
 AND2x2_ASAP7_75t_SL u0_g64205 (.A(w3[4]),
    .B(u0_n_32697),
    .Y(u0_n_31936));
 NAND2x1_ASAP7_75t_SL u0_g64206 (.A(n_8851),
    .B(w3[15]),
    .Y(u0_n_31938));
 NAND2xp5_ASAP7_75t_R u0_g64207 (.A(w3[24]),
    .B(u0_n_32687),
    .Y(u0_n_31939));
 NAND2xp5_ASAP7_75t_R u0_g64208 (.A(w3[0]),
    .B(u0_n_32695),
    .Y(u0_n_31941));
 NAND2xp5_ASAP7_75t_SL u0_g64209 (.A(u0_n_32706),
    .B(w3[31]),
    .Y(u0_n_31943));
 NAND2x1p5_ASAP7_75t_SL u0_g64210 (.A(w3[7]),
    .B(n_8742),
    .Y(u0_n_31945));
 NAND2xp5_ASAP7_75t_R u0_g64211 (.A(\u0_w[3] [16]),
    .B(u0_n_32741),
    .Y(u0_n_31949));
 AND2x2_ASAP7_75t_SL u0_g64212 (.A(\u0_w[3] [12]),
    .B(u0_n_32714),
    .Y(u0_n_31951));
 NAND2xp5_ASAP7_75t_SL u0_g64213 (.A(n_8833),
    .B(w3[20]),
    .Y(u0_n_31953));
 NOR2x1p5_ASAP7_75t_L u0_g64214 (.A(n_11401),
    .B(u0_n_32683),
    .Y(u0_n_31955));
 AND2x2_ASAP7_75t_SL u0_g64215 (.A(u0_n_32753),
    .B(w3[18]),
    .Y(u0_n_31957));
 NAND2x1_ASAP7_75t_L u0_g64216 (.A(n_8964),
    .B(u0_n_32704),
    .Y(u0_n_31959));
 NAND2x1_ASAP7_75t_SL u0_g64217 (.A(w3[23]),
    .B(u0_n_32735),
    .Y(u0_n_31961));
 NAND2xp5_ASAP7_75t_SL u0_g64218 (.A(w3[1]),
    .B(n_8623),
    .Y(u0_n_31963));
 NAND2xp5_ASAP7_75t_SL u0_g64219 (.A(w3[17]),
    .B(u0_n_33138),
    .Y(u0_n_31965));
 NOR2x1_ASAP7_75t_L u0_g64220 (.A(w3[0]),
    .B(u0_n_32695),
    .Y(u0_n_31967));
 NOR2x1_ASAP7_75t_SL u0_g64221 (.A(\u0_w[3] [12]),
    .B(n_8851),
    .Y(u0_n_31969));
 AND2x2_ASAP7_75t_SL u0_g64222 (.A(w3[28]),
    .B(u0_n_32715),
    .Y(u0_n_31971));
 NOR2x1_ASAP7_75t_L u0_g64223 (.A(w3[24]),
    .B(u0_n_32687),
    .Y(u0_n_31973));
 NOR2x1_ASAP7_75t_L u0_g64224 (.A(u0_n_32715),
    .B(w3[28]),
    .Y(u0_n_31975));
 NAND2xp5_ASAP7_75t_SL u0_g64225 (.A(w3[7]),
    .B(n_8623),
    .Y(u0_n_31981));
 AND2x2_ASAP7_75t_SL u0_g64226 (.A(w3[15]),
    .B(u0_n_32759),
    .Y(u0_n_31982));
 AND2x2_ASAP7_75t_SL u0_g64227 (.A(w3[23]),
    .B(u0_n_32761),
    .Y(u0_n_31984));
 NOR2x1p5_ASAP7_75t_SL u0_g64228 (.A(w3[19]),
    .B(u0_n_32795),
    .Y(u0_n_31998));
 NAND2xp5_ASAP7_75t_SL u0_g64229 (.A(n_8652),
    .B(u0_n_32795),
    .Y(u0_n_32011));
 NOR2x1p5_ASAP7_75t_SL u0_g64230 (.A(\u0_w[3] [27]),
    .B(u0_n_32793),
    .Y(u0_n_32040));
 NOR2x1p5_ASAP7_75t_SL u0_g64231 (.A(w3[3]),
    .B(u0_n_32766),
    .Y(u0_n_32080));
 AND2x2_ASAP7_75t_SL u0_g64232 (.A(w3[14]),
    .B(u0_n_32749),
    .Y(u0_n_32113));
 NAND2xp5_ASAP7_75t_SL u0_g64233 (.A(u0_n_32766),
    .B(w3[3]),
    .Y(u0_n_32160));
 NAND2x1p5_ASAP7_75t_L u0_g64234 (.A(u0_n_32749),
    .B(n_8801),
    .Y(u0_n_32174));
 AND2x6_ASAP7_75t_L u0_g64235 (.A(w3[22]),
    .B(w3[19]),
    .Y(u0_n_32208));
 OR2x4_ASAP7_75t_SL u0_g64236 (.A(w3[22]),
    .B(n_8652),
    .Y(u0_n_32254));
 AND2x6_ASAP7_75t_L u0_g64237 (.A(\u0_w[3] [30]),
    .B(\u0_w[3] [27]),
    .Y(u0_n_32273));
 OR2x2_ASAP7_75t_SL u0_g64238 (.A(\u0_w[3] [30]),
    .B(\u0_w[3] [27]),
    .Y(u0_n_32306));
 AND2x6_ASAP7_75t_L u0_g64239 (.A(w3[14]),
    .B(w3[11]),
    .Y(u0_n_32339));
 OR2x2_ASAP7_75t_SL u0_g64240 (.A(\u0_w[3] [30]),
    .B(u0_n_32751),
    .Y(u0_n_32372));
 OR2x2_ASAP7_75t_SL u0_g64241 (.A(w3[14]),
    .B(u0_n_32749),
    .Y(u0_n_32410));
 HB1xp67_ASAP7_75t_R u0_g64283 (.A(w2[21]),
    .Y(u0_n_32528));
 INVxp33_ASAP7_75t_R u0_g64305 (.A(w2[28]),
    .Y(u0_n_32571));
 INVxp33_ASAP7_75t_R u0_g64375 (.A(u0_r0_rcnt[0]),
    .Y(u0_n_32673));
 INVxp33_ASAP7_75t_R u0_g64376 (.A(w1[26]),
    .Y(u0_n_32675));
 INVx2_ASAP7_75t_L u0_g64382 (.A(w3[10]),
    .Y(u0_n_32683));
 INVx2_ASAP7_75t_L u0_g64383 (.A(w3[13]),
    .Y(u0_n_32685));
 INVx3_ASAP7_75t_SL u0_g64384 (.A(w3[26]),
    .Y(u0_n_32687));
 INVx1_ASAP7_75t_R u0_g64385 (.A(w3[29]),
    .Y(u0_n_32689));
 INVx1_ASAP7_75t_L u0_g64386 (.A(w3[5]),
    .Y(u0_n_32691));
 INVx3_ASAP7_75t_L u0_g64388 (.A(w3[2]),
    .Y(u0_n_32695));
 INVx1_ASAP7_75t_SL u0_g64389 (.A(w3[7]),
    .Y(u0_n_32697));
 INVx4_ASAP7_75t_SL u0_g64394 (.A(w3[25]),
    .Y(u0_n_32698));
 INVx1_ASAP7_75t_L u0_g64401 (.A(u0_n_32706),
    .Y(u0_n_32704));
 INVx2_ASAP7_75t_SL u0_g64402 (.A(w3[25]),
    .Y(u0_n_32706));
 INVx2_ASAP7_75t_SL u0_g64403 (.A(w3[15]),
    .Y(u0_n_32714));
 INVx1_ASAP7_75t_L u0_g64411 (.A(u0_n_32716),
    .Y(u0_n_32717));
 INVx2_ASAP7_75t_R u0_g64413 (.A(w3[31]),
    .Y(u0_n_32716));
 INVx4_ASAP7_75t_SL u0_g64414 (.A(w3[31]),
    .Y(u0_n_32715));
 INVx1_ASAP7_75t_SL u0_g64416 (.A(w3[21]),
    .Y(u0_n_32731));
 INVx6_ASAP7_75t_SL u0_g64418 (.A(w3[17]),
    .Y(u0_n_32735));
 INVx2_ASAP7_75t_L u0_g64419 (.A(w3[3]),
    .Y(u0_n_32737));
 INVx1_ASAP7_75t_L u0_g64421 (.A(w3[18]),
    .Y(u0_n_32741));
 INVx2_ASAP7_75t_L u0_g64422 (.A(w3[24]),
    .Y(u0_n_32743));
 INVxp67_ASAP7_75t_R u0_g64423 (.A(w3[8]),
    .Y(u0_n_32745));
 INVx1_ASAP7_75t_SL u0_g64424 (.A(w3[0]),
    .Y(u0_n_32747));
 INVx2_ASAP7_75t_SL u0_g64425 (.A(w3[11]),
    .Y(u0_n_32749));
 INVx2_ASAP7_75t_L u0_g64426 (.A(\u0_w[3] [27]),
    .Y(u0_n_32751));
 INVx2_ASAP7_75t_R u0_g64427 (.A(\u0_w[3] [16]),
    .Y(u0_n_32753));
 INVx2_ASAP7_75t_SL u0_g64430 (.A(\u0_w[3] [12]),
    .Y(u0_n_32759));
 INVx4_ASAP7_75t_SL u0_g64431 (.A(w3[20]),
    .Y(u0_n_32761));
 INVxp67_ASAP7_75t_L u0_g64446 (.A(u0_n_32774),
    .Y(u0_n_32773));
 HB1xp67_ASAP7_75t_SL u0_g64450 (.A(u0_n_32763),
    .Y(u0_n_32774));
 INVx2_ASAP7_75t_SL u0_g64451 (.A(u0_n_32766),
    .Y(u0_n_32763));
 INVx3_ASAP7_75t_SL u0_g64453 (.A(w3[6]),
    .Y(u0_n_32766));
 INVx3_ASAP7_75t_SL u0_g64456 (.A(\u0_w[3] [30]),
    .Y(u0_n_32793));
 INVx2_ASAP7_75t_L u0_g64457 (.A(\u0_w[3] [22]),
    .Y(u0_n_32795));
 INVxp33_ASAP7_75t_R u0_g64458 (.A(key[9]),
    .Y(u0_n_32796));
 INVxp33_ASAP7_75t_R u0_g64459 (.A(key[12]),
    .Y(u0_n_32797));
 INVxp33_ASAP7_75t_R u0_g64460 (.A(key[24]),
    .Y(u0_n_32798));
 INVxp33_ASAP7_75t_R u0_g64461 (.A(key[2]),
    .Y(u0_n_32799));
 INVxp33_ASAP7_75t_R u0_g64462 (.A(key[25]),
    .Y(u0_n_32800));
 INVxp33_ASAP7_75t_R u0_g64463 (.A(key[4]),
    .Y(u0_n_32801));
 INVxp33_ASAP7_75t_R u0_g64464 (.A(key[21]),
    .Y(u0_n_32802));
 INVxp33_ASAP7_75t_R u0_g64465 (.A(key[0]),
    .Y(u0_n_32803));
 INVxp33_ASAP7_75t_R u0_g64466 (.A(key[20]),
    .Y(u0_n_32804));
 INVxp33_ASAP7_75t_R u0_g64467 (.A(key[11]),
    .Y(u0_n_32805));
 INVxp33_ASAP7_75t_R u0_g64468 (.A(key[6]),
    .Y(u0_n_32806));
 INVxp33_ASAP7_75t_R u0_g64469 (.A(key[16]),
    .Y(u0_n_32807));
 INVxp33_ASAP7_75t_R u0_g64470 (.A(key[28]),
    .Y(u0_n_32808));
 INVxp33_ASAP7_75t_R u0_g64471 (.A(key[31]),
    .Y(u0_n_32809));
 INVxp33_ASAP7_75t_R u0_g64472 (.A(key[27]),
    .Y(u0_n_32810));
 INVxp33_ASAP7_75t_R u0_g64473 (.A(key[3]),
    .Y(u0_n_32811));
 INVxp33_ASAP7_75t_R u0_g64474 (.A(key[22]),
    .Y(u0_n_32812));
 INVxp33_ASAP7_75t_R u0_g64475 (.A(key[19]),
    .Y(u0_n_32813));
 INVxp33_ASAP7_75t_R u0_g64476 (.A(key[18]),
    .Y(u0_n_32814));
 INVxp33_ASAP7_75t_R u0_g64477 (.A(key[8]),
    .Y(u0_n_32815));
 INVxp33_ASAP7_75t_R u0_g64478 (.A(key[23]),
    .Y(u0_n_32816));
 INVxp33_ASAP7_75t_R u0_g64479 (.A(key[17]),
    .Y(u0_n_32817));
 INVxp33_ASAP7_75t_R u0_g64480 (.A(key[30]),
    .Y(u0_n_32818));
 INVxp33_ASAP7_75t_R u0_g64481 (.A(key[15]),
    .Y(u0_n_32819));
 INVxp33_ASAP7_75t_R u0_g64482 (.A(key[1]),
    .Y(u0_n_32820));
 INVxp33_ASAP7_75t_R u0_g64483 (.A(key[14]),
    .Y(u0_n_32821));
 INVxp33_ASAP7_75t_R u0_g64484 (.A(key[7]),
    .Y(u0_n_32822));
 HB1xp67_ASAP7_75t_R u0_g64486 (.A(u0_n_32843),
    .Y(u0_n_32825));
 INVx2_ASAP7_75t_L u0_g64489 (.A(u0_n_32835),
    .Y(u0_n_32836));
 BUFx2_ASAP7_75t_R u0_g64495 (.A(u0_n_32834),
    .Y(u0_n_32845));
 INVxp67_ASAP7_75t_R u0_g64503 (.A(u0_n_32836),
    .Y(u0_n_32879));
 INVx1_ASAP7_75t_L u0_g64504 (.A(u0_n_32834),
    .Y(u0_n_32877));
 INVx1_ASAP7_75t_SL u0_g64508 (.A(u0_n_32843),
    .Y(u0_n_32839));
 INVx2_ASAP7_75t_R u0_g64511 (.A(u0_n_32843),
    .Y(u0_n_32924));
 BUFx2_ASAP7_75t_R u0_g64513 (.A(u0_n_32836),
    .Y(u0_n_32934));
 BUFx2_ASAP7_75t_R u0_g64514 (.A(u0_n_32834),
    .Y(u0_n_32942));
 INVx1_ASAP7_75t_R u0_g64515 (.A(u0_n_32836),
    .Y(u0_n_32875));
 XNOR2xp5_ASAP7_75t_SL u0_g64681 (.A(u0_n_29681),
    .B(u0_n_31642),
    .Y(u0_n_33150));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[24]  (.CLK(clk),
    .D(u0_n_31188),
    .QN(u0_rcon[24]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[25]  (.CLK(clk),
    .D(u0_n_30046),
    .QN(u0_rcon[25]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[26]  (.CLK(clk),
    .D(u0_n_29890),
    .QN(u0_rcon[26]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[27]  (.CLK(clk),
    .D(u0_n_29892),
    .QN(u0_rcon[27]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[28]  (.CLK(clk),
    .D(u0_n_29898),
    .QN(u0_rcon[28]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[29]  (.CLK(clk),
    .D(u0_n_29904),
    .QN(u0_rcon[29]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[30]  (.CLK(clk),
    .D(u0_n_30047),
    .QN(u0_rcon[30]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_out_reg[31]  (.CLK(clk),
    .D(u0_n_29986),
    .QN(u0_rcon[31]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_rcnt_reg[0]  (.CLK(clk),
    .D(u0_n_31906),
    .QN(u0_r0_rcnt[0]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_rcnt_reg[1]  (.CLK(clk),
    .D(u0_n_31200),
    .QN(u0_r0_rcnt[1]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_rcnt_reg[2]  (.CLK(clk),
    .D(u0_n_30785),
    .QN(u0_r0_rcnt[2]));
 DFFHQNx1_ASAP7_75t_R \u0_r0_rcnt_reg[3]  (.CLK(clk),
    .D(u0_n_30383),
    .QN(u0_r0_rcnt[3]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][0]  (.CLK(clk),
    .D(u0_n_29544),
    .QN(w0[0]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[0][10]  (.CLK(clk),
    .D(u0_n_29533),
    .QN(w0[10]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][11]  (.CLK(clk),
    .D(u0_n_29534),
    .QN(w0[11]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][12]  (.CLK(clk),
    .D(u0_n_29462),
    .QN(w0[12]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][13]  (.CLK(clk),
    .D(u0_n_29538),
    .QN(w0[13]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][14]  (.CLK(clk),
    .D(u0_n_29539),
    .QN(w0[14]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][15]  (.CLK(clk),
    .D(u0_n_29489),
    .QN(w0[15]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][16]  (.CLK(clk),
    .D(u0_n_29536),
    .QN(w0[16]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][17]  (.CLK(clk),
    .D(u0_n_29526),
    .QN(w0[17]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][18]  (.CLK(clk),
    .D(u0_n_29527),
    .QN(w0[18]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][19]  (.CLK(clk),
    .D(u0_n_29529),
    .QN(w0[19]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][1]  (.CLK(clk),
    .D(u0_n_29461),
    .QN(w0[1]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][20]  (.CLK(clk),
    .D(u0_n_29624),
    .QN(w0[20]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][21]  (.CLK(clk),
    .D(u0_n_29530),
    .QN(w0[21]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][22]  (.CLK(clk),
    .D(u0_n_29531),
    .QN(w0[22]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][23]  (.CLK(clk),
    .D(u0_n_29623),
    .QN(w0[23]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][24]  (.CLK(clk),
    .D(u0_n_29380),
    .QN(w0[24]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[0][25]  (.CLK(clk),
    .D(u0_n_29373),
    .QN(w0[25]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[0][26]  (.CLK(clk),
    .D(u0_n_29379),
    .QN(w0[26]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][27]  (.CLK(clk),
    .D(u0_n_29535),
    .QN(w0[27]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][28]  (.CLK(clk),
    .D(u0_n_29483),
    .QN(w0[28]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][29]  (.CLK(clk),
    .D(u0_n_29537),
    .QN(w0[29]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][2]  (.CLK(clk),
    .D(u0_n_29484),
    .QN(w0[2]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[0][30]  (.CLK(clk),
    .D(u0_n_29334),
    .QN(w0[30]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][31]  (.CLK(clk),
    .D(u0_n_29540),
    .QN(w0[31]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][3]  (.CLK(clk),
    .D(u0_n_29532),
    .QN(w0[3]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[0][4]  (.CLK(clk),
    .D(u0_n_29485),
    .QN(w0[4]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][5]  (.CLK(clk),
    .D(u0_n_29523),
    .QN(w0[5]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[0][6]  (.CLK(clk),
    .D(u0_n_29491),
    .QN(w0[6]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[0][7]  (.CLK(clk),
    .D(u0_n_29493),
    .QN(w0[7]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][8]  (.CLK(clk),
    .D(u0_n_29528),
    .QN(w0[8]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[0][9]  (.CLK(clk),
    .D(u0_n_29459),
    .QN(w0[9]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][0]  (.CLK(clk),
    .D(u0_n_29378),
    .QN(w1[0]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][10]  (.CLK(clk),
    .D(u0_n_29541),
    .QN(w1[10]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][11]  (.CLK(clk),
    .D(u0_n_29376),
    .QN(w1[11]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][12]  (.CLK(clk),
    .D(u0_n_29488),
    .QN(w1[12]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][13]  (.CLK(clk),
    .D(u0_n_29375),
    .QN(w1[13]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][14]  (.CLK(clk),
    .D(u0_n_29386),
    .QN(w1[14]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][15]  (.CLK(clk),
    .D(u0_n_29337),
    .QN(w1[15]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][16]  (.CLK(clk),
    .D(u0_n_29374),
    .QN(w1[16]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][17]  (.CLK(clk),
    .D(u0_n_29542),
    .QN(w1[17]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][18]  (.CLK(clk),
    .D(u0_n_29417),
    .QN(w1[18]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][19]  (.CLK(clk),
    .D(u0_n_29385),
    .QN(w1[19]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][1]  (.CLK(clk),
    .D(u0_n_29486),
    .QN(w1[1]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][20]  (.CLK(clk),
    .D(u0_n_29490),
    .QN(w1[20]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][21]  (.CLK(clk),
    .D(u0_n_29398),
    .QN(w1[21]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][22]  (.CLK(clk),
    .D(u0_n_29384),
    .QN(w1[22]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][23]  (.CLK(clk),
    .D(u0_n_29460),
    .QN(w1[23]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][24]  (.CLK(clk),
    .D(u0_n_29297),
    .QN(w1[24]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][25]  (.CLK(clk),
    .D(u0_n_29543),
    .QN(w1[25]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[1][26]  (.CLK(clk),
    .D(u0_n_29288),
    .QN(w1[26]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][27]  (.CLK(clk),
    .D(u0_n_29399),
    .QN(w1[27]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][28]  (.CLK(clk),
    .D(u0_n_29326),
    .QN(w1[28]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][29]  (.CLK(clk),
    .D(u0_n_29400),
    .QN(w1[29]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[1][2]  (.CLK(clk),
    .D(u0_n_29335),
    .QN(w1[2]));
 DFFHQNx2_ASAP7_75t_SL \u0_w_reg[1][30]  (.CLK(clk),
    .D(u0_n_29286),
    .QN(w1[30]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][31]  (.CLK(clk),
    .D(u0_n_29402),
    .QN(w1[31]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][3]  (.CLK(clk),
    .D(u0_n_29388),
    .QN(w1[3]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[1][4]  (.CLK(clk),
    .D(u0_n_29336),
    .QN(w1[4]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][5]  (.CLK(clk),
    .D(u0_n_29387),
    .QN(w1[5]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][6]  (.CLK(clk),
    .D(u0_n_29321),
    .QN(w1[6]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[1][7]  (.CLK(clk),
    .D(u0_n_29371),
    .QN(w1[7]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][8]  (.CLK(clk),
    .D(u0_n_29377),
    .QN(w1[8]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[1][9]  (.CLK(clk),
    .D(u0_n_29487),
    .QN(w1[9]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][0]  (.CLK(clk),
    .D(u0_n_29298),
    .QN(w2[0]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][10]  (.CLK(clk),
    .D(u0_n_29383),
    .QN(w2[10]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][11]  (.CLK(clk),
    .D(u0_n_29287),
    .QN(w2[11]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][12]  (.CLK(clk),
    .D(u0_n_29343),
    .QN(w2[12]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][13]  (.CLK(clk),
    .D(u0_n_29300),
    .QN(w2[13]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][14]  (.CLK(clk),
    .D(u0_n_29382),
    .QN(w2[14]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][15]  (.CLK(clk),
    .D(u0_n_29328),
    .QN(w2[15]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][16]  (.CLK(clk),
    .D(u0_n_29301),
    .QN(w2[16]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][17]  (.CLK(clk),
    .D(u0_n_29406),
    .QN(w2[17]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][18]  (.CLK(clk),
    .D(u0_n_29290),
    .QN(w2[18]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][19]  (.CLK(clk),
    .D(u0_n_29407),
    .QN(w2[19]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][1]  (.CLK(clk),
    .D(u0_n_29338),
    .QN(w2[1]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][20]  (.CLK(clk),
    .D(u0_n_29329),
    .QN(w2[20]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[2][21]  (.CLK(clk),
    .D(u0_n_29302),
    .QN(w2[21]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[2][22]  (.CLK(clk),
    .D(u0_n_29408),
    .QN(w2[22]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][23]  (.CLK(clk),
    .D(u0_n_29492),
    .QN(w2[23]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][24]  (.CLK(clk),
    .D(u0_n_29279),
    .QN(w2[24]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][25]  (.CLK(clk),
    .D(u0_n_29409),
    .QN(w2[25]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][26]  (.CLK(clk),
    .D(u0_n_29291),
    .QN(w2[26]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][27]  (.CLK(clk),
    .D(u0_n_29292),
    .QN(w2[27]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][28]  (.CLK(clk),
    .D(u0_n_29303),
    .QN(w2[28]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][29]  (.CLK(clk),
    .D(u0_n_29293),
    .QN(w2[29]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][2]  (.CLK(clk),
    .D(u0_n_29285),
    .QN(w2[2]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][30]  (.CLK(clk),
    .D(u0_n_29283),
    .QN(w2[30]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][31]  (.CLK(clk),
    .D(u0_n_29294),
    .QN(w2[31]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][3]  (.CLK(clk),
    .D(u0_n_29403),
    .QN(w2[3]));
 DFFHQNx1_ASAP7_75t_SL \u0_w_reg[2][4]  (.CLK(clk),
    .D(u0_n_29284),
    .QN(w2[4]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][5]  (.CLK(clk),
    .D(u0_n_29404),
    .QN(w2[5]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[2][6]  (.CLK(clk),
    .D(u0_n_29339),
    .QN(w2[6]));
 DFFHQNx1_ASAP7_75t_L \u0_w_reg[2][7]  (.CLK(clk),
    .D(u0_n_29341),
    .QN(w2[7]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[2][8]  (.CLK(clk),
    .D(u0_n_29299),
    .QN(w2[8]));
 DFFHQNx1_ASAP7_75t_R \u0_w_reg[2][9]  (.CLK(clk),
    .D(u0_n_29342),
    .QN(w2[9]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][0]  (.CLK(clk),
    .D(u0_n_29308),
    .QN(w3[0]),
    .SE(u0_n_32834),
    .SI(u0_n_32803));
 DFFHQx4_ASAP7_75t_SL \u0_w_reg[3][10]  (.CLK(clk),
    .D(u0_n_29381),
    .Q(w3[10]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][11]  (.CLK(clk),
    .D(u0_n_32805),
    .QN(w3[11]),
    .SE(u0_n_32835),
    .SI(u0_n_29435));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][12]  (.CLK(clk),
    .D(u0_n_29360),
    .QN(\u0_w[3] [12]),
    .SE(u0_n_32845),
    .SI(u0_n_32797));
 DFFHQx4_ASAP7_75t_L \u0_w_reg[3][13]  (.CLK(clk),
    .D(u0_n_29280),
    .Q(w3[13]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][14]  (.CLK(clk),
    .D(u0_n_29570),
    .QN(w3[14]),
    .SE(u0_n_32825),
    .SI(u0_n_32821));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][15]  (.CLK(clk),
    .D(u0_n_32819),
    .QN(w3[15]),
    .SE(u0_n_32875),
    .SI(u0_n_29363));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][16]  (.CLK(clk),
    .D(u0_n_32807),
    .QN(\u0_w[3] [16]),
    .SE(u0_n_32835),
    .SI(u0_n_29314));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][17]  (.CLK(clk),
    .D(u0_n_32817),
    .QN(w3[17]),
    .SE(u0_n_32875),
    .SI(u0_n_29429));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][18]  (.CLK(clk),
    .D(u0_n_29431),
    .QN(w3[18]),
    .SE(u0_n_32834),
    .SI(u0_n_32814));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][19]  (.CLK(clk),
    .D(u0_n_32813),
    .QN(w3[19]),
    .SE(u0_n_32875),
    .SI(u0_n_29444));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][1]  (.CLK(clk),
    .D(u0_n_32820),
    .QN(w3[1]),
    .SE(u0_n_32839),
    .SI(u0_n_29353));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][20]  (.CLK(clk),
    .D(u0_n_29496),
    .QN(w3[20]),
    .SE(u0_n_32845),
    .SI(u0_n_32804));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][21]  (.CLK(clk),
    .D(u0_n_29317),
    .QN(w3[21]),
    .SE(u0_n_32845),
    .SI(u0_n_32802));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][22]  (.CLK(clk),
    .D(u0_n_29411),
    .QN(\u0_w[3] [22]),
    .SE(u0_n_32845),
    .SI(u0_n_32812));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][23]  (.CLK(clk),
    .D(u0_n_32816),
    .QN(w3[23]),
    .SE(u0_n_32875),
    .SI(u0_n_29494));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][24]  (.CLK(clk),
    .D(u0_n_29320),
    .QN(w3[24]),
    .SE(u0_n_32845),
    .SI(u0_n_32798));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][25]  (.CLK(clk),
    .D(u0_n_32800),
    .QN(w3[25]),
    .SE(u0_n_32875),
    .SI(u0_n_29432));
 DFFHQx4_ASAP7_75t_SL \u0_w_reg[3][26]  (.CLK(clk),
    .D(u0_n_29296),
    .Q(w3[26]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][27]  (.CLK(clk),
    .D(u0_n_29434),
    .QN(\u0_w[3] [27]),
    .SE(u0_n_32834),
    .SI(u0_n_32810));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][28]  (.CLK(clk),
    .D(u0_n_29348),
    .QN(w3[28]),
    .SE(u0_n_32834),
    .SI(u0_n_32808));
 DFFHQx4_ASAP7_75t_L \u0_w_reg[3][29]  (.CLK(clk),
    .D(u0_n_29289),
    .Q(w3[29]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][2]  (.CLK(clk),
    .D(u0_n_29355),
    .QN(w3[2]),
    .SE(u0_n_32834),
    .SI(u0_n_32799));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][30]  (.CLK(clk),
    .D(u0_n_29344),
    .QN(\u0_w[3] [30]),
    .SE(u0_n_32845),
    .SI(u0_n_32818));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][31]  (.CLK(clk),
    .D(u0_n_29410),
    .QN(w3[31]),
    .SE(u0_n_32834),
    .SI(u0_n_32809));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][3]  (.CLK(clk),
    .D(u0_n_29441),
    .QN(w3[3]),
    .SE(u0_n_32825),
    .SI(u0_n_32811));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][4]  (.CLK(clk),
    .D(u0_n_29356),
    .QN(w3[4]),
    .SE(u0_n_32834),
    .SI(u0_n_32801));
 DFFHQx4_ASAP7_75t_SL \u0_w_reg[3][5]  (.CLK(clk),
    .D(u0_n_29295),
    .Q(w3[5]));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][6]  (.CLK(clk),
    .D(u0_n_29324),
    .QN(w3[6]),
    .SE(u0_n_32845),
    .SI(u0_n_32806));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][7]  (.CLK(clk),
    .D(u0_n_32822),
    .QN(w3[7]),
    .SE(u0_n_32875),
    .SI(u0_n_29369));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][8]  (.CLK(clk),
    .D(u0_n_29311),
    .QN(w3[8]),
    .SE(u0_n_32845),
    .SI(u0_n_32815));
 SDFHx4_ASAP7_75t_SL \u0_w_reg[3][9]  (.CLK(clk),
    .D(u0_n_29357),
    .QN(w3[9]),
    .SE(u0_n_32834),
    .SI(u0_n_32796));
endmodule
