module NV_NVDLA_partition_m (cmac_a2csb_resp_valid,
    csb2cmac_a_req_pvld,
    direct_reset_,
    dla_reset_rstn,
    global_clk_ovr_on,
    mac2accu_pvld,
    nvdla_clk_ovr_on,
    nvdla_core_clk,
    csb2cmac_a_req_prdy,
    sc2mac_dat_pvld,
    sc2mac_wt_pvld,
    test_mode,
    tmc2slcg_disable_clock_gating,
    mac2accu_mode,
    cmac_a2csb_resp_pd,
    csb2cmac_a_req_pd,
    mac2accu_data0,
    mac2accu_data1,
    mac2accu_data2,
    mac2accu_data3,
    mac2accu_mask,
    mac2accu_pd,
    sc2mac_dat_data0,
    sc2mac_dat_data1,
    sc2mac_dat_data2,
    sc2mac_dat_data3,
    sc2mac_dat_data4,
    sc2mac_dat_data5,
    sc2mac_dat_data6,
    sc2mac_dat_data7,
    sc2mac_dat_mask,
    sc2mac_dat_pd,
    sc2mac_wt_data0,
    sc2mac_wt_data1,
    sc2mac_wt_data2,
    sc2mac_wt_data3,
    sc2mac_wt_data4,
    sc2mac_wt_data5,
    sc2mac_wt_data6,
    sc2mac_wt_data7,
    sc2mac_wt_mask,
    sc2mac_wt_sel);
 output cmac_a2csb_resp_valid;
 input csb2cmac_a_req_pvld;
 input direct_reset_;
 input dla_reset_rstn;
 input global_clk_ovr_on;
 output mac2accu_pvld;
 input nvdla_clk_ovr_on;
 input nvdla_core_clk;
 output csb2cmac_a_req_prdy;
 input sc2mac_dat_pvld;
 input sc2mac_wt_pvld;
 input test_mode;
 input tmc2slcg_disable_clock_gating;
 output mac2accu_mode;
 output [33:0] cmac_a2csb_resp_pd;
 input [62:0] csb2cmac_a_req_pd;
 output [18:0] mac2accu_data0;
 output [18:0] mac2accu_data1;
 output [18:0] mac2accu_data2;
 output [18:0] mac2accu_data3;
 output [3:0] mac2accu_mask;
 output [8:0] mac2accu_pd;
 input [7:0] sc2mac_dat_data0;
 input [7:0] sc2mac_dat_data1;
 input [7:0] sc2mac_dat_data2;
 input [7:0] sc2mac_dat_data3;
 input [7:0] sc2mac_dat_data4;
 input [7:0] sc2mac_dat_data5;
 input [7:0] sc2mac_dat_data6;
 input [7:0] sc2mac_dat_data7;
 input [7:0] sc2mac_dat_mask;
 input [8:0] sc2mac_dat_pd;
 input [7:0] sc2mac_wt_data0;
 input [7:0] sc2mac_wt_data1;
 input [7:0] sc2mac_wt_data2;
 input [7:0] sc2mac_wt_data3;
 input [7:0] sc2mac_wt_data4;
 input [7:0] sc2mac_wt_data5;
 input [7:0] sc2mac_wt_data6;
 input [7:0] sc2mac_wt_data7;
 input [7:0] sc2mac_wt_mask;
 input [3:0] sc2mac_wt_sel;

 wire UNCONNECTED;
 wire UNCONNECTED0;
 wire UNCONNECTED1;
 wire UNCONNECTED10;
 wire UNCONNECTED11;
 wire UNCONNECTED12;
 wire UNCONNECTED13;
 wire UNCONNECTED14;
 wire UNCONNECTED15;
 wire UNCONNECTED16;
 wire UNCONNECTED17;
 wire UNCONNECTED18;
 wire UNCONNECTED19;
 wire UNCONNECTED2;
 wire UNCONNECTED20;
 wire UNCONNECTED21;
 wire UNCONNECTED22;
 wire UNCONNECTED23;
 wire UNCONNECTED24;
 wire UNCONNECTED25;
 wire UNCONNECTED26;
 wire UNCONNECTED27;
 wire UNCONNECTED28;
 wire UNCONNECTED29;
 wire UNCONNECTED3;
 wire UNCONNECTED30;
 wire UNCONNECTED4;
 wire UNCONNECTED5;
 wire UNCONNECTED6;
 wire UNCONNECTED7;
 wire UNCONNECTED8;
 wire UNCONNECTED9;
 wire n_10;
 wire n_1000;
 wire n_10005;
 wire n_10009;
 wire n_1001;
 wire n_10012;
 wire n_10013;
 wire n_10014;
 wire n_1002;
 wire n_10029;
 wire n_1003;
 wire n_10032;
 wire n_10033;
 wire n_10038;
 wire n_10039;
 wire n_1004;
 wire n_10044;
 wire n_10046;
 wire n_1005;
 wire n_10053;
 wire n_10054;
 wire n_10055;
 wire n_10056;
 wire n_10057;
 wire n_1006;
 wire n_10068;
 wire n_10069;
 wire n_1007;
 wire n_10070;
 wire n_10071;
 wire n_10073;
 wire n_10078;
 wire n_1008;
 wire n_10081;
 wire n_10082;
 wire n_10083;
 wire n_10084;
 wire n_10085;
 wire n_10086;
 wire n_1009;
 wire n_10090;
 wire n_10091;
 wire n_10092;
 wire n_10093;
 wire n_10094;
 wire n_10097;
 wire n_10098;
 wire n_10099;
 wire n_101;
 wire n_1010;
 wire n_10100;
 wire n_10102;
 wire n_10103;
 wire n_10104;
 wire n_10106;
 wire n_1011;
 wire n_10114;
 wire n_10115;
 wire n_10116;
 wire n_10117;
 wire n_1012;
 wire n_10122;
 wire n_10125;
 wire n_10128;
 wire n_10129;
 wire n_1013;
 wire n_10130;
 wire n_10131;
 wire n_10136;
 wire n_10137;
 wire n_10138;
 wire n_10139;
 wire n_1014;
 wire n_10141;
 wire n_10142;
 wire n_10143;
 wire n_10144;
 wire n_1015;
 wire n_10153;
 wire n_10157;
 wire n_10159;
 wire n_1016;
 wire n_10161;
 wire n_10162;
 wire n_10163;
 wire n_10169;
 wire n_1017;
 wire n_10171;
 wire n_10172;
 wire n_10173;
 wire n_10174;
 wire n_10175;
 wire n_10176;
 wire n_10177;
 wire n_1018;
 wire n_10180;
 wire n_10181;
 wire n_10182;
 wire n_10185;
 wire n_10187;
 wire n_10188;
 wire n_1019;
 wire n_10195;
 wire n_102;
 wire n_1020;
 wire n_10200;
 wire n_10201;
 wire n_10202;
 wire n_10205;
 wire n_10208;
 wire n_1021;
 wire n_10212;
 wire n_1022;
 wire n_10220;
 wire n_10224;
 wire n_10225;
 wire n_1023;
 wire n_10234;
 wire n_10235;
 wire n_10236;
 wire n_10237;
 wire n_10238;
 wire n_10239;
 wire n_1024;
 wire n_10240;
 wire n_10241;
 wire n_10242;
 wire n_10243;
 wire n_10247;
 wire n_10248;
 wire n_10249;
 wire n_1025;
 wire n_10255;
 wire n_10256;
 wire n_10257;
 wire n_10258;
 wire n_1026;
 wire n_10260;
 wire n_10261;
 wire n_10262;
 wire n_10263;
 wire n_10264;
 wire n_10265;
 wire n_10266;
 wire n_10267;
 wire n_1027;
 wire n_10271;
 wire n_10272;
 wire n_10274;
 wire n_10276;
 wire n_10278;
 wire n_10279;
 wire n_1028;
 wire n_10280;
 wire n_10281;
 wire n_10283;
 wire n_10284;
 wire n_10286;
 wire n_1029;
 wire n_10290;
 wire n_10291;
 wire n_10294;
 wire n_10295;
 wire n_10298;
 wire n_10299;
 wire n_103;
 wire n_1030;
 wire n_10301;
 wire n_10302;
 wire n_10303;
 wire n_10305;
 wire n_10307;
 wire n_10309;
 wire n_1031;
 wire n_10311;
 wire n_10318;
 wire n_10319;
 wire n_1032;
 wire n_10320;
 wire n_10321;
 wire n_10322;
 wire n_10324;
 wire n_10325;
 wire n_10326;
 wire n_10327;
 wire n_10328;
 wire n_10329;
 wire n_1033;
 wire n_10333;
 wire n_10334;
 wire n_10338;
 wire n_1034;
 wire n_10340;
 wire n_10344;
 wire n_10346;
 wire n_10348;
 wire n_1035;
 wire n_10350;
 wire n_10355;
 wire n_10356;
 wire n_10359;
 wire n_1036;
 wire n_10360;
 wire n_10368;
 wire n_10369;
 wire n_1037;
 wire n_10370;
 wire n_10374;
 wire n_10375;
 wire n_10376;
 wire n_10378;
 wire n_10379;
 wire n_1038;
 wire n_10387;
 wire n_10389;
 wire n_1039;
 wire n_10393;
 wire n_10394;
 wire n_10395;
 wire n_104;
 wire n_1040;
 wire n_10408;
 wire n_1041;
 wire n_10411;
 wire n_10414;
 wire n_10416;
 wire n_10417;
 wire n_10419;
 wire n_1042;
 wire n_10421;
 wire n_10423;
 wire n_10427;
 wire n_10429;
 wire n_1043;
 wire n_1044;
 wire n_10442;
 wire n_10443;
 wire n_10444;
 wire n_10445;
 wire n_10446;
 wire n_1045;
 wire n_10455;
 wire n_10456;
 wire n_1046;
 wire n_10465;
 wire n_10466;
 wire n_10469;
 wire n_1047;
 wire n_10470;
 wire n_10471;
 wire n_10472;
 wire n_10475;
 wire n_10476;
 wire n_10477;
 wire n_10478;
 wire n_10479;
 wire n_1048;
 wire n_10480;
 wire n_10481;
 wire n_10482;
 wire n_10483;
 wire n_1049;
 wire n_10490;
 wire n_10492;
 wire n_10499;
 wire n_105;
 wire n_1050;
 wire n_10500;
 wire n_10501;
 wire n_10503;
 wire n_10505;
 wire n_10506;
 wire n_10509;
 wire n_10512;
 wire n_10513;
 wire n_10515;
 wire n_10516;
 wire n_10520;
 wire n_10521;
 wire n_10522;
 wire n_10523;
 wire n_10527;
 wire n_10532;
 wire n_10533;
 wire n_10536;
 wire n_10537;
 wire n_10538;
 wire n_10541;
 wire n_10542;
 wire n_10543;
 wire n_10544;
 wire n_1055;
 wire n_10557;
 wire n_10558;
 wire n_1056;
 wire n_10560;
 wire n_10561;
 wire n_10563;
 wire n_10564;
 wire n_10567;
 wire n_10568;
 wire n_10569;
 wire n_1057;
 wire n_1058;
 wire n_10582;
 wire n_10585;
 wire n_10588;
 wire n_1059;
 wire n_10591;
 wire n_10592;
 wire n_10593;
 wire n_10594;
 wire n_10595;
 wire n_106;
 wire n_10601;
 wire n_10608;
 wire n_1061;
 wire n_10611;
 wire n_10612;
 wire n_10613;
 wire n_10617;
 wire n_10618;
 wire n_1062;
 wire n_10621;
 wire n_10622;
 wire n_10623;
 wire n_10627;
 wire n_10628;
 wire n_10629;
 wire n_1063;
 wire n_10635;
 wire n_1064;
 wire n_10640;
 wire n_10641;
 wire n_10642;
 wire n_10643;
 wire n_10645;
 wire n_10646;
 wire n_10647;
 wire n_10648;
 wire n_1065;
 wire n_10650;
 wire n_10657;
 wire n_1066;
 wire n_10665;
 wire n_10666;
 wire n_1067;
 wire n_10676;
 wire n_10677;
 wire n_1068;
 wire n_10684;
 wire n_10685;
 wire n_10686;
 wire n_10693;
 wire n_10694;
 wire n_10696;
 wire n_10697;
 wire n_107;
 wire n_1070;
 wire n_1071;
 wire n_10711;
 wire n_10713;
 wire n_10718;
 wire n_10719;
 wire n_1072;
 wire n_10720;
 wire n_10721;
 wire n_10723;
 wire n_10725;
 wire n_10728;
 wire n_1073;
 wire n_10730;
 wire n_10731;
 wire n_10732;
 wire n_10734;
 wire n_10736;
 wire n_10737;
 wire n_10738;
 wire n_10739;
 wire n_1074;
 wire n_10740;
 wire n_10741;
 wire n_10742;
 wire n_10744;
 wire n_10745;
 wire n_1075;
 wire n_10752;
 wire n_10753;
 wire n_10754;
 wire n_10755;
 wire n_10756;
 wire n_10757;
 wire n_10758;
 wire n_10759;
 wire n_1076;
 wire n_10760;
 wire n_10762;
 wire n_10765;
 wire n_1077;
 wire n_10771;
 wire n_10773;
 wire n_10774;
 wire n_10775;
 wire n_10776;
 wire n_10777;
 wire n_10778;
 wire n_1078;
 wire n_10788;
 wire n_10789;
 wire n_1079;
 wire n_10790;
 wire n_10791;
 wire n_10792;
 wire n_10793;
 wire n_10795;
 wire n_10796;
 wire n_10797;
 wire n_10798;
 wire n_10799;
 wire n_1080;
 wire n_10801;
 wire n_10802;
 wire n_10803;
 wire n_1081;
 wire n_10814;
 wire n_10816;
 wire n_1082;
 wire n_1083;
 wire n_10838;
 wire n_10839;
 wire n_1084;
 wire n_10840;
 wire n_10841;
 wire n_10842;
 wire n_10847;
 wire n_10848;
 wire n_1085;
 wire n_10856;
 wire n_10859;
 wire n_1086;
 wire n_10860;
 wire n_10862;
 wire n_10863;
 wire n_10864;
 wire n_10865;
 wire n_10866;
 wire n_1087;
 wire n_10878;
 wire n_1088;
 wire n_10882;
 wire n_10883;
 wire n_10885;
 wire n_10886;
 wire n_10887;
 wire n_10888;
 wire n_1089;
 wire n_10891;
 wire n_10892;
 wire n_10894;
 wire n_10895;
 wire n_1090;
 wire n_10901;
 wire n_10902;
 wire n_10903;
 wire n_10904;
 wire n_10905;
 wire n_10908;
 wire n_1091;
 wire n_10912;
 wire n_10913;
 wire n_10915;
 wire n_10916;
 wire n_10917;
 wire n_10918;
 wire n_1092;
 wire n_10922;
 wire n_1093;
 wire n_10933;
 wire n_1094;
 wire n_10947;
 wire n_1095;
 wire n_10953;
 wire n_10954;
 wire n_1096;
 wire n_10963;
 wire n_10964;
 wire n_10965;
 wire n_10968;
 wire n_10969;
 wire n_1097;
 wire n_10970;
 wire n_10971;
 wire n_10972;
 wire n_10973;
 wire n_1098;
 wire n_10981;
 wire n_10982;
 wire n_10983;
 wire n_1099;
 wire n_10990;
 wire n_10992;
 wire n_10993;
 wire n_10994;
 wire n_10995;
 wire n_10998;
 wire n_10999;
 wire n_11;
 wire n_1100;
 wire n_11000;
 wire n_1101;
 wire n_1102;
 wire n_11021;
 wire n_11022;
 wire n_11023;
 wire n_11026;
 wire n_11027;
 wire n_11028;
 wire n_11029;
 wire n_1103;
 wire n_11031;
 wire n_11032;
 wire n_11033;
 wire n_11036;
 wire n_11039;
 wire n_1104;
 wire n_11040;
 wire n_11041;
 wire n_11042;
 wire n_11043;
 wire n_11044;
 wire n_11045;
 wire n_1105;
 wire n_11054;
 wire n_11056;
 wire n_11058;
 wire n_1106;
 wire n_11062;
 wire n_11063;
 wire n_11064;
 wire n_11065;
 wire n_11066;
 wire n_11067;
 wire n_11069;
 wire n_1107;
 wire n_11070;
 wire n_11071;
 wire n_11072;
 wire n_11077;
 wire n_11084;
 wire n_11085;
 wire n_11088;
 wire n_11090;
 wire n_11091;
 wire n_11092;
 wire n_11093;
 wire n_11094;
 wire n_11095;
 wire n_11096;
 wire n_11097;
 wire n_11098;
 wire n_111;
 wire n_11105;
 wire n_11108;
 wire n_1111;
 wire n_11112;
 wire n_11116;
 wire n_11120;
 wire n_11121;
 wire n_11124;
 wire n_11125;
 wire n_11126;
 wire n_11127;
 wire n_11128;
 wire n_11129;
 wire n_11130;
 wire n_11131;
 wire n_11132;
 wire n_11133;
 wire n_11134;
 wire n_11135;
 wire n_11136;
 wire n_11137;
 wire n_11138;
 wire n_11142;
 wire n_11145;
 wire n_1115;
 wire n_11151;
 wire n_11152;
 wire n_1116;
 wire n_11164;
 wire n_11165;
 wire n_11168;
 wire n_11169;
 wire n_1117;
 wire n_11175;
 wire n_11176;
 wire n_11177;
 wire n_11178;
 wire n_1118;
 wire n_11189;
 wire n_1119;
 wire n_11192;
 wire n_11193;
 wire n_11194;
 wire n_11195;
 wire n_11196;
 wire n_11197;
 wire n_11198;
 wire n_112;
 wire n_1120;
 wire n_11200;
 wire n_11201;
 wire n_11204;
 wire n_11208;
 wire n_11209;
 wire n_1121;
 wire n_11212;
 wire n_11213;
 wire n_11215;
 wire n_11216;
 wire n_11218;
 wire n_11219;
 wire n_1122;
 wire n_11220;
 wire n_1123;
 wire n_11235;
 wire n_11236;
 wire n_11238;
 wire n_1124;
 wire n_11241;
 wire n_11242;
 wire n_11243;
 wire n_11246;
 wire n_11248;
 wire n_11249;
 wire n_1126;
 wire n_11264;
 wire n_11266;
 wire n_11267;
 wire n_11268;
 wire n_11269;
 wire n_1127;
 wire n_11270;
 wire n_11277;
 wire n_1128;
 wire n_11289;
 wire n_1129;
 wire n_11295;
 wire n_11298;
 wire n_11299;
 wire n_113;
 wire n_1130;
 wire n_11300;
 wire n_11302;
 wire n_11304;
 wire n_11307;
 wire n_11308;
 wire n_11309;
 wire n_1131;
 wire n_11310;
 wire n_11315;
 wire n_11316;
 wire n_11317;
 wire n_11318;
 wire n_1132;
 wire n_11320;
 wire n_11321;
 wire n_11322;
 wire n_11323;
 wire n_11324;
 wire n_11325;
 wire n_11326;
 wire n_11327;
 wire n_11328;
 wire n_1133;
 wire n_11332;
 wire n_11333;
 wire n_11334;
 wire n_11338;
 wire n_11339;
 wire n_1134;
 wire n_11340;
 wire n_11341;
 wire n_11343;
 wire n_11346;
 wire n_11348;
 wire n_1135;
 wire n_11350;
 wire n_11356;
 wire n_11357;
 wire n_11359;
 wire n_1136;
 wire n_11361;
 wire n_1137;
 wire n_11374;
 wire n_11375;
 wire n_11376;
 wire n_11377;
 wire n_11379;
 wire n_1138;
 wire n_11381;
 wire n_11382;
 wire n_11383;
 wire n_11384;
 wire n_11385;
 wire n_11386;
 wire n_11387;
 wire n_11388;
 wire n_11389;
 wire n_1139;
 wire n_114;
 wire n_1140;
 wire n_11401;
 wire n_11403;
 wire n_11404;
 wire n_11405;
 wire n_11409;
 wire n_1141;
 wire n_11411;
 wire n_11412;
 wire n_11413;
 wire n_11417;
 wire n_11418;
 wire n_11419;
 wire n_1142;
 wire n_11421;
 wire n_11423;
 wire n_11424;
 wire n_11425;
 wire n_11427;
 wire n_11428;
 wire n_11429;
 wire n_1143;
 wire n_11430;
 wire n_11431;
 wire n_11433;
 wire n_11438;
 wire n_1144;
 wire n_11444;
 wire n_11445;
 wire n_11446;
 wire n_11449;
 wire n_11450;
 wire n_11451;
 wire n_11452;
 wire n_11453;
 wire n_11454;
 wire n_11455;
 wire n_11456;
 wire n_11458;
 wire n_1146;
 wire n_11462;
 wire n_11463;
 wire n_11469;
 wire n_1147;
 wire n_11471;
 wire n_11472;
 wire n_11473;
 wire n_11474;
 wire n_11475;
 wire n_11476;
 wire n_11477;
 wire n_11479;
 wire n_1148;
 wire n_11480;
 wire n_11481;
 wire n_11483;
 wire n_11487;
 wire n_11489;
 wire n_1149;
 wire n_11490;
 wire n_11492;
 wire n_11493;
 wire n_11495;
 wire n_11496;
 wire n_1150;
 wire n_11501;
 wire n_11502;
 wire n_11509;
 wire n_1151;
 wire n_11510;
 wire n_11515;
 wire n_11517;
 wire n_11519;
 wire n_1152;
 wire n_11520;
 wire n_11521;
 wire n_11525;
 wire n_11526;
 wire n_11527;
 wire n_11528;
 wire n_11529;
 wire n_1153;
 wire n_11533;
 wire n_11534;
 wire n_11535;
 wire n_11536;
 wire n_11537;
 wire n_11538;
 wire n_11539;
 wire n_1154;
 wire n_11540;
 wire n_11541;
 wire n_11542;
 wire n_11543;
 wire n_11544;
 wire n_11545;
 wire n_11546;
 wire n_11547;
 wire n_1155;
 wire n_11550;
 wire n_1156;
 wire n_11568;
 wire n_1157;
 wire n_11570;
 wire n_11571;
 wire n_11573;
 wire n_11574;
 wire n_11575;
 wire n_11576;
 wire n_11578;
 wire n_11579;
 wire n_1158;
 wire n_11580;
 wire n_11581;
 wire n_11582;
 wire n_11583;
 wire n_11584;
 wire n_11585;
 wire n_11586;
 wire n_11587;
 wire n_1159;
 wire n_11590;
 wire n_11592;
 wire n_11593;
 wire n_11596;
 wire n_11597;
 wire n_11598;
 wire n_11599;
 wire n_116;
 wire n_1160;
 wire n_1161;
 wire n_11610;
 wire n_11611;
 wire n_11612;
 wire n_11618;
 wire n_1162;
 wire n_11620;
 wire n_11621;
 wire n_11622;
 wire n_11625;
 wire n_11627;
 wire n_1163;
 wire n_11630;
 wire n_11638;
 wire n_1164;
 wire n_11644;
 wire n_1165;
 wire n_1166;
 wire n_1167;
 wire n_1168;
 wire n_1169;
 wire n_117;
 wire n_11722;
 wire n_11723;
 wire n_11725;
 wire n_11726;
 wire n_11729;
 wire n_11739;
 wire n_11742;
 wire n_11743;
 wire n_11746;
 wire n_11751;
 wire n_11752;
 wire n_11753;
 wire n_1176;
 wire n_11760;
 wire n_11761;
 wire n_11762;
 wire n_11763;
 wire n_11767;
 wire n_11768;
 wire n_11770;
 wire n_11771;
 wire n_1178;
 wire n_11781;
 wire n_11783;
 wire n_11787;
 wire n_11788;
 wire n_11789;
 wire n_11790;
 wire n_11791;
 wire n_11793;
 wire n_118;
 wire n_1180;
 wire n_11800;
 wire n_11808;
 wire n_1181;
 wire n_11812;
 wire n_11818;
 wire n_11819;
 wire n_1182;
 wire n_11821;
 wire n_11822;
 wire n_11823;
 wire n_11826;
 wire n_11827;
 wire n_11828;
 wire n_11829;
 wire n_1183;
 wire n_11830;
 wire n_11832;
 wire n_11833;
 wire n_11835;
 wire n_1184;
 wire n_11845;
 wire n_11846;
 wire n_1185;
 wire n_11852;
 wire n_11854;
 wire n_11855;
 wire n_11856;
 wire n_11857;
 wire n_11858;
 wire n_1186;
 wire n_11865;
 wire n_11867;
 wire n_11868;
 wire n_11869;
 wire n_1187;
 wire n_11871;
 wire n_11872;
 wire n_1188;
 wire n_11887;
 wire n_1189;
 wire n_11891;
 wire n_11892;
 wire n_11896;
 wire n_119;
 wire n_1190;
 wire n_11904;
 wire n_1191;
 wire n_11912;
 wire n_11913;
 wire n_11914;
 wire n_11915;
 wire n_11916;
 wire n_11918;
 wire n_11919;
 wire n_1192;
 wire n_11920;
 wire n_11924;
 wire n_11925;
 wire n_11928;
 wire n_1193;
 wire n_11930;
 wire n_11931;
 wire n_11932;
 wire n_11936;
 wire n_11937;
 wire n_1194;
 wire n_11941;
 wire n_11942;
 wire n_11943;
 wire n_11944;
 wire n_11945;
 wire n_1195;
 wire n_1196;
 wire n_11960;
 wire n_11961;
 wire n_11962;
 wire n_11963;
 wire n_11964;
 wire n_11965;
 wire n_11966;
 wire n_11967;
 wire n_11968;
 wire n_1197;
 wire n_11970;
 wire n_11972;
 wire n_1198;
 wire n_11984;
 wire n_1199;
 wire n_11995;
 wire n_11996;
 wire n_11997;
 wire n_11998;
 wire n_11999;
 wire n_12;
 wire n_120;
 wire n_1200;
 wire n_12000;
 wire n_12001;
 wire n_1201;
 wire n_12013;
 wire n_12016;
 wire n_12017;
 wire n_12018;
 wire n_1202;
 wire n_12023;
 wire n_12025;
 wire n_12026;
 wire n_12027;
 wire n_12028;
 wire n_1203;
 wire n_12033;
 wire n_12035;
 wire n_12036;
 wire n_12038;
 wire n_12039;
 wire n_1204;
 wire n_1205;
 wire n_12050;
 wire n_12051;
 wire n_12056;
 wire n_1206;
 wire n_12061;
 wire n_12062;
 wire n_12063;
 wire n_12064;
 wire n_12065;
 wire n_12066;
 wire n_12067;
 wire n_12068;
 wire n_12069;
 wire n_1207;
 wire n_12073;
 wire n_12077;
 wire n_12079;
 wire n_1208;
 wire n_12080;
 wire n_12087;
 wire n_12088;
 wire n_1209;
 wire n_12091;
 wire n_1210;
 wire n_12101;
 wire n_12107;
 wire n_12108;
 wire n_1211;
 wire n_12110;
 wire n_12111;
 wire n_12114;
 wire n_1212;
 wire n_12120;
 wire n_12124;
 wire n_12129;
 wire n_1213;
 wire n_12134;
 wire n_1214;
 wire n_1215;
 wire n_12152;
 wire n_12154;
 wire n_1216;
 wire n_1217;
 wire n_1218;
 wire n_12186;
 wire n_12187;
 wire n_12188;
 wire n_1219;
 wire n_12190;
 wire n_12191;
 wire n_122;
 wire n_1220;
 wire n_1221;
 wire n_12213;
 wire n_12214;
 wire n_12215;
 wire n_12216;
 wire n_12217;
 wire n_12218;
 wire n_12219;
 wire n_1222;
 wire n_1223;
 wire n_1224;
 wire n_12245;
 wire n_12246;
 wire n_1225;
 wire n_12250;
 wire n_12251;
 wire n_12252;
 wire n_12254;
 wire n_12255;
 wire n_12257;
 wire n_12258;
 wire n_12259;
 wire n_1226;
 wire n_12260;
 wire n_12261;
 wire n_12262;
 wire n_12263;
 wire n_12264;
 wire n_12265;
 wire n_12266;
 wire n_12267;
 wire n_12271;
 wire n_12272;
 wire n_12276;
 wire n_12278;
 wire n_12279;
 wire n_1228;
 wire n_12281;
 wire n_12283;
 wire n_12284;
 wire n_12285;
 wire n_12286;
 wire n_12287;
 wire n_12288;
 wire n_12289;
 wire n_1229;
 wire n_12290;
 wire n_12293;
 wire n_123;
 wire n_1230;
 wire n_12301;
 wire n_12303;
 wire n_12304;
 wire n_12306;
 wire n_12307;
 wire n_12308;
 wire n_1236;
 wire n_1237;
 wire n_12374;
 wire n_12375;
 wire n_12376;
 wire n_12377;
 wire n_12379;
 wire n_1238;
 wire n_12380;
 wire n_12381;
 wire n_12382;
 wire n_12383;
 wire n_12384;
 wire n_12385;
 wire n_12386;
 wire n_12387;
 wire n_12388;
 wire n_12389;
 wire n_12390;
 wire n_12391;
 wire n_12392;
 wire n_12393;
 wire n_12394;
 wire n_12395;
 wire n_12397;
 wire n_12398;
 wire n_124;
 wire n_1240;
 wire n_12400;
 wire n_12402;
 wire n_1241;
 wire n_12411;
 wire n_12412;
 wire n_12414;
 wire n_12418;
 wire n_12419;
 wire n_1242;
 wire n_12420;
 wire n_12422;
 wire n_12424;
 wire n_12425;
 wire n_12427;
 wire n_12428;
 wire n_1243;
 wire n_1244;
 wire n_1245;
 wire n_1246;
 wire n_1247;
 wire n_1248;
 wire n_1249;
 wire n_12492;
 wire n_12494;
 wire n_12498;
 wire n_12499;
 wire n_125;
 wire n_12500;
 wire n_12503;
 wire n_12504;
 wire n_12508;
 wire n_1251;
 wire n_12510;
 wire n_12511;
 wire n_12512;
 wire n_12513;
 wire n_12514;
 wire n_12516;
 wire n_12518;
 wire n_1252;
 wire n_12520;
 wire n_12525;
 wire n_12526;
 wire n_12527;
 wire n_12528;
 wire n_1253;
 wire n_12530;
 wire n_12531;
 wire n_12532;
 wire n_1254;
 wire n_12540;
 wire n_12546;
 wire n_12547;
 wire n_12548;
 wire n_12549;
 wire n_1255;
 wire n_12550;
 wire n_12559;
 wire n_1256;
 wire n_12560;
 wire n_12561;
 wire n_12562;
 wire n_12563;
 wire n_12564;
 wire n_12565;
 wire n_12567;
 wire n_1257;
 wire n_12570;
 wire n_12571;
 wire n_12575;
 wire n_12576;
 wire n_12578;
 wire n_12579;
 wire n_1258;
 wire n_12580;
 wire n_12581;
 wire n_12583;
 wire n_12584;
 wire n_12589;
 wire n_1259;
 wire n_12591;
 wire n_12592;
 wire n_12593;
 wire n_12594;
 wire n_12595;
 wire n_12597;
 wire n_12598;
 wire n_126;
 wire n_1260;
 wire n_12603;
 wire n_12604;
 wire n_12605;
 wire n_12606;
 wire n_1261;
 wire n_12616;
 wire n_12618;
 wire n_1262;
 wire n_12620;
 wire n_12621;
 wire n_12622;
 wire n_12623;
 wire n_12624;
 wire n_12625;
 wire n_1263;
 wire n_12631;
 wire n_12632;
 wire n_12634;
 wire n_12637;
 wire n_12639;
 wire n_1264;
 wire n_12640;
 wire n_12641;
 wire n_12642;
 wire n_12643;
 wire n_12644;
 wire n_12648;
 wire n_12649;
 wire n_1265;
 wire n_12652;
 wire n_12653;
 wire n_12658;
 wire n_12659;
 wire n_1266;
 wire n_12661;
 wire n_12662;
 wire n_12663;
 wire n_12664;
 wire n_12665;
 wire n_12666;
 wire n_12667;
 wire n_12669;
 wire n_1267;
 wire n_12672;
 wire n_12674;
 wire n_12676;
 wire n_1268;
 wire n_12680;
 wire n_12681;
 wire n_12696;
 wire n_12697;
 wire n_12698;
 wire n_1270;
 wire n_12700;
 wire n_12701;
 wire n_12702;
 wire n_12703;
 wire n_12704;
 wire n_12705;
 wire n_12706;
 wire n_12707;
 wire n_12708;
 wire n_12709;
 wire n_1271;
 wire n_12712;
 wire n_12715;
 wire n_12717;
 wire n_12719;
 wire n_12720;
 wire n_1273;
 wire n_12738;
 wire n_12739;
 wire n_1274;
 wire n_12740;
 wire n_12744;
 wire n_12745;
 wire n_12746;
 wire n_12747;
 wire n_12748;
 wire n_12749;
 wire n_1275;
 wire n_12750;
 wire n_12752;
 wire n_12754;
 wire n_1276;
 wire n_1277;
 wire n_12774;
 wire n_12775;
 wire n_12778;
 wire n_12779;
 wire n_1278;
 wire n_12780;
 wire n_12781;
 wire n_12782;
 wire n_12785;
 wire n_12786;
 wire n_12787;
 wire n_1279;
 wire n_1280;
 wire n_12800;
 wire n_12801;
 wire n_12802;
 wire n_12803;
 wire n_12806;
 wire n_1281;
 wire n_12813;
 wire n_12814;
 wire n_12817;
 wire n_12818;
 wire n_12819;
 wire n_1282;
 wire n_12820;
 wire n_1283;
 wire n_12831;
 wire n_12833;
 wire n_12834;
 wire n_12839;
 wire n_1284;
 wire n_1285;
 wire n_1286;
 wire n_1287;
 wire n_12878;
 wire n_1288;
 wire n_12882;
 wire n_12884;
 wire n_12887;
 wire n_12888;
 wire n_1289;
 wire n_12892;
 wire n_12893;
 wire n_12894;
 wire n_12895;
 wire n_12896;
 wire n_12897;
 wire n_12899;
 wire n_129;
 wire n_1290;
 wire n_12900;
 wire n_12901;
 wire n_12902;
 wire n_12903;
 wire n_12904;
 wire n_12905;
 wire n_12906;
 wire n_1291;
 wire n_12917;
 wire n_12918;
 wire n_1292;
 wire n_12922;
 wire n_12923;
 wire n_12924;
 wire n_12926;
 wire n_12927;
 wire n_12928;
 wire n_12929;
 wire n_1293;
 wire n_12930;
 wire n_12931;
 wire n_12932;
 wire n_12933;
 wire n_12934;
 wire n_12935;
 wire n_12938;
 wire n_12939;
 wire n_1294;
 wire n_12940;
 wire n_12945;
 wire n_12948;
 wire n_1295;
 wire n_12956;
 wire n_12959;
 wire n_1296;
 wire n_12962;
 wire n_1297;
 wire n_12975;
 wire n_12978;
 wire n_12979;
 wire n_1298;
 wire n_12980;
 wire n_12981;
 wire n_12982;
 wire n_12984;
 wire n_12985;
 wire n_12986;
 wire n_12987;
 wire n_12988;
 wire n_1299;
 wire n_12990;
 wire n_12991;
 wire n_12993;
 wire n_12995;
 wire n_12996;
 wire n_12997;
 wire n_13;
 wire n_130;
 wire n_1300;
 wire n_13007;
 wire n_13008;
 wire n_13009;
 wire n_1301;
 wire n_13010;
 wire n_13011;
 wire n_13012;
 wire n_13013;
 wire n_13014;
 wire n_13015;
 wire n_13016;
 wire n_13017;
 wire n_1302;
 wire n_13021;
 wire n_13022;
 wire n_13023;
 wire n_13025;
 wire n_13028;
 wire n_1303;
 wire n_13030;
 wire n_13031;
 wire n_13033;
 wire n_13034;
 wire n_13036;
 wire n_13038;
 wire n_1304;
 wire n_13040;
 wire n_1305;
 wire n_13052;
 wire n_13053;
 wire n_13054;
 wire n_13056;
 wire n_13057;
 wire n_13059;
 wire n_1306;
 wire n_13060;
 wire n_13061;
 wire n_13065;
 wire n_13067;
 wire n_13069;
 wire n_1307;
 wire n_13071;
 wire n_13072;
 wire n_13079;
 wire n_1308;
 wire n_13080;
 wire n_13081;
 wire n_13082;
 wire n_13087;
 wire n_13088;
 wire n_13089;
 wire n_1309;
 wire n_13090;
 wire n_13091;
 wire n_13097;
 wire n_13098;
 wire n_131;
 wire n_1310;
 wire n_13100;
 wire n_13103;
 wire n_13104;
 wire n_13106;
 wire n_13107;
 wire n_1311;
 wire n_13111;
 wire n_13112;
 wire n_1312;
 wire n_13123;
 wire n_13124;
 wire n_13125;
 wire n_13126;
 wire n_13127;
 wire n_13128;
 wire n_13129;
 wire n_1313;
 wire n_13130;
 wire n_13133;
 wire n_13138;
 wire n_1314;
 wire n_13141;
 wire n_13142;
 wire n_13143;
 wire n_13144;
 wire n_13148;
 wire n_13149;
 wire n_1315;
 wire n_1316;
 wire n_1317;
 wire n_13172;
 wire n_13173;
 wire n_13175;
 wire n_13176;
 wire n_13178;
 wire n_1318;
 wire n_13181;
 wire n_13185;
 wire n_13186;
 wire n_13188;
 wire n_1319;
 wire n_13190;
 wire n_13191;
 wire n_13193;
 wire n_13196;
 wire n_132;
 wire n_1320;
 wire n_13201;
 wire n_13203;
 wire n_13204;
 wire n_1321;
 wire n_1322;
 wire n_13227;
 wire n_13228;
 wire n_1323;
 wire n_13230;
 wire n_13231;
 wire n_13233;
 wire n_13234;
 wire n_13235;
 wire n_13236;
 wire n_13237;
 wire n_13238;
 wire n_13239;
 wire n_1324;
 wire n_13240;
 wire n_13241;
 wire n_13242;
 wire n_13243;
 wire n_13244;
 wire n_13245;
 wire n_13247;
 wire n_13248;
 wire n_13249;
 wire n_1325;
 wire n_13250;
 wire n_13251;
 wire n_1326;
 wire n_1327;
 wire n_1328;
 wire n_13289;
 wire n_1329;
 wire n_13291;
 wire n_13292;
 wire n_13293;
 wire n_13294;
 wire n_13295;
 wire n_1330;
 wire n_1331;
 wire n_13319;
 wire n_1332;
 wire n_13321;
 wire n_13324;
 wire n_13327;
 wire n_13328;
 wire n_1333;
 wire n_13330;
 wire n_13331;
 wire n_13332;
 wire n_13333;
 wire n_1334;
 wire n_1335;
 wire n_13358;
 wire n_13359;
 wire n_1336;
 wire n_13360;
 wire n_13361;
 wire n_13362;
 wire n_13363;
 wire n_13364;
 wire n_1337;
 wire n_1338;
 wire n_13387;
 wire n_13389;
 wire n_1339;
 wire n_13390;
 wire n_13393;
 wire n_13397;
 wire n_134;
 wire n_1340;
 wire n_13401;
 wire n_13404;
 wire n_13405;
 wire n_13406;
 wire n_1341;
 wire n_13412;
 wire n_13413;
 wire n_13415;
 wire n_13416;
 wire n_13417;
 wire n_13418;
 wire n_13419;
 wire n_1342;
 wire n_13420;
 wire n_13423;
 wire n_1343;
 wire n_13435;
 wire n_13437;
 wire n_13439;
 wire n_1344;
 wire n_13440;
 wire n_13441;
 wire n_13447;
 wire n_13448;
 wire n_13449;
 wire n_1345;
 wire n_13450;
 wire n_13451;
 wire n_13456;
 wire n_13458;
 wire n_13459;
 wire n_1346;
 wire n_13464;
 wire n_13465;
 wire n_13467;
 wire n_1347;
 wire n_13474;
 wire n_13475;
 wire n_13476;
 wire n_13477;
 wire n_1348;
 wire n_13480;
 wire n_13481;
 wire n_13482;
 wire n_13483;
 wire n_13487;
 wire n_1349;
 wire n_13495;
 wire n_13498;
 wire n_13499;
 wire n_135;
 wire n_1350;
 wire n_13502;
 wire n_13504;
 wire n_13505;
 wire n_13508;
 wire n_1351;
 wire n_13519;
 wire n_1352;
 wire n_13521;
 wire n_13522;
 wire n_13523;
 wire n_13524;
 wire n_13525;
 wire n_1353;
 wire n_13530;
 wire n_13537;
 wire n_13538;
 wire n_13539;
 wire n_1354;
 wire n_13540;
 wire n_13541;
 wire n_13542;
 wire n_13543;
 wire n_13544;
 wire n_13546;
 wire n_1355;
 wire n_13551;
 wire n_13552;
 wire n_1356;
 wire n_13566;
 wire n_13567;
 wire n_1357;
 wire n_13570;
 wire n_13571;
 wire n_13572;
 wire n_13573;
 wire n_13574;
 wire n_13575;
 wire n_13576;
 wire n_13577;
 wire n_13578;
 wire n_1358;
 wire n_13586;
 wire n_13588;
 wire n_13589;
 wire n_1359;
 wire n_13590;
 wire n_13593;
 wire n_13596;
 wire n_13597;
 wire n_13598;
 wire n_13599;
 wire n_1360;
 wire n_13600;
 wire n_13602;
 wire n_13603;
 wire n_13605;
 wire n_13606;
 wire n_13608;
 wire n_13609;
 wire n_1361;
 wire n_13612;
 wire n_13616;
 wire n_13617;
 wire n_13619;
 wire n_1362;
 wire n_13621;
 wire n_13622;
 wire n_13623;
 wire n_13625;
 wire n_13627;
 wire n_13628;
 wire n_13629;
 wire n_1363;
 wire n_13631;
 wire n_13634;
 wire n_13635;
 wire n_13637;
 wire n_1364;
 wire n_13640;
 wire n_13641;
 wire n_13644;
 wire n_13645;
 wire n_13646;
 wire n_13647;
 wire n_13648;
 wire n_13649;
 wire n_1365;
 wire n_13650;
 wire n_13651;
 wire n_13652;
 wire n_13653;
 wire n_13654;
 wire n_13655;
 wire n_13656;
 wire n_13657;
 wire n_13658;
 wire n_1366;
 wire n_13667;
 wire n_1367;
 wire n_13674;
 wire n_13676;
 wire n_13678;
 wire n_1368;
 wire n_13681;
 wire n_13685;
 wire n_13687;
 wire n_13688;
 wire n_1369;
 wire n_13694;
 wire n_13697;
 wire n_13699;
 wire n_1370;
 wire n_13701;
 wire n_13702;
 wire n_13707;
 wire n_13708;
 wire n_13709;
 wire n_1371;
 wire n_13710;
 wire n_13711;
 wire n_13712;
 wire n_13716;
 wire n_13717;
 wire n_13718;
 wire n_13719;
 wire n_1372;
 wire n_13720;
 wire n_13721;
 wire n_13723;
 wire n_13724;
 wire n_13725;
 wire n_13726;
 wire n_13727;
 wire n_13728;
 wire n_1373;
 wire n_1374;
 wire n_1375;
 wire n_1376;
 wire n_13766;
 wire n_13767;
 wire n_13769;
 wire n_1377;
 wire n_13770;
 wire n_13771;
 wire n_13772;
 wire n_13773;
 wire n_13774;
 wire n_13776;
 wire n_13777;
 wire n_13778;
 wire n_13779;
 wire n_1378;
 wire n_13782;
 wire n_13784;
 wire n_13785;
 wire n_13786;
 wire n_13787;
 wire n_13788;
 wire n_13789;
 wire n_1379;
 wire n_13790;
 wire n_13791;
 wire n_13792;
 wire n_13793;
 wire n_13794;
 wire n_13795;
 wire n_13796;
 wire n_13797;
 wire n_138;
 wire n_1380;
 wire n_1381;
 wire n_1382;
 wire n_1383;
 wire n_1384;
 wire n_13843;
 wire n_13844;
 wire n_13845;
 wire n_13846;
 wire n_13848;
 wire n_1385;
 wire n_1386;
 wire n_1387;
 wire n_13873;
 wire n_13874;
 wire n_13877;
 wire n_13878;
 wire n_1388;
 wire n_13880;
 wire n_1389;
 wire n_139;
 wire n_1390;
 wire n_1391;
 wire n_1392;
 wire n_13929;
 wire n_1393;
 wire n_13930;
 wire n_13931;
 wire n_13932;
 wire n_13933;
 wire n_13934;
 wire n_13936;
 wire n_1394;
 wire n_13945;
 wire n_13946;
 wire n_13947;
 wire n_1395;
 wire n_13951;
 wire n_13952;
 wire n_13953;
 wire n_13958;
 wire n_13959;
 wire n_1396;
 wire n_13960;
 wire n_13966;
 wire n_13968;
 wire n_13969;
 wire n_1397;
 wire n_13970;
 wire n_13971;
 wire n_13975;
 wire n_1398;
 wire n_1399;
 wire n_14;
 wire n_140;
 wire n_1400;
 wire n_1401;
 wire n_14017;
 wire n_14018;
 wire n_14019;
 wire n_1402;
 wire n_14020;
 wire n_14021;
 wire n_14022;
 wire n_14024;
 wire n_14025;
 wire n_14029;
 wire n_1403;
 wire n_14031;
 wire n_14033;
 wire n_14035;
 wire n_14038;
 wire n_1404;
 wire n_14045;
 wire n_14048;
 wire n_14049;
 wire n_1405;
 wire n_14050;
 wire n_14059;
 wire n_1406;
 wire n_14061;
 wire n_14062;
 wire n_14063;
 wire n_14064;
 wire n_14067;
 wire n_1407;
 wire n_1408;
 wire n_14087;
 wire n_14088;
 wire n_14089;
 wire n_1409;
 wire n_14090;
 wire n_14091;
 wire n_14092;
 wire n_1410;
 wire n_14100;
 wire n_14101;
 wire n_14102;
 wire n_14103;
 wire n_14105;
 wire n_14106;
 wire n_14108;
 wire n_14109;
 wire n_1411;
 wire n_14110;
 wire n_14111;
 wire n_14115;
 wire n_14116;
 wire n_14117;
 wire n_14118;
 wire n_14120;
 wire n_14121;
 wire n_14122;
 wire n_14123;
 wire n_14124;
 wire n_14125;
 wire n_1413;
 wire n_14135;
 wire n_14136;
 wire n_14137;
 wire n_1414;
 wire n_14140;
 wire n_14141;
 wire n_14143;
 wire n_14147;
 wire n_1415;
 wire n_14151;
 wire n_14152;
 wire n_14153;
 wire n_14158;
 wire n_14159;
 wire n_1416;
 wire n_14162;
 wire n_1417;
 wire n_14172;
 wire n_14174;
 wire n_14176;
 wire n_14177;
 wire n_14179;
 wire n_1418;
 wire n_14181;
 wire n_14183;
 wire n_14186;
 wire n_1419;
 wire n_142;
 wire n_1420;
 wire n_14203;
 wire n_14204;
 wire n_14208;
 wire n_1421;
 wire n_14211;
 wire n_14213;
 wire n_1422;
 wire n_1423;
 wire n_14237;
 wire n_14238;
 wire n_1424;
 wire n_14241;
 wire n_14242;
 wire n_14243;
 wire n_14244;
 wire n_1425;
 wire n_1426;
 wire n_1427;
 wire n_1428;
 wire n_1429;
 wire n_14298;
 wire n_14299;
 wire n_143;
 wire n_1430;
 wire n_14300;
 wire n_14301;
 wire n_1431;
 wire n_1432;
 wire n_14327;
 wire n_14329;
 wire n_1433;
 wire n_14330;
 wire n_14333;
 wire n_14334;
 wire n_14335;
 wire n_14336;
 wire n_14339;
 wire n_1434;
 wire n_14340;
 wire n_14344;
 wire n_1435;
 wire n_14353;
 wire n_14354;
 wire n_14355;
 wire n_1436;
 wire n_14364;
 wire n_14367;
 wire n_14368;
 wire n_1437;
 wire n_14372;
 wire n_14373;
 wire n_1438;
 wire n_14382;
 wire n_14383;
 wire n_14384;
 wire n_14386;
 wire n_14388;
 wire n_1439;
 wire n_14394;
 wire n_144;
 wire n_1440;
 wire n_14407;
 wire n_14408;
 wire n_1441;
 wire n_14411;
 wire n_14412;
 wire n_14413;
 wire n_14414;
 wire n_14415;
 wire n_14416;
 wire n_14417;
 wire n_14418;
 wire n_1442;
 wire n_14425;
 wire n_14427;
 wire n_14429;
 wire n_1443;
 wire n_14430;
 wire n_14431;
 wire n_14434;
 wire n_14436;
 wire n_14437;
 wire n_14438;
 wire n_14439;
 wire n_1444;
 wire n_14440;
 wire n_14441;
 wire n_14442;
 wire n_14443;
 wire n_14444;
 wire n_14445;
 wire n_1445;
 wire n_14451;
 wire n_14452;
 wire n_14454;
 wire n_14456;
 wire n_14457;
 wire n_1446;
 wire n_1447;
 wire n_1448;
 wire n_1449;
 wire n_145;
 wire n_1450;
 wire n_1451;
 wire n_1452;
 wire n_14523;
 wire n_1453;
 wire n_14537;
 wire n_1454;
 wire n_1455;
 wire n_1456;
 wire n_1457;
 wire n_1458;
 wire n_1459;
 wire n_146;
 wire n_1460;
 wire n_1461;
 wire n_1462;
 wire n_1463;
 wire n_1464;
 wire n_14643;
 wire n_14645;
 wire n_1465;
 wire n_14652;
 wire n_14653;
 wire n_1466;
 wire n_14664;
 wire n_14669;
 wire n_1467;
 wire n_14671;
 wire n_14674;
 wire n_14675;
 wire n_1468;
 wire n_14683;
 wire n_14684;
 wire n_14687;
 wire n_14688;
 wire n_14689;
 wire n_1469;
 wire n_14695;
 wire n_14698;
 wire n_147;
 wire n_1470;
 wire n_14701;
 wire n_14702;
 wire n_14703;
 wire n_14704;
 wire n_14705;
 wire n_14706;
 wire n_14708;
 wire n_14709;
 wire n_1471;
 wire n_14713;
 wire n_14716;
 wire n_14717;
 wire n_14718;
 wire n_1472;
 wire n_14720;
 wire n_14721;
 wire n_14722;
 wire n_14723;
 wire n_14724;
 wire n_14725;
 wire n_14729;
 wire n_1473;
 wire n_14730;
 wire n_14731;
 wire n_14732;
 wire n_14733;
 wire n_14734;
 wire n_14735;
 wire n_14736;
 wire n_14739;
 wire n_1474;
 wire n_14740;
 wire n_14741;
 wire n_14742;
 wire n_14746;
 wire n_14748;
 wire n_14749;
 wire n_1475;
 wire n_14758;
 wire n_14759;
 wire n_1476;
 wire n_14760;
 wire n_14761;
 wire n_14762;
 wire n_14763;
 wire n_14764;
 wire n_14768;
 wire n_14769;
 wire n_1477;
 wire n_14770;
 wire n_14771;
 wire n_14772;
 wire n_14773;
 wire n_14774;
 wire n_1478;
 wire n_14781;
 wire n_14783;
 wire n_14784;
 wire n_14785;
 wire n_14786;
 wire n_14788;
 wire n_1479;
 wire n_14791;
 wire n_14798;
 wire n_14799;
 wire n_148;
 wire n_1480;
 wire n_14800;
 wire n_14802;
 wire n_14803;
 wire n_14804;
 wire n_14805;
 wire n_14806;
 wire n_14807;
 wire n_14808;
 wire n_14809;
 wire n_1481;
 wire n_14810;
 wire n_14811;
 wire n_14812;
 wire n_14813;
 wire n_14814;
 wire n_14815;
 wire n_14819;
 wire n_1482;
 wire n_14820;
 wire n_14822;
 wire n_14823;
 wire n_14824;
 wire n_14825;
 wire n_14826;
 wire n_14827;
 wire n_14829;
 wire n_1483;
 wire n_14831;
 wire n_14832;
 wire n_14835;
 wire n_14836;
 wire n_14837;
 wire n_14838;
 wire n_1484;
 wire n_1485;
 wire n_14857;
 wire n_1486;
 wire n_14864;
 wire n_14867;
 wire n_14868;
 wire n_1487;
 wire n_14871;
 wire n_14872;
 wire n_14873;
 wire n_14874;
 wire n_14877;
 wire n_14878;
 wire n_1488;
 wire n_14880;
 wire n_14881;
 wire n_14883;
 wire n_14887;
 wire n_1489;
 wire n_14891;
 wire n_14893;
 wire n_14894;
 wire n_14896;
 wire n_14897;
 wire n_149;
 wire n_1490;
 wire n_14902;
 wire n_14903;
 wire n_14904;
 wire n_14905;
 wire n_14906;
 wire n_14907;
 wire n_14908;
 wire n_14909;
 wire n_1491;
 wire n_14910;
 wire n_14911;
 wire n_14912;
 wire n_14914;
 wire n_14915;
 wire n_1492;
 wire n_14920;
 wire n_14921;
 wire n_14925;
 wire n_14926;
 wire n_14927;
 wire n_14928;
 wire n_14929;
 wire n_1493;
 wire n_14931;
 wire n_14932;
 wire n_14933;
 wire n_14934;
 wire n_14935;
 wire n_14936;
 wire n_14937;
 wire n_14938;
 wire n_14939;
 wire n_1494;
 wire n_14940;
 wire n_14941;
 wire n_14943;
 wire n_14944;
 wire n_14945;
 wire n_14946;
 wire n_14947;
 wire n_14948;
 wire n_14949;
 wire n_1495;
 wire n_14950;
 wire n_14951;
 wire n_1496;
 wire n_1497;
 wire n_14975;
 wire n_14977;
 wire n_14978;
 wire n_1498;
 wire n_14981;
 wire n_14984;
 wire n_14985;
 wire n_14986;
 wire n_14987;
 wire n_1499;
 wire n_14998;
 wire n_15;
 wire n_150;
 wire n_1500;
 wire n_15000;
 wire n_15001;
 wire n_15003;
 wire n_1501;
 wire n_15013;
 wire n_15014;
 wire n_1502;
 wire n_1503;
 wire n_1504;
 wire n_15045;
 wire n_15046;
 wire n_1505;
 wire n_1506;
 wire n_15060;
 wire n_15067;
 wire n_15068;
 wire n_1507;
 wire n_15070;
 wire n_15071;
 wire n_15077;
 wire n_15079;
 wire n_1508;
 wire n_15081;
 wire n_15084;
 wire n_15085;
 wire n_15086;
 wire n_15087;
 wire n_15088;
 wire n_1509;
 wire n_15090;
 wire n_15091;
 wire n_15092;
 wire n_15093;
 wire n_15094;
 wire n_15095;
 wire n_15096;
 wire n_15097;
 wire n_15098;
 wire n_151;
 wire n_1510;
 wire n_1511;
 wire n_1512;
 wire n_1513;
 wire n_1514;
 wire n_15142;
 wire n_15144;
 wire n_15145;
 wire n_15149;
 wire n_1515;
 wire n_15150;
 wire n_15151;
 wire n_15153;
 wire n_15156;
 wire n_15157;
 wire n_15158;
 wire n_1516;
 wire n_15163;
 wire n_15164;
 wire n_15166;
 wire n_15167;
 wire n_15168;
 wire n_15169;
 wire n_1517;
 wire n_15171;
 wire n_15172;
 wire n_15173;
 wire n_15174;
 wire n_15175;
 wire n_15176;
 wire n_15177;
 wire n_15178;
 wire n_15179;
 wire n_1518;
 wire n_15180;
 wire n_15181;
 wire n_15185;
 wire n_15186;
 wire n_15187;
 wire n_15188;
 wire n_1519;
 wire n_15191;
 wire n_15192;
 wire n_152;
 wire n_1520;
 wire n_15200;
 wire n_15201;
 wire n_1521;
 wire n_15210;
 wire n_15213;
 wire n_15215;
 wire n_15217;
 wire n_15218;
 wire n_1522;
 wire n_15223;
 wire n_15226;
 wire n_15227;
 wire n_1523;
 wire n_15231;
 wire n_15233;
 wire n_15235;
 wire n_15239;
 wire n_1524;
 wire n_15240;
 wire n_1525;
 wire n_1526;
 wire n_1527;
 wire n_1528;
 wire n_15289;
 wire n_1529;
 wire n_15290;
 wire n_153;
 wire n_1530;
 wire n_1531;
 wire n_1532;
 wire n_15324;
 wire n_15325;
 wire n_1533;
 wire n_15332;
 wire n_15334;
 wire n_1534;
 wire n_1535;
 wire n_15353;
 wire n_15355;
 wire n_15358;
 wire n_1536;
 wire n_15361;
 wire n_1537;
 wire n_1538;
 wire n_15380;
 wire n_15384;
 wire n_15386;
 wire n_1539;
 wire n_154;
 wire n_1540;
 wire n_1541;
 wire n_1542;
 wire n_1543;
 wire n_1544;
 wire n_15449;
 wire n_1545;
 wire n_15450;
 wire n_15451;
 wire n_15453;
 wire n_15456;
 wire n_15457;
 wire n_1546;
 wire n_15462;
 wire n_15464;
 wire n_1547;
 wire n_1548;
 wire n_1549;
 wire n_155;
 wire n_1550;
 wire n_1551;
 wire n_1552;
 wire n_1553;
 wire n_1554;
 wire n_15549;
 wire n_1555;
 wire n_15551;
 wire n_15552;
 wire n_15553;
 wire n_15559;
 wire n_1556;
 wire n_15560;
 wire n_15561;
 wire n_15567;
 wire n_15568;
 wire n_15569;
 wire n_1557;
 wire n_15570;
 wire n_15571;
 wire n_15572;
 wire n_15573;
 wire n_15574;
 wire n_15575;
 wire n_15576;
 wire n_15577;
 wire n_15578;
 wire n_15579;
 wire n_1558;
 wire n_15581;
 wire n_15584;
 wire n_15585;
 wire n_15588;
 wire n_15589;
 wire n_1559;
 wire n_15590;
 wire n_15591;
 wire n_156;
 wire n_1560;
 wire n_1561;
 wire n_1562;
 wire n_15626;
 wire n_1563;
 wire n_1564;
 wire n_15641;
 wire n_15645;
 wire n_1565;
 wire n_15651;
 wire n_1566;
 wire n_1567;
 wire n_1568;
 wire n_1569;
 wire n_157;
 wire n_1570;
 wire n_1571;
 wire n_15719;
 wire n_1572;
 wire n_15720;
 wire n_1573;
 wire n_1574;
 wire n_15740;
 wire n_1575;
 wire n_1576;
 wire n_1577;
 wire n_1578;
 wire n_1579;
 wire n_15794;
 wire n_15795;
 wire n_15796;
 wire n_15798;
 wire n_15799;
 wire n_158;
 wire n_1580;
 wire n_1581;
 wire n_15813;
 wire n_15815;
 wire n_15816;
 wire n_1582;
 wire n_1583;
 wire n_1584;
 wire n_1585;
 wire n_1586;
 wire n_1587;
 wire n_1588;
 wire n_15886;
 wire n_1589;
 wire n_159;
 wire n_1590;
 wire n_1591;
 wire n_1592;
 wire n_15920;
 wire n_15921;
 wire n_15922;
 wire n_1593;
 wire n_15939;
 wire n_1594;
 wire n_1595;
 wire n_1596;
 wire n_15960;
 wire n_15962;
 wire n_1597;
 wire n_1598;
 wire n_1599;
 wire n_15999;
 wire n_160;
 wire n_1600;
 wire n_16000;
 wire n_1601;
 wire n_1602;
 wire n_1603;
 wire n_1604;
 wire n_1605;
 wire n_16058;
 wire n_16059;
 wire n_1606;
 wire n_16060;
 wire n_16062;
 wire n_16063;
 wire n_16069;
 wire n_1607;
 wire n_16070;
 wire n_16071;
 wire n_1608;
 wire n_1609;
 wire n_161;
 wire n_1610;
 wire n_1611;
 wire n_1612;
 wire n_1613;
 wire n_1614;
 wire n_16140;
 wire n_16142;
 wire n_16149;
 wire n_1615;
 wire n_16155;
 wire n_16156;
 wire n_16158;
 wire n_1616;
 wire n_16160;
 wire n_16162;
 wire n_1617;
 wire n_1618;
 wire n_1619;
 wire n_162;
 wire n_1620;
 wire n_1621;
 wire n_1622;
 wire n_16226;
 wire n_16227;
 wire n_16228;
 wire n_1623;
 wire n_16230;
 wire n_1624;
 wire n_16247;
 wire n_1625;
 wire n_16253;
 wire n_16255;
 wire n_16256;
 wire n_16257;
 wire n_16258;
 wire n_16259;
 wire n_1626;
 wire n_1627;
 wire n_1628;
 wire n_1629;
 wire n_163;
 wire n_1630;
 wire n_1631;
 wire n_16316;
 wire n_16319;
 wire n_1632;
 wire n_16324;
 wire n_16325;
 wire n_16326;
 wire n_16327;
 wire n_1633;
 wire n_1634;
 wire n_16347;
 wire n_16348;
 wire n_16349;
 wire n_1635;
 wire n_16352;
 wire n_1636;
 wire n_16365;
 wire n_16367;
 wire n_1637;
 wire n_1638;
 wire n_1639;
 wire n_16397;
 wire n_164;
 wire n_1640;
 wire n_1641;
 wire n_16418;
 wire n_1642;
 wire n_1643;
 wire n_1644;
 wire n_1645;
 wire n_16456;
 wire n_16458;
 wire n_16459;
 wire n_1646;
 wire n_16466;
 wire n_1647;
 wire n_16475;
 wire n_16476;
 wire n_16477;
 wire n_1648;
 wire n_1649;
 wire n_165;
 wire n_1650;
 wire n_1651;
 wire n_1652;
 wire n_16528;
 wire n_16529;
 wire n_1653;
 wire n_16530;
 wire n_16532;
 wire n_16533;
 wire n_16534;
 wire n_16535;
 wire n_16536;
 wire n_1654;
 wire n_16540;
 wire n_16541;
 wire n_1655;
 wire n_16557;
 wire n_16558;
 wire n_16559;
 wire n_1656;
 wire n_16561;
 wire n_16563;
 wire n_16564;
 wire n_16565;
 wire n_1657;
 wire n_16579;
 wire n_1658;
 wire n_1659;
 wire n_16596;
 wire n_16597;
 wire n_166;
 wire n_1660;
 wire n_1661;
 wire n_16614;
 wire n_16615;
 wire n_16616;
 wire n_1662;
 wire n_1663;
 wire n_1664;
 wire n_1665;
 wire n_1666;
 wire n_16663;
 wire n_16664;
 wire n_1667;
 wire n_16676;
 wire n_1668;
 wire n_16681;
 wire n_16684;
 wire n_16685;
 wire n_1669;
 wire n_1670;
 wire n_16705;
 wire n_16706;
 wire n_16707;
 wire n_1671;
 wire n_1672;
 wire n_1673;
 wire n_1674;
 wire n_16749;
 wire n_1675;
 wire n_16751;
 wire n_16753;
 wire n_16757;
 wire n_1676;
 wire n_16763;
 wire n_16764;
 wire n_16769;
 wire n_1677;
 wire n_16772;
 wire n_16779;
 wire n_1678;
 wire n_16780;
 wire n_16781;
 wire n_16782;
 wire n_16784;
 wire n_16785;
 wire n_1679;
 wire n_168;
 wire n_1680;
 wire n_1681;
 wire n_1682;
 wire n_1683;
 wire n_1684;
 wire n_1685;
 wire n_1686;
 wire n_1687;
 wire n_1688;
 wire n_1689;
 wire n_169;
 wire n_1690;
 wire n_1691;
 wire n_1692;
 wire n_1693;
 wire n_1694;
 wire n_1695;
 wire n_1696;
 wire n_1697;
 wire n_1698;
 wire n_1699;
 wire n_17;
 wire n_170;
 wire n_1700;
 wire n_1701;
 wire n_17019;
 wire n_1702;
 wire n_17020;
 wire n_17024;
 wire n_1703;
 wire n_1704;
 wire n_1705;
 wire n_17057;
 wire n_1706;
 wire n_17063;
 wire n_17064;
 wire n_17066;
 wire n_1707;
 wire n_17072;
 wire n_17073;
 wire n_17074;
 wire n_17075;
 wire n_17076;
 wire n_17077;
 wire n_17078;
 wire n_1708;
 wire n_1709;
 wire n_1710;
 wire n_1711;
 wire n_1712;
 wire n_1713;
 wire n_1714;
 wire n_1715;
 wire n_1716;
 wire n_1717;
 wire n_1718;
 wire n_1719;
 wire n_172;
 wire n_1720;
 wire n_1721;
 wire n_1722;
 wire n_1723;
 wire n_1724;
 wire n_17240;
 wire n_17241;
 wire n_17242;
 wire n_17243;
 wire n_17244;
 wire n_17245;
 wire n_17246;
 wire n_17248;
 wire n_17249;
 wire n_1725;
 wire n_17250;
 wire n_1726;
 wire n_1727;
 wire n_1728;
 wire n_1729;
 wire n_173;
 wire n_1730;
 wire n_1731;
 wire n_1732;
 wire n_1733;
 wire n_1734;
 wire n_1735;
 wire n_1736;
 wire n_1737;
 wire n_1738;
 wire n_1739;
 wire n_17397;
 wire n_17398;
 wire n_174;
 wire n_1740;
 wire n_17400;
 wire n_17401;
 wire n_17403;
 wire n_17404;
 wire n_1741;
 wire n_17413;
 wire n_17414;
 wire n_17416;
 wire n_17417;
 wire n_17418;
 wire n_17419;
 wire n_1742;
 wire n_17420;
 wire n_1743;
 wire n_17438;
 wire n_1744;
 wire n_17440;
 wire n_17441;
 wire n_17442;
 wire n_17443;
 wire n_1745;
 wire n_1746;
 wire n_1747;
 wire n_17470;
 wire n_17471;
 wire n_17472;
 wire n_17473;
 wire n_17474;
 wire n_17475;
 wire n_1748;
 wire n_17486;
 wire n_17487;
 wire n_17488;
 wire n_17489;
 wire n_1749;
 wire n_17490;
 wire n_17491;
 wire n_17492;
 wire n_175;
 wire n_1750;
 wire n_1751;
 wire n_1752;
 wire n_1753;
 wire n_1754;
 wire n_1755;
 wire n_17551;
 wire n_17552;
 wire n_17553;
 wire n_17559;
 wire n_1756;
 wire n_17560;
 wire n_1757;
 wire n_1758;
 wire n_17587;
 wire n_1759;
 wire n_176;
 wire n_1760;
 wire n_1761;
 wire n_1762;
 wire n_1763;
 wire n_1764;
 wire n_1765;
 wire n_17651;
 wire n_17654;
 wire n_17655;
 wire n_1766;
 wire n_17661;
 wire n_17663;
 wire n_17665;
 wire n_17669;
 wire n_1767;
 wire n_17670;
 wire n_17672;
 wire n_17673;
 wire n_1768;
 wire n_1769;
 wire n_177;
 wire n_1770;
 wire n_17707;
 wire n_17709;
 wire n_1771;
 wire n_17710;
 wire n_17712;
 wire n_1772;
 wire n_1773;
 wire n_17732;
 wire n_17733;
 wire n_17734;
 wire n_17735;
 wire n_1774;
 wire n_1775;
 wire n_17754;
 wire n_1776;
 wire n_1777;
 wire n_17772;
 wire n_17773;
 wire n_17774;
 wire n_17775;
 wire n_1778;
 wire n_1779;
 wire n_178;
 wire n_1780;
 wire n_17808;
 wire n_1781;
 wire n_1782;
 wire n_17829;
 wire n_1783;
 wire n_17830;
 wire n_17831;
 wire n_17832;
 wire n_1784;
 wire n_1785;
 wire n_1786;
 wire n_17863;
 wire n_17865;
 wire n_17866;
 wire n_17867;
 wire n_17868;
 wire n_17869;
 wire n_1787;
 wire n_17870;
 wire n_17871;
 wire n_17872;
 wire n_17873;
 wire n_17874;
 wire n_17875;
 wire n_17876;
 wire n_17877;
 wire n_17878;
 wire n_17879;
 wire n_1788;
 wire n_17880;
 wire n_17882;
 wire n_17883;
 wire n_17884;
 wire n_17885;
 wire n_17886;
 wire n_1789;
 wire n_179;
 wire n_1790;
 wire n_17907;
 wire n_17908;
 wire n_17909;
 wire n_1791;
 wire n_17910;
 wire n_1792;
 wire n_1793;
 wire n_17936;
 wire n_17938;
 wire n_17939;
 wire n_1794;
 wire n_17940;
 wire n_1795;
 wire n_1796;
 wire n_1797;
 wire n_17976;
 wire n_17977;
 wire n_17978;
 wire n_17979;
 wire n_1798;
 wire n_1799;
 wire n_17997;
 wire n_17998;
 wire n_18;
 wire n_1800;
 wire n_18002;
 wire n_18003;
 wire n_18004;
 wire n_18008;
 wire n_18009;
 wire n_1801;
 wire n_1802;
 wire n_1803;
 wire n_18031;
 wire n_18034;
 wire n_18039;
 wire n_1804;
 wire n_18041;
 wire n_18049;
 wire n_1805;
 wire n_18050;
 wire n_1806;
 wire n_18063;
 wire n_18064;
 wire n_18065;
 wire n_18067;
 wire n_18068;
 wire n_18069;
 wire n_1807;
 wire n_1808;
 wire n_18084;
 wire n_18085;
 wire n_1809;
 wire n_18091;
 wire n_18092;
 wire n_18093;
 wire n_18094;
 wire n_181;
 wire n_1810;
 wire n_1811;
 wire n_1812;
 wire n_18124;
 wire n_1813;
 wire n_1814;
 wire n_18141;
 wire n_18144;
 wire n_1815;
 wire n_18154;
 wire n_18155;
 wire n_18157;
 wire n_1816;
 wire n_18165;
 wire n_18166;
 wire n_18167;
 wire n_18168;
 wire n_1817;
 wire n_18175;
 wire n_1818;
 wire n_1819;
 wire n_182;
 wire n_1820;
 wire n_1821;
 wire n_1822;
 wire n_1823;
 wire n_1824;
 wire n_1825;
 wire n_1826;
 wire n_1827;
 wire n_1828;
 wire n_1829;
 wire n_183;
 wire n_1830;
 wire n_1831;
 wire n_1832;
 wire n_1833;
 wire n_1834;
 wire n_1835;
 wire n_1836;
 wire n_1837;
 wire n_1838;
 wire n_1839;
 wire n_184;
 wire n_1840;
 wire n_1841;
 wire n_1842;
 wire n_1843;
 wire n_18430;
 wire n_18431;
 wire n_18432;
 wire n_1844;
 wire n_1845;
 wire n_18458;
 wire n_1846;
 wire n_1847;
 wire n_1848;
 wire n_1849;
 wire n_185;
 wire n_1850;
 wire n_1851;
 wire n_1852;
 wire n_1853;
 wire n_1854;
 wire n_1855;
 wire n_1856;
 wire n_1857;
 wire n_18577;
 wire n_18578;
 wire n_18579;
 wire n_1858;
 wire n_18580;
 wire n_18581;
 wire n_18582;
 wire n_1859;
 wire n_18597;
 wire n_186;
 wire n_1860;
 wire n_18605;
 wire n_1861;
 wire n_1862;
 wire n_1863;
 wire n_1864;
 wire n_18648;
 wire n_1865;
 wire n_1866;
 wire n_18663;
 wire n_18664;
 wire n_18665;
 wire n_18666;
 wire n_18667;
 wire n_1867;
 wire n_1868;
 wire n_1869;
 wire n_18692;
 wire n_18695;
 wire n_18698;
 wire n_18699;
 wire n_187;
 wire n_1870;
 wire n_18700;
 wire n_18701;
 wire n_18702;
 wire n_18703;
 wire n_18704;
 wire n_18707;
 wire n_1871;
 wire n_18710;
 wire n_18711;
 wire n_18712;
 wire n_18716;
 wire n_18717;
 wire n_18718;
 wire n_18719;
 wire n_1872;
 wire n_18720;
 wire n_18721;
 wire n_18726;
 wire n_18729;
 wire n_1873;
 wire n_18730;
 wire n_18731;
 wire n_18732;
 wire n_18737;
 wire n_18738;
 wire n_18739;
 wire n_1874;
 wire n_18740;
 wire n_18748;
 wire n_18749;
 wire n_1875;
 wire n_18751;
 wire n_18752;
 wire n_18753;
 wire n_18754;
 wire n_18756;
 wire n_18757;
 wire n_18758;
 wire n_1876;
 wire n_18760;
 wire n_18761;
 wire n_18763;
 wire n_18764;
 wire n_18765;
 wire n_18766;
 wire n_18767;
 wire n_18769;
 wire n_1877;
 wire n_18770;
 wire n_18771;
 wire n_18774;
 wire n_18775;
 wire n_18776;
 wire n_18778;
 wire n_18779;
 wire n_1878;
 wire n_18780;
 wire n_18781;
 wire n_18782;
 wire n_18783;
 wire n_18785;
 wire n_18786;
 wire n_18787;
 wire n_1879;
 wire n_18790;
 wire n_18791;
 wire n_18793;
 wire n_18794;
 wire n_18795;
 wire n_18797;
 wire n_18798;
 wire n_18799;
 wire n_188;
 wire n_1880;
 wire n_18800;
 wire n_18802;
 wire n_18803;
 wire n_18804;
 wire n_18806;
 wire n_18807;
 wire n_18809;
 wire n_1881;
 wire n_18811;
 wire n_18812;
 wire n_18815;
 wire n_18819;
 wire n_1882;
 wire n_18820;
 wire n_18822;
 wire n_18823;
 wire n_18825;
 wire n_18826;
 wire n_18827;
 wire n_18828;
 wire n_1883;
 wire n_18831;
 wire n_18832;
 wire n_18835;
 wire n_18836;
 wire n_18838;
 wire n_18839;
 wire n_1884;
 wire n_18842;
 wire n_18843;
 wire n_18846;
 wire n_18848;
 wire n_18849;
 wire n_1885;
 wire n_18850;
 wire n_18851;
 wire n_18856;
 wire n_18857;
 wire n_18858;
 wire n_1886;
 wire n_18862;
 wire n_18863;
 wire n_18865;
 wire n_18866;
 wire n_18867;
 wire n_18868;
 wire n_1887;
 wire n_18870;
 wire n_18871;
 wire n_18874;
 wire n_18875;
 wire n_1888;
 wire n_18881;
 wire n_18883;
 wire n_18884;
 wire n_18885;
 wire n_18886;
 wire n_18889;
 wire n_1889;
 wire n_18891;
 wire n_18896;
 wire n_18897;
 wire n_18899;
 wire n_189;
 wire n_1890;
 wire n_18900;
 wire n_18901;
 wire n_18902;
 wire n_18903;
 wire n_18904;
 wire n_18907;
 wire n_1891;
 wire n_18914;
 wire n_18915;
 wire n_18916;
 wire n_18919;
 wire n_1892;
 wire n_18925;
 wire n_18926;
 wire n_18927;
 wire n_18928;
 wire n_18929;
 wire n_1893;
 wire n_18930;
 wire n_18933;
 wire n_18934;
 wire n_18935;
 wire n_18938;
 wire n_18939;
 wire n_1894;
 wire n_18940;
 wire n_18941;
 wire n_18942;
 wire n_18943;
 wire n_18945;
 wire n_18947;
 wire n_18948;
 wire n_18949;
 wire n_1895;
 wire n_18952;
 wire n_18953;
 wire n_18954;
 wire n_18956;
 wire n_18957;
 wire n_1896;
 wire n_18960;
 wire n_18961;
 wire n_18964;
 wire n_18967;
 wire n_18968;
 wire n_18969;
 wire n_1897;
 wire n_18970;
 wire n_18972;
 wire n_18973;
 wire n_18974;
 wire n_18978;
 wire n_1898;
 wire n_18983;
 wire n_18985;
 wire n_18986;
 wire n_18987;
 wire n_18988;
 wire n_1899;
 wire n_18992;
 wire n_18993;
 wire n_18996;
 wire n_18997;
 wire n_18999;
 wire n_19;
 wire n_190;
 wire n_1900;
 wire n_19001;
 wire n_19002;
 wire n_19006;
 wire n_19007;
 wire n_19008;
 wire n_1901;
 wire n_19011;
 wire n_19012;
 wire n_19013;
 wire n_19014;
 wire n_19015;
 wire n_19016;
 wire n_19017;
 wire n_19018;
 wire n_19019;
 wire n_1902;
 wire n_19020;
 wire n_19021;
 wire n_19022;
 wire n_19023;
 wire n_19024;
 wire n_19027;
 wire n_19028;
 wire n_19029;
 wire n_1903;
 wire n_19032;
 wire n_19033;
 wire n_19034;
 wire n_19035;
 wire n_19036;
 wire n_19037;
 wire n_19038;
 wire n_19039;
 wire n_1904;
 wire n_19041;
 wire n_19043;
 wire n_19044;
 wire n_19045;
 wire n_19049;
 wire n_1905;
 wire n_19050;
 wire n_19052;
 wire n_19053;
 wire n_19054;
 wire n_19055;
 wire n_19056;
 wire n_19057;
 wire n_19058;
 wire n_19059;
 wire n_1906;
 wire n_19060;
 wire n_19061;
 wire n_19062;
 wire n_19063;
 wire n_19064;
 wire n_19065;
 wire n_19067;
 wire n_19068;
 wire n_19069;
 wire n_1907;
 wire n_19070;
 wire n_19071;
 wire n_19072;
 wire n_19073;
 wire n_19075;
 wire n_19076;
 wire n_19077;
 wire n_19078;
 wire n_19079;
 wire n_1908;
 wire n_19080;
 wire n_19083;
 wire n_19084;
 wire n_19085;
 wire n_19086;
 wire n_19088;
 wire n_19089;
 wire n_1909;
 wire n_19090;
 wire n_19091;
 wire n_19093;
 wire n_19095;
 wire n_19096;
 wire n_19097;
 wire n_19098;
 wire n_19099;
 wire n_191;
 wire n_1910;
 wire n_19101;
 wire n_19102;
 wire n_19103;
 wire n_19104;
 wire n_19105;
 wire n_19106;
 wire n_19108;
 wire n_19109;
 wire n_1911;
 wire n_19111;
 wire n_19112;
 wire n_19113;
 wire n_19114;
 wire n_19115;
 wire n_19117;
 wire n_1912;
 wire n_19120;
 wire n_19122;
 wire n_19123;
 wire n_19124;
 wire n_19126;
 wire n_19128;
 wire n_19129;
 wire n_1913;
 wire n_19131;
 wire n_19132;
 wire n_19133;
 wire n_19134;
 wire n_19135;
 wire n_19136;
 wire n_19137;
 wire n_19138;
 wire n_1914;
 wire n_19141;
 wire n_19142;
 wire n_19143;
 wire n_19144;
 wire n_19145;
 wire n_19146;
 wire n_19147;
 wire n_19149;
 wire n_1915;
 wire n_19150;
 wire n_1916;
 wire n_19160;
 wire n_19164;
 wire n_19165;
 wire n_19168;
 wire n_19169;
 wire n_1917;
 wire n_19170;
 wire n_19172;
 wire n_19174;
 wire n_19175;
 wire n_19177;
 wire n_1918;
 wire n_19181;
 wire n_19182;
 wire n_19183;
 wire n_19185;
 wire n_19186;
 wire n_19187;
 wire n_19188;
 wire n_19189;
 wire n_1919;
 wire n_19190;
 wire n_19191;
 wire n_19193;
 wire n_19194;
 wire n_19195;
 wire n_19197;
 wire n_19199;
 wire n_192;
 wire n_1920;
 wire n_19200;
 wire n_19201;
 wire n_19205;
 wire n_19206;
 wire n_19207;
 wire n_19208;
 wire n_1921;
 wire n_19218;
 wire n_19219;
 wire n_1922;
 wire n_19222;
 wire n_19228;
 wire n_1923;
 wire n_19230;
 wire n_19232;
 wire n_19234;
 wire n_19235;
 wire n_19236;
 wire n_19237;
 wire n_1924;
 wire n_19240;
 wire n_19241;
 wire n_19242;
 wire n_19243;
 wire n_19248;
 wire n_19249;
 wire n_1925;
 wire n_19252;
 wire n_19253;
 wire n_19254;
 wire n_19259;
 wire n_1926;
 wire n_19261;
 wire n_19263;
 wire n_19264;
 wire n_19265;
 wire n_19267;
 wire n_19268;
 wire n_19269;
 wire n_1927;
 wire n_19270;
 wire n_19271;
 wire n_19272;
 wire n_19273;
 wire n_19274;
 wire n_19275;
 wire n_19276;
 wire n_19277;
 wire n_19278;
 wire n_19279;
 wire n_1928;
 wire n_19280;
 wire n_19281;
 wire n_19282;
 wire n_19283;
 wire n_19288;
 wire n_19289;
 wire n_1929;
 wire n_19290;
 wire n_19291;
 wire n_193;
 wire n_1930;
 wire n_19304;
 wire n_19305;
 wire n_19306;
 wire n_19307;
 wire n_19308;
 wire n_19309;
 wire n_1931;
 wire n_19310;
 wire n_19314;
 wire n_19316;
 wire n_1932;
 wire n_19323;
 wire n_19324;
 wire n_19325;
 wire n_19326;
 wire n_19327;
 wire n_1933;
 wire n_19330;
 wire n_19331;
 wire n_19332;
 wire n_19333;
 wire n_19334;
 wire n_19335;
 wire n_19336;
 wire n_19337;
 wire n_19338;
 wire n_19339;
 wire n_1934;
 wire n_19340;
 wire n_19341;
 wire n_19342;
 wire n_1935;
 wire n_19353;
 wire n_19354;
 wire n_19355;
 wire n_19356;
 wire n_19357;
 wire n_19358;
 wire n_19359;
 wire n_1936;
 wire n_19360;
 wire n_19363;
 wire n_19365;
 wire n_19366;
 wire n_19367;
 wire n_19368;
 wire n_19369;
 wire n_1937;
 wire n_19370;
 wire n_19371;
 wire n_19372;
 wire n_19374;
 wire n_19375;
 wire n_19376;
 wire n_19377;
 wire n_19378;
 wire n_1938;
 wire n_19380;
 wire n_19381;
 wire n_19382;
 wire n_19385;
 wire n_19386;
 wire n_19387;
 wire n_1939;
 wire n_19390;
 wire n_19391;
 wire n_19393;
 wire n_19394;
 wire n_19395;
 wire n_19396;
 wire n_19398;
 wire n_194;
 wire n_1940;
 wire n_19400;
 wire n_19404;
 wire n_19407;
 wire n_19408;
 wire n_1941;
 wire n_19410;
 wire n_19411;
 wire n_1942;
 wire n_19428;
 wire n_19429;
 wire n_1943;
 wire n_19430;
 wire n_19431;
 wire n_19432;
 wire n_19433;
 wire n_19435;
 wire n_19436;
 wire n_19437;
 wire n_19438;
 wire n_19439;
 wire n_1944;
 wire n_19440;
 wire n_19441;
 wire n_19442;
 wire n_19443;
 wire n_19444;
 wire n_19445;
 wire n_19446;
 wire n_19447;
 wire n_19448;
 wire n_19449;
 wire n_1945;
 wire n_19453;
 wire n_19454;
 wire n_19457;
 wire n_1946;
 wire n_19461;
 wire n_19462;
 wire n_1947;
 wire n_19471;
 wire n_19472;
 wire n_19478;
 wire n_1948;
 wire n_19480;
 wire n_19484;
 wire n_19485;
 wire n_19486;
 wire n_19487;
 wire n_19488;
 wire n_19489;
 wire n_1949;
 wire n_19490;
 wire n_19491;
 wire n_19492;
 wire n_19493;
 wire n_19494;
 wire n_19495;
 wire n_19496;
 wire n_19497;
 wire n_19498;
 wire n_19499;
 wire n_195;
 wire n_1950;
 wire n_19500;
 wire n_19501;
 wire n_19502;
 wire n_19503;
 wire n_19504;
 wire n_19505;
 wire n_1951;
 wire n_19515;
 wire n_19516;
 wire n_19517;
 wire n_1952;
 wire n_19522;
 wire n_19523;
 wire n_19525;
 wire n_1953;
 wire n_19530;
 wire n_19531;
 wire n_19532;
 wire n_19533;
 wire n_19534;
 wire n_19538;
 wire n_19539;
 wire n_1954;
 wire n_19540;
 wire n_19541;
 wire n_19542;
 wire n_19543;
 wire n_1955;
 wire n_19550;
 wire n_19551;
 wire n_19552;
 wire n_19553;
 wire n_19554;
 wire n_19555;
 wire n_19556;
 wire n_19557;
 wire n_19558;
 wire n_19559;
 wire n_1956;
 wire n_19563;
 wire n_19564;
 wire n_19565;
 wire n_19566;
 wire n_19567;
 wire n_19568;
 wire n_1957;
 wire n_19570;
 wire n_19571;
 wire n_19572;
 wire n_19573;
 wire n_19575;
 wire n_1958;
 wire n_19582;
 wire n_19583;
 wire n_19584;
 wire n_1959;
 wire n_19594;
 wire n_19595;
 wire n_19597;
 wire n_19598;
 wire n_19599;
 wire n_196;
 wire n_1960;
 wire n_19600;
 wire n_19601;
 wire n_19602;
 wire n_19604;
 wire n_19605;
 wire n_19607;
 wire n_1961;
 wire n_19612;
 wire n_19613;
 wire n_19614;
 wire n_19615;
 wire n_1962;
 wire n_19621;
 wire n_19622;
 wire n_19623;
 wire n_19625;
 wire n_1963;
 wire n_1964;
 wire n_19644;
 wire n_19645;
 wire n_19646;
 wire n_19647;
 wire n_19648;
 wire n_19649;
 wire n_1965;
 wire n_19650;
 wire n_19656;
 wire n_19657;
 wire n_19658;
 wire n_1966;
 wire n_19660;
 wire n_19661;
 wire n_19662;
 wire n_19663;
 wire n_19664;
 wire n_19665;
 wire n_19666;
 wire n_19667;
 wire n_19669;
 wire n_1967;
 wire n_19670;
 wire n_19672;
 wire n_19673;
 wire n_19674;
 wire n_19675;
 wire n_19676;
 wire n_19677;
 wire n_19679;
 wire n_1968;
 wire n_19680;
 wire n_19681;
 wire n_19682;
 wire n_19685;
 wire n_19686;
 wire n_19688;
 wire n_1969;
 wire n_19695;
 wire n_19696;
 wire n_19697;
 wire n_19698;
 wire n_19699;
 wire n_1970;
 wire n_19700;
 wire n_19701;
 wire n_19702;
 wire n_19703;
 wire n_19704;
 wire n_19705;
 wire n_19706;
 wire n_1971;
 wire n_19710;
 wire n_19711;
 wire n_19712;
 wire n_19714;
 wire n_19718;
 wire n_19719;
 wire n_1972;
 wire n_19722;
 wire n_19729;
 wire n_1973;
 wire n_19730;
 wire n_19732;
 wire n_19734;
 wire n_19736;
 wire n_19737;
 wire n_1974;
 wire n_19746;
 wire n_1975;
 wire n_19752;
 wire n_19753;
 wire n_19754;
 wire n_1976;
 wire n_19764;
 wire n_19767;
 wire n_19768;
 wire n_19769;
 wire n_1977;
 wire n_19773;
 wire n_19774;
 wire n_19775;
 wire n_19776;
 wire n_19777;
 wire n_19778;
 wire n_19779;
 wire n_1978;
 wire n_19783;
 wire n_19785;
 wire n_19787;
 wire n_19789;
 wire n_1979;
 wire n_19790;
 wire n_19792;
 wire n_19795;
 wire n_19796;
 wire n_19797;
 wire n_19799;
 wire n_198;
 wire n_1980;
 wire n_19800;
 wire n_19801;
 wire n_19802;
 wire n_19803;
 wire n_19804;
 wire n_19808;
 wire n_19809;
 wire n_1981;
 wire n_19810;
 wire n_19814;
 wire n_19815;
 wire n_19816;
 wire n_1982;
 wire n_19820;
 wire n_19821;
 wire n_19825;
 wire n_19826;
 wire n_19827;
 wire n_19829;
 wire n_1983;
 wire n_19830;
 wire n_19831;
 wire n_19832;
 wire n_19833;
 wire n_19834;
 wire n_19835;
 wire n_19838;
 wire n_1984;
 wire n_19840;
 wire n_19844;
 wire n_1985;
 wire n_19850;
 wire n_19851;
 wire n_19855;
 wire n_19856;
 wire n_19857;
 wire n_19858;
 wire n_19859;
 wire n_1986;
 wire n_19860;
 wire n_19861;
 wire n_19862;
 wire n_19863;
 wire n_19864;
 wire n_19865;
 wire n_19866;
 wire n_19867;
 wire n_19868;
 wire n_19869;
 wire n_1987;
 wire n_19877;
 wire n_19878;
 wire n_1988;
 wire n_19882;
 wire n_19884;
 wire n_19886;
 wire n_1989;
 wire n_19890;
 wire n_19892;
 wire n_19893;
 wire n_19894;
 wire n_19898;
 wire n_19899;
 wire n_199;
 wire n_1990;
 wire n_19900;
 wire n_19901;
 wire n_19903;
 wire n_19904;
 wire n_19905;
 wire n_19907;
 wire n_19908;
 wire n_19909;
 wire n_1991;
 wire n_19910;
 wire n_19911;
 wire n_19912;
 wire n_19913;
 wire n_19914;
 wire n_19915;
 wire n_19917;
 wire n_19918;
 wire n_1992;
 wire n_19928;
 wire n_19929;
 wire n_1993;
 wire n_19930;
 wire n_1994;
 wire n_19945;
 wire n_19948;
 wire n_19949;
 wire n_1995;
 wire n_19950;
 wire n_19951;
 wire n_19952;
 wire n_19953;
 wire n_19954;
 wire n_19955;
 wire n_19956;
 wire n_19957;
 wire n_19958;
 wire n_19959;
 wire n_1996;
 wire n_19963;
 wire n_19964;
 wire n_19965;
 wire n_19967;
 wire n_19969;
 wire n_1997;
 wire n_19970;
 wire n_19971;
 wire n_1998;
 wire n_19981;
 wire n_19982;
 wire n_19983;
 wire n_19985;
 wire n_19989;
 wire n_1999;
 wire n_200;
 wire n_2000;
 wire n_20006;
 wire n_20008;
 wire n_2001;
 wire n_20012;
 wire n_20013;
 wire n_20016;
 wire n_20017;
 wire n_20018;
 wire n_2002;
 wire n_20022;
 wire n_20023;
 wire n_20025;
 wire n_20026;
 wire n_20027;
 wire n_20028;
 wire n_20029;
 wire n_2003;
 wire n_20030;
 wire n_20034;
 wire n_20035;
 wire n_20036;
 wire n_20037;
 wire n_20038;
 wire n_20039;
 wire n_2004;
 wire n_20040;
 wire n_20041;
 wire n_20043;
 wire n_20044;
 wire n_20045;
 wire n_20046;
 wire n_20047;
 wire n_2005;
 wire n_20054;
 wire n_2006;
 wire n_20066;
 wire n_2007;
 wire n_20071;
 wire n_20072;
 wire n_20073;
 wire n_20074;
 wire n_20075;
 wire n_20076;
 wire n_20077;
 wire n_20078;
 wire n_2008;
 wire n_20082;
 wire n_20083;
 wire n_20087;
 wire n_20088;
 wire n_2009;
 wire n_20093;
 wire n_20094;
 wire n_20095;
 wire n_20096;
 wire n_20097;
 wire n_20098;
 wire n_20099;
 wire n_201;
 wire n_2010;
 wire n_20101;
 wire n_20103;
 wire n_20106;
 wire n_20107;
 wire n_20108;
 wire n_20109;
 wire n_2011;
 wire n_20110;
 wire n_20111;
 wire n_20112;
 wire n_20113;
 wire n_20114;
 wire n_20115;
 wire n_20116;
 wire n_20117;
 wire n_20118;
 wire n_2012;
 wire n_20120;
 wire n_20121;
 wire n_20122;
 wire n_20123;
 wire n_20124;
 wire n_20125;
 wire n_20126;
 wire n_20127;
 wire n_20128;
 wire n_20129;
 wire n_2013;
 wire n_20130;
 wire n_20131;
 wire n_20132;
 wire n_20133;
 wire n_20134;
 wire n_20135;
 wire n_20136;
 wire n_20137;
 wire n_20138;
 wire n_20139;
 wire n_2014;
 wire n_20140;
 wire n_20141;
 wire n_20142;
 wire n_20143;
 wire n_20148;
 wire n_20149;
 wire n_2015;
 wire n_20151;
 wire n_20152;
 wire n_20156;
 wire n_20157;
 wire n_20158;
 wire n_2016;
 wire n_20160;
 wire n_20161;
 wire n_20162;
 wire n_20163;
 wire n_20164;
 wire n_2017;
 wire n_2018;
 wire n_2019;
 wire n_20195;
 wire n_20198;
 wire n_20199;
 wire n_202;
 wire n_2020;
 wire n_20200;
 wire n_2021;
 wire n_20210;
 wire n_20214;
 wire n_20215;
 wire n_20216;
 wire n_20217;
 wire n_20218;
 wire n_20219;
 wire n_2022;
 wire n_20220;
 wire n_20221;
 wire n_20222;
 wire n_20223;
 wire n_2023;
 wire n_20231;
 wire n_20232;
 wire n_20233;
 wire n_20234;
 wire n_20235;
 wire n_20236;
 wire n_20237;
 wire n_20238;
 wire n_20239;
 wire n_2024;
 wire n_20248;
 wire n_2025;
 wire n_2026;
 wire n_2027;
 wire n_20274;
 wire n_20275;
 wire n_20276;
 wire n_20277;
 wire n_20279;
 wire n_2028;
 wire n_20280;
 wire n_20281;
 wire n_20282;
 wire n_20283;
 wire n_20285;
 wire n_20287;
 wire n_20288;
 wire n_2029;
 wire n_20290;
 wire n_20291;
 wire n_20292;
 wire n_20293;
 wire n_20294;
 wire n_20295;
 wire n_20296;
 wire n_20297;
 wire n_203;
 wire n_2030;
 wire n_20301;
 wire n_20302;
 wire n_20303;
 wire n_20304;
 wire n_20305;
 wire n_20306;
 wire n_20307;
 wire n_20309;
 wire n_2031;
 wire n_20310;
 wire n_20311;
 wire n_20312;
 wire n_20313;
 wire n_20314;
 wire n_2032;
 wire n_20321;
 wire n_20322;
 wire n_20324;
 wire n_20326;
 wire n_20327;
 wire n_20328;
 wire n_20329;
 wire n_20330;
 wire n_20331;
 wire n_20332;
 wire n_20333;
 wire n_20334;
 wire n_20335;
 wire n_20336;
 wire n_20343;
 wire n_20344;
 wire n_20345;
 wire n_20346;
 wire n_20347;
 wire n_20353;
 wire n_20354;
 wire n_20355;
 wire n_20356;
 wire n_20357;
 wire n_20358;
 wire n_20359;
 wire n_20360;
 wire n_20361;
 wire n_20362;
 wire n_20363;
 wire n_20365;
 wire n_20369;
 wire n_2037;
 wire n_20370;
 wire n_20371;
 wire n_20372;
 wire n_20373;
 wire n_20374;
 wire n_20375;
 wire n_20376;
 wire n_20377;
 wire n_20379;
 wire n_2038;
 wire n_20380;
 wire n_20383;
 wire n_20384;
 wire n_20385;
 wire n_2039;
 wire n_20390;
 wire n_20393;
 wire n_20395;
 wire n_20396;
 wire n_20397;
 wire n_20398;
 wire n_20399;
 wire n_2040;
 wire n_20400;
 wire n_20401;
 wire n_20405;
 wire n_2041;
 wire n_20413;
 wire n_2042;
 wire n_20421;
 wire n_20422;
 wire n_2043;
 wire n_2044;
 wire n_2045;
 wire n_20459;
 wire n_2046;
 wire n_20463;
 wire n_20464;
 wire n_2047;
 wire n_20478;
 wire n_2048;
 wire n_20480;
 wire n_20481;
 wire n_20488;
 wire n_2049;
 wire n_20494;
 wire n_20496;
 wire n_205;
 wire n_2050;
 wire n_20500;
 wire n_20501;
 wire n_20503;
 wire n_20504;
 wire n_2051;
 wire n_20510;
 wire n_20512;
 wire n_20514;
 wire n_20519;
 wire n_2052;
 wire n_20520;
 wire n_2053;
 wire n_2054;
 wire n_2055;
 wire n_2056;
 wire n_2057;
 wire n_2058;
 wire n_20588;
 wire n_20589;
 wire n_2059;
 wire n_20590;
 wire n_20591;
 wire n_206;
 wire n_2060;
 wire n_2061;
 wire n_2062;
 wire n_20621;
 wire n_20623;
 wire n_20624;
 wire n_20625;
 wire n_20629;
 wire n_2063;
 wire n_20630;
 wire n_20633;
 wire n_20637;
 wire n_20638;
 wire n_20639;
 wire n_2064;
 wire n_20640;
 wire n_20641;
 wire n_20642;
 wire n_20643;
 wire n_20644;
 wire n_20645;
 wire n_20646;
 wire n_20649;
 wire n_2065;
 wire n_20650;
 wire n_20651;
 wire n_20652;
 wire n_20653;
 wire n_20654;
 wire n_20656;
 wire n_20659;
 wire n_2066;
 wire n_20660;
 wire n_2067;
 wire n_20670;
 wire n_20671;
 wire n_20673;
 wire n_20674;
 wire n_20675;
 wire n_2068;
 wire n_20680;
 wire n_20681;
 wire n_20682;
 wire n_20683;
 wire n_20684;
 wire n_20687;
 wire n_20688;
 wire n_20689;
 wire n_2069;
 wire n_20696;
 wire n_207;
 wire n_2070;
 wire n_20700;
 wire n_2071;
 wire n_20716;
 wire n_20717;
 wire n_20718;
 wire n_20719;
 wire n_2072;
 wire n_20720;
 wire n_20721;
 wire n_20723;
 wire n_20724;
 wire n_20725;
 wire n_20726;
 wire n_20727;
 wire n_20728;
 wire n_20729;
 wire n_2073;
 wire n_20730;
 wire n_20731;
 wire n_20737;
 wire n_20738;
 wire n_20739;
 wire n_2074;
 wire n_20740;
 wire n_20741;
 wire n_20742;
 wire n_2075;
 wire n_20752;
 wire n_20758;
 wire n_20759;
 wire n_2076;
 wire n_20764;
 wire n_20765;
 wire n_20767;
 wire n_20769;
 wire n_2077;
 wire n_20770;
 wire n_20771;
 wire n_20773;
 wire n_20776;
 wire n_20777;
 wire n_20778;
 wire n_2078;
 wire n_20782;
 wire n_20783;
 wire n_20784;
 wire n_20785;
 wire n_20786;
 wire n_20787;
 wire n_20788;
 wire n_20789;
 wire n_2079;
 wire n_20793;
 wire n_20794;
 wire n_20795;
 wire n_20796;
 wire n_208;
 wire n_2080;
 wire n_20809;
 wire n_2081;
 wire n_20810;
 wire n_20811;
 wire n_20812;
 wire n_20813;
 wire n_20814;
 wire n_2082;
 wire n_20823;
 wire n_20824;
 wire n_20825;
 wire n_20828;
 wire n_20829;
 wire n_2083;
 wire n_20830;
 wire n_20831;
 wire n_20832;
 wire n_20833;
 wire n_2084;
 wire n_20841;
 wire n_20842;
 wire n_20843;
 wire n_20844;
 wire n_20845;
 wire n_20847;
 wire n_20849;
 wire n_2085;
 wire n_20850;
 wire n_20851;
 wire n_20852;
 wire n_20853;
 wire n_20855;
 wire n_20856;
 wire n_20857;
 wire n_20859;
 wire n_2086;
 wire n_20860;
 wire n_20861;
 wire n_20862;
 wire n_20863;
 wire n_20864;
 wire n_20865;
 wire n_20866;
 wire n_20867;
 wire n_20868;
 wire n_20869;
 wire n_2087;
 wire n_20870;
 wire n_20871;
 wire n_20872;
 wire n_20873;
 wire n_20874;
 wire n_20875;
 wire n_20876;
 wire n_20877;
 wire n_20878;
 wire n_2088;
 wire n_20881;
 wire n_20882;
 wire n_20883;
 wire n_20884;
 wire n_20885;
 wire n_20886;
 wire n_20887;
 wire n_20888;
 wire n_2089;
 wire n_20893;
 wire n_20894;
 wire n_20895;
 wire n_20896;
 wire n_20897;
 wire n_20898;
 wire n_20899;
 wire n_209;
 wire n_2090;
 wire n_20900;
 wire n_20901;
 wire n_20902;
 wire n_20903;
 wire n_20904;
 wire n_20905;
 wire n_20909;
 wire n_2091;
 wire n_20911;
 wire n_20912;
 wire n_20913;
 wire n_20914;
 wire n_20916;
 wire n_20917;
 wire n_2092;
 wire n_20921;
 wire n_20922;
 wire n_20923;
 wire n_20924;
 wire n_20925;
 wire n_20926;
 wire n_20927;
 wire n_20928;
 wire n_2093;
 wire n_20931;
 wire n_20932;
 wire n_20933;
 wire n_20934;
 wire n_20935;
 wire n_20936;
 wire n_20938;
 wire n_20939;
 wire n_2094;
 wire n_20943;
 wire n_20945;
 wire n_20946;
 wire n_20949;
 wire n_2095;
 wire n_20950;
 wire n_20951;
 wire n_20953;
 wire n_20954;
 wire n_20956;
 wire n_20957;
 wire n_20959;
 wire n_2096;
 wire n_20961;
 wire n_20963;
 wire n_20964;
 wire n_20965;
 wire n_20966;
 wire n_20967;
 wire n_20968;
 wire n_20969;
 wire n_2097;
 wire n_20971;
 wire n_20972;
 wire n_20973;
 wire n_20974;
 wire n_20975;
 wire n_20976;
 wire n_20977;
 wire n_20979;
 wire n_2098;
 wire n_20981;
 wire n_20982;
 wire n_20983;
 wire n_20984;
 wire n_20985;
 wire n_20986;
 wire n_20987;
 wire n_20988;
 wire n_20989;
 wire n_2099;
 wire n_20990;
 wire n_20993;
 wire n_20994;
 wire n_20996;
 wire n_20997;
 wire n_20998;
 wire n_20999;
 wire n_21;
 wire n_210;
 wire n_2100;
 wire n_21000;
 wire n_21002;
 wire n_21004;
 wire n_21007;
 wire n_2101;
 wire n_21010;
 wire n_21013;
 wire n_21014;
 wire n_21015;
 wire n_21016;
 wire n_2102;
 wire n_21020;
 wire n_21023;
 wire n_21025;
 wire n_21026;
 wire n_21028;
 wire n_2103;
 wire n_21036;
 wire n_21038;
 wire n_2104;
 wire n_21042;
 wire n_21043;
 wire n_21044;
 wire n_21045;
 wire n_21046;
 wire n_21047;
 wire n_21048;
 wire n_21049;
 wire n_2105;
 wire n_21050;
 wire n_21051;
 wire n_21052;
 wire n_21056;
 wire n_21058;
 wire n_21059;
 wire n_2106;
 wire n_21061;
 wire n_21062;
 wire n_21064;
 wire n_21065;
 wire n_21066;
 wire n_21067;
 wire n_21069;
 wire n_2107;
 wire n_21071;
 wire n_21072;
 wire n_21073;
 wire n_21074;
 wire n_21075;
 wire n_21077;
 wire n_21078;
 wire n_21079;
 wire n_2108;
 wire n_21080;
 wire n_21081;
 wire n_21082;
 wire n_21083;
 wire n_21084;
 wire n_2109;
 wire n_21091;
 wire n_21092;
 wire n_21093;
 wire n_21097;
 wire n_21098;
 wire n_211;
 wire n_2110;
 wire n_2111;
 wire n_21110;
 wire n_21111;
 wire n_21112;
 wire n_21113;
 wire n_21117;
 wire n_21118;
 wire n_2112;
 wire n_21126;
 wire n_21129;
 wire n_2113;
 wire n_21130;
 wire n_21131;
 wire n_21134;
 wire n_21135;
 wire n_21136;
 wire n_21137;
 wire n_21139;
 wire n_2114;
 wire n_21140;
 wire n_21141;
 wire n_21142;
 wire n_21143;
 wire n_21144;
 wire n_21146;
 wire n_21147;
 wire n_21148;
 wire n_2115;
 wire n_21151;
 wire n_21152;
 wire n_21157;
 wire n_21159;
 wire n_2116;
 wire n_21160;
 wire n_21161;
 wire n_21162;
 wire n_21163;
 wire n_21164;
 wire n_21165;
 wire n_21166;
 wire n_21167;
 wire n_21168;
 wire n_21169;
 wire n_2117;
 wire n_21170;
 wire n_21177;
 wire n_2118;
 wire n_21183;
 wire n_21184;
 wire n_21185;
 wire n_2119;
 wire n_21191;
 wire n_21192;
 wire n_21197;
 wire n_21198;
 wire n_21199;
 wire n_2120;
 wire n_21200;
 wire n_21201;
 wire n_21202;
 wire n_21203;
 wire n_21204;
 wire n_21205;
 wire n_21206;
 wire n_21207;
 wire n_2121;
 wire n_21210;
 wire n_21211;
 wire n_21212;
 wire n_21214;
 wire n_21215;
 wire n_21217;
 wire n_21218;
 wire n_21219;
 wire n_21220;
 wire n_21222;
 wire n_21224;
 wire n_21229;
 wire n_2123;
 wire n_21230;
 wire n_21240;
 wire n_21241;
 wire n_21242;
 wire n_21243;
 wire n_21244;
 wire n_21245;
 wire n_21246;
 wire n_21247;
 wire n_21248;
 wire n_21249;
 wire n_2125;
 wire n_21250;
 wire n_21251;
 wire n_21254;
 wire n_21255;
 wire n_21256;
 wire n_21257;
 wire n_21258;
 wire n_2126;
 wire n_21266;
 wire n_21267;
 wire n_21268;
 wire n_21269;
 wire n_21270;
 wire n_21276;
 wire n_21277;
 wire n_21278;
 wire n_2128;
 wire n_21282;
 wire n_21283;
 wire n_21284;
 wire n_21285;
 wire n_21286;
 wire n_21287;
 wire n_21288;
 wire n_21289;
 wire n_2129;
 wire n_21290;
 wire n_21291;
 wire n_21293;
 wire n_21294;
 wire n_21295;
 wire n_213;
 wire n_2130;
 wire n_21306;
 wire n_21307;
 wire n_21308;
 wire n_21309;
 wire n_2131;
 wire n_21311;
 wire n_21317;
 wire n_21318;
 wire n_21319;
 wire n_2132;
 wire n_21322;
 wire n_2133;
 wire n_21331;
 wire n_21332;
 wire n_21333;
 wire n_21334;
 wire n_21335;
 wire n_21336;
 wire n_21337;
 wire n_21338;
 wire n_21339;
 wire n_21340;
 wire n_2135;
 wire n_21350;
 wire n_21351;
 wire n_21352;
 wire n_21353;
 wire n_21354;
 wire n_21355;
 wire n_21357;
 wire n_21359;
 wire n_2136;
 wire n_21361;
 wire n_21362;
 wire n_21363;
 wire n_21364;
 wire n_21365;
 wire n_21367;
 wire n_21368;
 wire n_21369;
 wire n_2137;
 wire n_21370;
 wire n_21371;
 wire n_21372;
 wire n_21373;
 wire n_21374;
 wire n_21375;
 wire n_21376;
 wire n_21377;
 wire n_21378;
 wire n_21379;
 wire n_2138;
 wire n_21380;
 wire n_21381;
 wire n_21382;
 wire n_21383;
 wire n_21384;
 wire n_21385;
 wire n_21386;
 wire n_21387;
 wire n_21388;
 wire n_21389;
 wire n_2139;
 wire n_21390;
 wire n_21391;
 wire n_21392;
 wire n_21393;
 wire n_21394;
 wire n_21395;
 wire n_21397;
 wire n_21398;
 wire n_21399;
 wire n_214;
 wire n_2140;
 wire n_21400;
 wire n_21401;
 wire n_21404;
 wire n_21407;
 wire n_21409;
 wire n_21410;
 wire n_21411;
 wire n_21413;
 wire n_21414;
 wire n_21415;
 wire n_21419;
 wire n_21420;
 wire n_21421;
 wire n_21422;
 wire n_21423;
 wire n_21424;
 wire n_21425;
 wire n_21426;
 wire n_21427;
 wire n_21429;
 wire n_21430;
 wire n_21434;
 wire n_21435;
 wire n_21436;
 wire n_21437;
 wire n_21438;
 wire n_21439;
 wire n_2144;
 wire n_21446;
 wire n_21447;
 wire n_21448;
 wire n_21449;
 wire n_21450;
 wire n_21452;
 wire n_21454;
 wire n_21458;
 wire n_21459;
 wire n_2146;
 wire n_21460;
 wire n_21461;
 wire n_21462;
 wire n_21463;
 wire n_21464;
 wire n_21467;
 wire n_21469;
 wire n_21471;
 wire n_21473;
 wire n_21474;
 wire n_21475;
 wire n_21476;
 wire n_21477;
 wire n_21478;
 wire n_21479;
 wire n_21480;
 wire n_21481;
 wire n_21482;
 wire n_21483;
 wire n_21484;
 wire n_21485;
 wire n_21486;
 wire n_21487;
 wire n_21489;
 wire n_21492;
 wire n_21493;
 wire n_21495;
 wire n_21496;
 wire n_21497;
 wire n_215;
 wire n_2150;
 wire n_21503;
 wire n_21504;
 wire n_21505;
 wire n_21506;
 wire n_21507;
 wire n_21508;
 wire n_21509;
 wire n_2151;
 wire n_21510;
 wire n_21511;
 wire n_21512;
 wire n_21513;
 wire n_21514;
 wire n_21515;
 wire n_21516;
 wire n_21517;
 wire n_21518;
 wire n_21519;
 wire n_21520;
 wire n_21524;
 wire n_21526;
 wire n_21527;
 wire n_21529;
 wire n_21530;
 wire n_21531;
 wire n_21532;
 wire n_21534;
 wire n_2154;
 wire n_21541;
 wire n_21543;
 wire n_21544;
 wire n_21545;
 wire n_21546;
 wire n_2155;
 wire n_21551;
 wire n_21552;
 wire n_21553;
 wire n_21554;
 wire n_21556;
 wire n_21557;
 wire n_21559;
 wire n_21560;
 wire n_21570;
 wire n_21571;
 wire n_21572;
 wire n_21573;
 wire n_21576;
 wire n_21577;
 wire n_21578;
 wire n_21579;
 wire n_2158;
 wire n_21580;
 wire n_21581;
 wire n_21582;
 wire n_21583;
 wire n_21588;
 wire n_2159;
 wire n_21593;
 wire n_21595;
 wire n_21596;
 wire n_21598;
 wire n_21599;
 wire n_216;
 wire n_2160;
 wire n_21600;
 wire n_21601;
 wire n_21606;
 wire n_21607;
 wire n_2161;
 wire n_21611;
 wire n_21612;
 wire n_21613;
 wire n_21617;
 wire n_21618;
 wire n_21619;
 wire n_2162;
 wire n_21620;
 wire n_21621;
 wire n_21622;
 wire n_21623;
 wire n_21624;
 wire n_21625;
 wire n_21626;
 wire n_21627;
 wire n_21628;
 wire n_21629;
 wire n_2163;
 wire n_21630;
 wire n_21631;
 wire n_21632;
 wire n_21633;
 wire n_21634;
 wire n_21635;
 wire n_21636;
 wire n_21637;
 wire n_21638;
 wire n_21639;
 wire n_21643;
 wire n_21644;
 wire n_21645;
 wire n_21646;
 wire n_21648;
 wire n_21649;
 wire n_2165;
 wire n_21650;
 wire n_21651;
 wire n_21654;
 wire n_21655;
 wire n_21656;
 wire n_21657;
 wire n_21658;
 wire n_21659;
 wire n_21660;
 wire n_21661;
 wire n_21662;
 wire n_21663;
 wire n_21664;
 wire n_21665;
 wire n_21666;
 wire n_21667;
 wire n_21668;
 wire n_21669;
 wire n_21673;
 wire n_21675;
 wire n_21676;
 wire n_21677;
 wire n_21678;
 wire n_21679;
 wire n_2168;
 wire n_21684;
 wire n_21685;
 wire n_21686;
 wire n_21687;
 wire n_21688;
 wire n_21689;
 wire n_2169;
 wire n_21690;
 wire n_21691;
 wire n_21692;
 wire n_21694;
 wire n_21696;
 wire n_21697;
 wire n_21698;
 wire n_21699;
 wire n_217;
 wire n_2173;
 wire n_2174;
 wire n_2176;
 wire n_2177;
 wire n_21789;
 wire n_2179;
 wire n_21793;
 wire n_21795;
 wire n_21796;
 wire n_21797;
 wire n_21798;
 wire n_218;
 wire n_2180;
 wire n_21800;
 wire n_21801;
 wire n_21802;
 wire n_21803;
 wire n_21804;
 wire n_21805;
 wire n_2181;
 wire n_2182;
 wire n_21826;
 wire n_21827;
 wire n_21828;
 wire n_21829;
 wire n_21830;
 wire n_21832;
 wire n_21835;
 wire n_21836;
 wire n_21837;
 wire n_21838;
 wire n_21839;
 wire n_21840;
 wire n_21841;
 wire n_21842;
 wire n_21845;
 wire n_21846;
 wire n_21847;
 wire n_21848;
 wire n_21849;
 wire n_21850;
 wire n_21851;
 wire n_21852;
 wire n_21853;
 wire n_21855;
 wire n_21856;
 wire n_21857;
 wire n_21858;
 wire n_21859;
 wire n_21860;
 wire n_21861;
 wire n_21862;
 wire n_21863;
 wire n_21864;
 wire n_21865;
 wire n_21866;
 wire n_21867;
 wire n_21869;
 wire n_21873;
 wire n_21875;
 wire n_21876;
 wire n_21880;
 wire n_21881;
 wire n_21882;
 wire n_21883;
 wire n_21892;
 wire n_219;
 wire n_2191;
 wire n_21911;
 wire n_21912;
 wire n_21913;
 wire n_21918;
 wire n_21919;
 wire n_21920;
 wire n_21922;
 wire n_21923;
 wire n_21924;
 wire n_21925;
 wire n_21926;
 wire n_21927;
 wire n_21928;
 wire n_21929;
 wire n_21930;
 wire n_21931;
 wire n_21932;
 wire n_21936;
 wire n_21937;
 wire n_21939;
 wire n_21941;
 wire n_21942;
 wire n_21943;
 wire n_21944;
 wire n_21945;
 wire n_21946;
 wire n_21947;
 wire n_21948;
 wire n_21949;
 wire n_21951;
 wire n_21952;
 wire n_21956;
 wire n_2196;
 wire n_21960;
 wire n_21961;
 wire n_21962;
 wire n_21963;
 wire n_21965;
 wire n_21966;
 wire n_21967;
 wire n_21968;
 wire n_21970;
 wire n_21971;
 wire n_21972;
 wire n_21973;
 wire n_21974;
 wire n_21976;
 wire n_21977;
 wire n_21978;
 wire n_21979;
 wire n_21980;
 wire n_21983;
 wire n_21984;
 wire n_21985;
 wire n_21986;
 wire n_21987;
 wire n_21988;
 wire n_21989;
 wire n_21990;
 wire n_21991;
 wire n_21994;
 wire n_21995;
 wire n_21996;
 wire n_21997;
 wire n_21998;
 wire n_21999;
 wire n_22;
 wire n_220;
 wire n_22000;
 wire n_22001;
 wire n_22002;
 wire n_22003;
 wire n_22004;
 wire n_22005;
 wire n_22011;
 wire n_22012;
 wire n_22013;
 wire n_22016;
 wire n_22017;
 wire n_22019;
 wire n_22020;
 wire n_22021;
 wire n_22022;
 wire n_22023;
 wire n_22024;
 wire n_22025;
 wire n_22026;
 wire n_22027;
 wire n_22028;
 wire n_22034;
 wire n_22035;
 wire n_22036;
 wire n_22037;
 wire n_22040;
 wire n_22041;
 wire n_22042;
 wire n_22043;
 wire n_22044;
 wire n_22045;
 wire n_22046;
 wire n_22047;
 wire n_22048;
 wire n_22049;
 wire n_22050;
 wire n_22051;
 wire n_22052;
 wire n_22053;
 wire n_22054;
 wire n_22055;
 wire n_22056;
 wire n_22057;
 wire n_22061;
 wire n_22062;
 wire n_22063;
 wire n_22064;
 wire n_22066;
 wire n_22068;
 wire n_22069;
 wire n_22071;
 wire n_22072;
 wire n_22073;
 wire n_22074;
 wire n_22076;
 wire n_22077;
 wire n_22078;
 wire n_22079;
 wire n_22080;
 wire n_22081;
 wire n_22082;
 wire n_22083;
 wire n_22084;
 wire n_22087;
 wire n_22089;
 wire n_22090;
 wire n_22092;
 wire n_22093;
 wire n_22094;
 wire n_22095;
 wire n_22096;
 wire n_22097;
 wire n_22099;
 wire n_221;
 wire n_22100;
 wire n_22101;
 wire n_22103;
 wire n_22104;
 wire n_22105;
 wire n_22110;
 wire n_22112;
 wire n_22113;
 wire n_22120;
 wire n_22121;
 wire n_22123;
 wire n_22128;
 wire n_22129;
 wire n_22138;
 wire n_22141;
 wire n_22142;
 wire n_22143;
 wire n_22147;
 wire n_22151;
 wire n_22152;
 wire n_22153;
 wire n_22154;
 wire n_22155;
 wire n_22156;
 wire n_22157;
 wire n_22158;
 wire n_22159;
 wire n_22161;
 wire n_22162;
 wire n_22164;
 wire n_22166;
 wire n_22167;
 wire n_22169;
 wire n_22170;
 wire n_22171;
 wire n_22172;
 wire n_22173;
 wire n_22174;
 wire n_22175;
 wire n_22176;
 wire n_22177;
 wire n_22178;
 wire n_22179;
 wire n_22180;
 wire n_22182;
 wire n_22183;
 wire n_22185;
 wire n_22186;
 wire n_22187;
 wire n_22188;
 wire n_22190;
 wire n_222;
 wire n_22214;
 wire n_22215;
 wire n_22216;
 wire n_22217;
 wire n_22218;
 wire n_22219;
 wire n_22220;
 wire n_22221;
 wire n_22222;
 wire n_22224;
 wire n_22229;
 wire n_22230;
 wire n_22231;
 wire n_22232;
 wire n_22234;
 wire n_22235;
 wire n_22236;
 wire n_22241;
 wire n_22242;
 wire n_22243;
 wire n_22244;
 wire n_22245;
 wire n_22246;
 wire n_22247;
 wire n_22250;
 wire n_22251;
 wire n_22252;
 wire n_22256;
 wire n_22257;
 wire n_22258;
 wire n_22259;
 wire n_22260;
 wire n_22261;
 wire n_22287;
 wire n_22290;
 wire n_22291;
 wire n_22292;
 wire n_22293;
 wire n_22294;
 wire n_22295;
 wire n_22296;
 wire n_223;
 wire n_22306;
 wire n_22307;
 wire n_22308;
 wire n_22309;
 wire n_22311;
 wire n_22312;
 wire n_22314;
 wire n_22315;
 wire n_22316;
 wire n_22317;
 wire n_22318;
 wire n_22319;
 wire n_22320;
 wire n_22321;
 wire n_22323;
 wire n_22324;
 wire n_22325;
 wire n_22326;
 wire n_22331;
 wire n_22332;
 wire n_22333;
 wire n_22334;
 wire n_22335;
 wire n_22379;
 wire n_224;
 wire n_22412;
 wire n_22413;
 wire n_22414;
 wire n_22416;
 wire n_22417;
 wire n_22418;
 wire n_22419;
 wire n_22420;
 wire n_22421;
 wire n_22422;
 wire n_22423;
 wire n_22424;
 wire n_22425;
 wire n_22426;
 wire n_22427;
 wire n_22428;
 wire n_22429;
 wire n_22430;
 wire n_22431;
 wire n_22435;
 wire n_22436;
 wire n_22437;
 wire n_22438;
 wire n_22439;
 wire n_22440;
 wire n_22441;
 wire n_22442;
 wire n_22443;
 wire n_22448;
 wire n_22451;
 wire n_22456;
 wire n_22457;
 wire n_22458;
 wire n_22459;
 wire n_22460;
 wire n_22461;
 wire n_22462;
 wire n_22463;
 wire n_22464;
 wire n_22465;
 wire n_22477;
 wire n_22478;
 wire n_22479;
 wire n_22480;
 wire n_22481;
 wire n_22482;
 wire n_22485;
 wire n_22486;
 wire n_22487;
 wire n_22488;
 wire n_22489;
 wire n_22490;
 wire n_22494;
 wire n_22495;
 wire n_22496;
 wire n_22497;
 wire n_22498;
 wire n_22499;
 wire n_225;
 wire n_22500;
 wire n_22503;
 wire n_22504;
 wire n_22506;
 wire n_22508;
 wire n_22509;
 wire n_22510;
 wire n_22511;
 wire n_22512;
 wire n_22514;
 wire n_22515;
 wire n_22516;
 wire n_22517;
 wire n_22518;
 wire n_22519;
 wire n_22520;
 wire n_22521;
 wire n_22522;
 wire n_22523;
 wire n_22524;
 wire n_22525;
 wire n_22533;
 wire n_22534;
 wire n_22535;
 wire n_22536;
 wire n_22537;
 wire n_22538;
 wire n_22539;
 wire n_22540;
 wire n_22541;
 wire n_22542;
 wire n_22543;
 wire n_22557;
 wire n_22558;
 wire n_22559;
 wire n_22560;
 wire n_22561;
 wire n_22562;
 wire n_22564;
 wire n_22565;
 wire n_22566;
 wire n_22567;
 wire n_22568;
 wire n_22594;
 wire n_22596;
 wire n_226;
 wire n_22604;
 wire n_22606;
 wire n_22608;
 wire n_22609;
 wire n_22610;
 wire n_22611;
 wire n_22612;
 wire n_22614;
 wire n_22615;
 wire n_22616;
 wire n_22617;
 wire n_22618;
 wire n_22619;
 wire n_22620;
 wire n_22621;
 wire n_22622;
 wire n_22623;
 wire n_22624;
 wire n_22625;
 wire n_22626;
 wire n_22628;
 wire n_22629;
 wire n_22630;
 wire n_22631;
 wire n_22632;
 wire n_22633;
 wire n_22634;
 wire n_22635;
 wire n_22636;
 wire n_22637;
 wire n_22638;
 wire n_2271;
 wire n_22712;
 wire n_22713;
 wire n_22714;
 wire n_22715;
 wire n_22716;
 wire n_22717;
 wire n_22718;
 wire n_22719;
 wire n_22720;
 wire n_22721;
 wire n_22724;
 wire n_22725;
 wire n_22726;
 wire n_22727;
 wire n_22728;
 wire n_22731;
 wire n_22732;
 wire n_22733;
 wire n_22734;
 wire n_22735;
 wire n_22736;
 wire n_22737;
 wire n_22738;
 wire n_22739;
 wire n_22740;
 wire n_22741;
 wire n_22742;
 wire n_22743;
 wire n_22744;
 wire n_22745;
 wire n_2275;
 wire n_2277;
 wire n_22779;
 wire n_22780;
 wire n_22781;
 wire n_22783;
 wire n_22784;
 wire n_22785;
 wire n_22786;
 wire n_22787;
 wire n_22790;
 wire n_22791;
 wire n_22792;
 wire n_22793;
 wire n_22794;
 wire n_22795;
 wire n_22796;
 wire n_22797;
 wire n_22798;
 wire n_22799;
 wire n_228;
 wire n_22800;
 wire n_22801;
 wire n_22802;
 wire n_22803;
 wire n_22804;
 wire n_22805;
 wire n_22806;
 wire n_22807;
 wire n_22808;
 wire n_22812;
 wire n_22813;
 wire n_22814;
 wire n_22815;
 wire n_22816;
 wire n_22817;
 wire n_22818;
 wire n_22819;
 wire n_22820;
 wire n_22821;
 wire n_22822;
 wire n_22823;
 wire n_22824;
 wire n_22825;
 wire n_2283;
 wire n_22834;
 wire n_22836;
 wire n_22837;
 wire n_22838;
 wire n_22839;
 wire n_22840;
 wire n_22841;
 wire n_22842;
 wire n_22843;
 wire n_22844;
 wire n_22845;
 wire n_22846;
 wire n_22847;
 wire n_22848;
 wire n_22849;
 wire n_22850;
 wire n_22851;
 wire n_22852;
 wire n_22853;
 wire n_22854;
 wire n_22856;
 wire n_22858;
 wire n_22859;
 wire n_22860;
 wire n_22861;
 wire n_22862;
 wire n_22863;
 wire n_22864;
 wire n_22865;
 wire n_22866;
 wire n_22867;
 wire n_22868;
 wire n_22869;
 wire n_22870;
 wire n_22871;
 wire n_22872;
 wire n_22873;
 wire n_22874;
 wire n_22875;
 wire n_22876;
 wire n_22877;
 wire n_22878;
 wire n_22879;
 wire n_22880;
 wire n_22881;
 wire n_22882;
 wire n_22883;
 wire n_22884;
 wire n_22885;
 wire n_22886;
 wire n_22888;
 wire n_22889;
 wire n_22890;
 wire n_22891;
 wire n_22892;
 wire n_22893;
 wire n_22894;
 wire n_22895;
 wire n_22896;
 wire n_229;
 wire n_2293;
 wire n_22948;
 wire n_22949;
 wire n_22950;
 wire n_22951;
 wire n_22952;
 wire n_22953;
 wire n_22954;
 wire n_22955;
 wire n_22956;
 wire n_22958;
 wire n_22959;
 wire n_22960;
 wire n_22962;
 wire n_22966;
 wire n_22967;
 wire n_22968;
 wire n_22969;
 wire n_22970;
 wire n_22971;
 wire n_22972;
 wire n_22973;
 wire n_22974;
 wire n_22975;
 wire n_22976;
 wire n_22977;
 wire n_22978;
 wire n_22979;
 wire n_2298;
 wire n_22980;
 wire n_22983;
 wire n_22987;
 wire n_22988;
 wire n_22989;
 wire n_22994;
 wire n_22995;
 wire n_22997;
 wire n_23;
 wire n_230;
 wire n_23000;
 wire n_23001;
 wire n_23002;
 wire n_23009;
 wire n_23010;
 wire n_23011;
 wire n_23012;
 wire n_23014;
 wire n_23015;
 wire n_23016;
 wire n_23018;
 wire n_23019;
 wire n_23020;
 wire n_23021;
 wire n_23031;
 wire n_23032;
 wire n_23033;
 wire n_23035;
 wire n_23036;
 wire n_23037;
 wire n_23038;
 wire n_23039;
 wire n_23041;
 wire n_23042;
 wire n_23043;
 wire n_23045;
 wire n_23046;
 wire n_23047;
 wire n_23049;
 wire n_23050;
 wire n_23051;
 wire n_23052;
 wire n_23053;
 wire n_23054;
 wire n_23056;
 wire n_23057;
 wire n_23058;
 wire n_23059;
 wire n_23060;
 wire n_23062;
 wire n_23063;
 wire n_23064;
 wire n_23065;
 wire n_23066;
 wire n_23067;
 wire n_23068;
 wire n_23069;
 wire n_2307;
 wire n_23070;
 wire n_23071;
 wire n_23072;
 wire n_23073;
 wire n_23074;
 wire n_23075;
 wire n_23076;
 wire n_23077;
 wire n_23078;
 wire n_23079;
 wire n_23083;
 wire n_23084;
 wire n_23085;
 wire n_23086;
 wire n_23087;
 wire n_23088;
 wire n_23090;
 wire n_23091;
 wire n_23092;
 wire n_23093;
 wire n_23094;
 wire n_23095;
 wire n_23097;
 wire n_23098;
 wire n_23099;
 wire n_231;
 wire n_23100;
 wire n_23101;
 wire n_23102;
 wire n_23103;
 wire n_23104;
 wire n_23105;
 wire n_23106;
 wire n_23108;
 wire n_23109;
 wire n_23110;
 wire n_23111;
 wire n_23112;
 wire n_23113;
 wire n_23114;
 wire n_23115;
 wire n_23116;
 wire n_23118;
 wire n_23119;
 wire n_2312;
 wire n_23120;
 wire n_23121;
 wire n_23122;
 wire n_23123;
 wire n_23124;
 wire n_23125;
 wire n_23126;
 wire n_23127;
 wire n_23128;
 wire n_23129;
 wire n_23130;
 wire n_23131;
 wire n_23132;
 wire n_23133;
 wire n_23134;
 wire n_23135;
 wire n_23138;
 wire n_23139;
 wire n_23165;
 wire n_23166;
 wire n_23167;
 wire n_23168;
 wire n_23169;
 wire n_23170;
 wire n_23174;
 wire n_23175;
 wire n_23192;
 wire n_23193;
 wire n_23194;
 wire n_23195;
 wire n_23196;
 wire n_23197;
 wire n_232;
 wire n_23219;
 wire n_23220;
 wire n_23221;
 wire n_23222;
 wire n_23223;
 wire n_23224;
 wire n_23225;
 wire n_23226;
 wire n_23227;
 wire n_23228;
 wire n_23229;
 wire n_23230;
 wire n_23231;
 wire n_23232;
 wire n_23233;
 wire n_23234;
 wire n_23235;
 wire n_23236;
 wire n_2325;
 wire n_23266;
 wire n_23268;
 wire n_23272;
 wire n_23276;
 wire n_23277;
 wire n_23278;
 wire n_23280;
 wire n_23289;
 wire n_23290;
 wire n_23291;
 wire n_23296;
 wire n_2331;
 wire n_2335;
 wire n_23365;
 wire n_23366;
 wire n_23367;
 wire n_23368;
 wire n_2337;
 wire n_23372;
 wire n_23373;
 wire n_23374;
 wire n_23375;
 wire n_23376;
 wire n_23378;
 wire n_23379;
 wire n_23380;
 wire n_23385;
 wire n_23386;
 wire n_23387;
 wire n_23388;
 wire n_23389;
 wire n_2339;
 wire n_23390;
 wire n_23391;
 wire n_23392;
 wire n_23393;
 wire n_23394;
 wire n_23398;
 wire n_23399;
 wire n_23400;
 wire n_23401;
 wire n_23402;
 wire n_23403;
 wire n_23404;
 wire n_23407;
 wire n_23408;
 wire n_23409;
 wire n_23410;
 wire n_23411;
 wire n_23412;
 wire n_23413;
 wire n_23414;
 wire n_23415;
 wire n_23416;
 wire n_23417;
 wire n_23418;
 wire n_23419;
 wire n_23420;
 wire n_23421;
 wire n_23422;
 wire n_23423;
 wire n_23424;
 wire n_23425;
 wire n_23426;
 wire n_23427;
 wire n_23428;
 wire n_23429;
 wire n_23430;
 wire n_23431;
 wire n_23432;
 wire n_23433;
 wire n_23434;
 wire n_23435;
 wire n_23436;
 wire n_23437;
 wire n_23438;
 wire n_23439;
 wire n_23440;
 wire n_23441;
 wire n_23442;
 wire n_23443;
 wire n_23444;
 wire n_23445;
 wire n_23446;
 wire n_23447;
 wire n_23448;
 wire n_23449;
 wire n_23450;
 wire n_23451;
 wire n_23461;
 wire n_23462;
 wire n_23463;
 wire n_23466;
 wire n_23467;
 wire n_23468;
 wire n_23469;
 wire n_23470;
 wire n_23471;
 wire n_23493;
 wire n_23495;
 wire n_23497;
 wire n_23541;
 wire n_23546;
 wire n_23547;
 wire n_23548;
 wire n_23549;
 wire n_23550;
 wire n_23551;
 wire n_23552;
 wire n_23553;
 wire n_23554;
 wire n_23555;
 wire n_23557;
 wire n_23559;
 wire n_23560;
 wire n_23561;
 wire n_23562;
 wire n_23563;
 wire n_23564;
 wire n_23565;
 wire n_23566;
 wire n_23567;
 wire n_23568;
 wire n_23569;
 wire n_23573;
 wire n_23578;
 wire n_23579;
 wire n_23580;
 wire n_23581;
 wire n_23582;
 wire n_2359;
 wire n_236;
 wire n_2364;
 wire n_23658;
 wire n_23659;
 wire n_2366;
 wire n_23660;
 wire n_23661;
 wire n_23662;
 wire n_23663;
 wire n_23664;
 wire n_23665;
 wire n_23666;
 wire n_23667;
 wire n_23668;
 wire n_23669;
 wire n_23670;
 wire n_23682;
 wire n_23683;
 wire n_23684;
 wire n_23685;
 wire n_237;
 wire n_23738;
 wire n_23753;
 wire n_2377;
 wire n_23772;
 wire n_23776;
 wire n_23789;
 wire n_23790;
 wire n_238;
 wire n_2381;
 wire n_23818;
 wire n_23819;
 wire n_23820;
 wire n_23824;
 wire n_23825;
 wire n_23829;
 wire n_23830;
 wire n_23832;
 wire n_23833;
 wire n_23834;
 wire n_23835;
 wire n_23837;
 wire n_2384;
 wire n_23894;
 wire n_23895;
 wire n_2392;
 wire n_23931;
 wire n_23932;
 wire n_23934;
 wire n_23935;
 wire n_23936;
 wire n_23941;
 wire n_23942;
 wire n_23972;
 wire n_23973;
 wire n_23974;
 wire n_23975;
 wire n_23976;
 wire n_2398;
 wire n_23985;
 wire n_23986;
 wire n_23987;
 wire n_23988;
 wire n_24;
 wire n_240;
 wire n_2400;
 wire n_24021;
 wire n_24022;
 wire n_24024;
 wire n_24025;
 wire n_24027;
 wire n_24028;
 wire n_24029;
 wire n_24033;
 wire n_24034;
 wire n_24035;
 wire n_24102;
 wire n_24103;
 wire n_24104;
 wire n_24105;
 wire n_24106;
 wire n_24107;
 wire n_24152;
 wire n_24153;
 wire n_24166;
 wire n_24167;
 wire n_24168;
 wire n_24169;
 wire n_24171;
 wire n_24172;
 wire n_24173;
 wire n_24174;
 wire n_24175;
 wire n_24176;
 wire n_24177;
 wire n_24178;
 wire n_24179;
 wire n_24181;
 wire n_242;
 wire n_24200;
 wire n_24201;
 wire n_24202;
 wire n_24203;
 wire n_24204;
 wire n_24206;
 wire n_24207;
 wire n_24208;
 wire n_24210;
 wire n_24212;
 wire n_24213;
 wire n_24230;
 wire n_24231;
 wire n_2429;
 wire n_243;
 wire n_2431;
 wire n_2435;
 wire n_2437;
 wire n_2439;
 wire n_244;
 wire n_24402;
 wire n_24403;
 wire n_24404;
 wire n_24405;
 wire n_2441;
 wire n_2442;
 wire n_2444;
 wire n_2445;
 wire n_245;
 wire n_246;
 wire n_2465;
 wire n_2466;
 wire n_24669;
 wire n_24670;
 wire n_24671;
 wire n_24678;
 wire n_24679;
 wire n_24680;
 wire n_24681;
 wire n_24682;
 wire n_24683;
 wire n_24684;
 wire n_24710;
 wire n_24711;
 wire n_24712;
 wire n_24751;
 wire n_24752;
 wire n_24753;
 wire n_24754;
 wire n_24766;
 wire n_24767;
 wire n_24768;
 wire n_24769;
 wire n_24770;
 wire n_24912;
 wire n_24913;
 wire n_24914;
 wire n_24915;
 wire n_24916;
 wire n_24917;
 wire n_24976;
 wire n_24977;
 wire n_24978;
 wire n_24979;
 wire n_2499;
 wire n_25;
 wire n_250;
 wire n_2507;
 wire n_251;
 wire n_25128;
 wire n_25130;
 wire n_25131;
 wire n_25132;
 wire n_252;
 wire n_2524;
 wire n_2525;
 wire n_25292;
 wire n_25294;
 wire n_25295;
 wire n_25296;
 wire n_25298;
 wire n_25299;
 wire n_253;
 wire n_25300;
 wire n_25301;
 wire n_25302;
 wire n_25303;
 wire n_25311;
 wire n_25312;
 wire n_25313;
 wire n_25335;
 wire n_25336;
 wire n_25337;
 wire n_254;
 wire n_25425;
 wire n_25426;
 wire n_25427;
 wire n_25428;
 wire n_25429;
 wire n_25430;
 wire n_25431;
 wire n_2544;
 wire n_25445;
 wire n_25446;
 wire n_25447;
 wire n_25448;
 wire n_25449;
 wire n_25450;
 wire n_25499;
 wire n_255;
 wire n_25500;
 wire n_25502;
 wire n_25503;
 wire n_25504;
 wire n_2552;
 wire n_25596;
 wire n_25597;
 wire n_25598;
 wire n_25599;
 wire n_256;
 wire n_25602;
 wire n_25603;
 wire n_25604;
 wire n_25605;
 wire n_25606;
 wire n_25607;
 wire n_2562;
 wire n_2564;
 wire n_2566;
 wire n_257;
 wire n_2578;
 wire n_258;
 wire n_2580;
 wire n_2582;
 wire n_25833;
 wire n_2588;
 wire n_25881;
 wire n_25882;
 wire n_259;
 wire n_2591;
 wire n_2592;
 wire n_25921;
 wire n_25963;
 wire n_25971;
 wire n_25976;
 wire n_25977;
 wire n_25978;
 wire n_25979;
 wire n_25980;
 wire n_25981;
 wire n_25982;
 wire n_25983;
 wire n_25984;
 wire n_25987;
 wire n_25988;
 wire n_25989;
 wire n_25990;
 wire n_25992;
 wire n_25996;
 wire n_25999;
 wire n_26;
 wire n_260;
 wire n_26000;
 wire n_26003;
 wire n_26004;
 wire n_26005;
 wire n_26008;
 wire n_26009;
 wire n_26010;
 wire n_26011;
 wire n_26012;
 wire n_26015;
 wire n_26016;
 wire n_26017;
 wire n_26021;
 wire n_26024;
 wire n_26026;
 wire n_26028;
 wire n_26029;
 wire n_26030;
 wire n_26031;
 wire n_26032;
 wire n_26033;
 wire n_26035;
 wire n_26037;
 wire n_26038;
 wire n_26039;
 wire n_26040;
 wire n_26041;
 wire n_26044;
 wire n_26045;
 wire n_26046;
 wire n_26049;
 wire n_26051;
 wire n_26052;
 wire n_26053;
 wire n_26054;
 wire n_26055;
 wire n_26057;
 wire n_26058;
 wire n_26059;
 wire n_26060;
 wire n_26062;
 wire n_26063;
 wire n_26066;
 wire n_26068;
 wire n_26071;
 wire n_26073;
 wire n_26074;
 wire n_26076;
 wire n_26077;
 wire n_26078;
 wire n_26079;
 wire n_26080;
 wire n_26081;
 wire n_26083;
 wire n_26089;
 wire n_26091;
 wire n_26093;
 wire n_26097;
 wire n_26098;
 wire n_26099;
 wire n_261;
 wire n_26100;
 wire n_26101;
 wire n_26102;
 wire n_26103;
 wire n_26105;
 wire n_26107;
 wire n_26108;
 wire n_26109;
 wire n_26110;
 wire n_26111;
 wire n_26112;
 wire n_26113;
 wire n_26114;
 wire n_26117;
 wire n_26118;
 wire n_26119;
 wire n_26120;
 wire n_26121;
 wire n_26122;
 wire n_26123;
 wire n_26124;
 wire n_26125;
 wire n_26126;
 wire n_26127;
 wire n_26128;
 wire n_26129;
 wire n_26130;
 wire n_26131;
 wire n_26132;
 wire n_26133;
 wire n_26134;
 wire n_26135;
 wire n_26137;
 wire n_26138;
 wire n_26139;
 wire n_26140;
 wire n_26141;
 wire n_26142;
 wire n_26143;
 wire n_26144;
 wire n_26145;
 wire n_26146;
 wire n_26147;
 wire n_26148;
 wire n_26149;
 wire n_26150;
 wire n_26151;
 wire n_26152;
 wire n_26153;
 wire n_26159;
 wire n_26164;
 wire n_26166;
 wire n_26167;
 wire n_26168;
 wire n_26169;
 wire n_26170;
 wire n_26172;
 wire n_26173;
 wire n_26174;
 wire n_26175;
 wire n_26177;
 wire n_26178;
 wire n_26179;
 wire n_26180;
 wire n_26181;
 wire n_26183;
 wire n_26184;
 wire n_26186;
 wire n_26187;
 wire n_26189;
 wire n_26190;
 wire n_26191;
 wire n_26193;
 wire n_26194;
 wire n_26196;
 wire n_262;
 wire n_2620;
 wire n_26200;
 wire n_26202;
 wire n_26207;
 wire n_26208;
 wire n_26210;
 wire n_26212;
 wire n_26213;
 wire n_26214;
 wire n_26215;
 wire n_26216;
 wire n_26218;
 wire n_26221;
 wire n_26222;
 wire n_26224;
 wire n_26226;
 wire n_26227;
 wire n_26228;
 wire n_26231;
 wire n_26235;
 wire n_26236;
 wire n_26237;
 wire n_26238;
 wire n_26239;
 wire n_26241;
 wire n_26242;
 wire n_26243;
 wire n_26244;
 wire n_26245;
 wire n_26247;
 wire n_26249;
 wire n_26250;
 wire n_26251;
 wire n_26252;
 wire n_26255;
 wire n_26256;
 wire n_26257;
 wire n_26258;
 wire n_26264;
 wire n_26266;
 wire n_26267;
 wire n_263;
 wire n_2634;
 wire n_2642;
 wire n_265;
 wire n_2657;
 wire n_266;
 wire n_2663;
 wire n_267;
 wire n_2673;
 wire n_268;
 wire n_2685;
 wire n_2686;
 wire n_2689;
 wire n_269;
 wire n_2694;
 wire n_2697;
 wire n_27;
 wire n_2700;
 wire n_2711;
 wire n_2718;
 wire n_272;
 wire n_2728;
 wire n_273;
 wire n_2735;
 wire n_2741;
 wire n_2744;
 wire n_2746;
 wire n_2747;
 wire n_275;
 wire n_276;
 wire n_2764;
 wire n_2766;
 wire n_277;
 wire n_2781;
 wire n_2785;
 wire n_2789;
 wire n_279;
 wire n_2791;
 wire n_2793;
 wire n_28;
 wire n_280;
 wire n_2801;
 wire n_2805;
 wire n_281;
 wire n_2820;
 wire n_2821;
 wire n_2825;
 wire n_2827;
 wire n_283;
 wire n_2831;
 wire n_2836;
 wire n_284;
 wire n_2841;
 wire n_2848;
 wire n_285;
 wire n_2850;
 wire n_2852;
 wire n_2855;
 wire n_286;
 wire n_2864;
 wire n_2865;
 wire n_287;
 wire n_2873;
 wire n_2877;
 wire n_288;
 wire n_2883;
 wire n_2887;
 wire n_289;
 wire n_2891;
 wire n_2893;
 wire n_2897;
 wire n_29;
 wire n_290;
 wire n_2901;
 wire n_2903;
 wire n_291;
 wire n_292;
 wire n_2922;
 wire n_2927;
 wire n_293;
 wire n_2930;
 wire n_2934;
 wire n_2939;
 wire n_294;
 wire n_2940;
 wire n_2943;
 wire n_2944;
 wire n_2945;
 wire n_295;
 wire n_2958;
 wire n_296;
 wire n_2962;
 wire n_2965;
 wire n_2966;
 wire n_297;
 wire n_298;
 wire n_2985;
 wire n_299;
 wire n_2990;
 wire n_3;
 wire n_30;
 wire n_300;
 wire n_301;
 wire n_3011;
 wire n_3030;
 wire n_3032;
 wire n_304;
 wire n_305;
 wire n_306;
 wire n_307;
 wire n_308;
 wire n_3088;
 wire n_309;
 wire n_3090;
 wire n_31;
 wire n_310;
 wire n_3107;
 wire n_311;
 wire n_3112;
 wire n_3113;
 wire n_312;
 wire n_313;
 wire n_314;
 wire n_3148;
 wire n_3149;
 wire n_315;
 wire n_3150;
 wire n_316;
 wire n_3168;
 wire n_317;
 wire n_3170;
 wire n_318;
 wire n_3181;
 wire n_319;
 wire n_3190;
 wire n_32;
 wire n_320;
 wire n_3204;
 wire n_3206;
 wire n_3208;
 wire n_321;
 wire n_3210;
 wire n_3212;
 wire n_3214;
 wire n_3218;
 wire n_322;
 wire n_3224;
 wire n_3229;
 wire n_323;
 wire n_3231;
 wire n_3233;
 wire n_3235;
 wire n_3237;
 wire n_3239;
 wire n_324;
 wire n_3243;
 wire n_3246;
 wire n_325;
 wire n_326;
 wire n_3260;
 wire n_3265;
 wire n_3266;
 wire n_327;
 wire n_3275;
 wire n_3279;
 wire n_328;
 wire n_329;
 wire n_33;
 wire n_330;
 wire n_3309;
 wire n_331;
 wire n_3314;
 wire n_3317;
 wire n_332;
 wire n_333;
 wire n_3331;
 wire n_3332;
 wire n_334;
 wire n_335;
 wire n_3358;
 wire n_336;
 wire n_3360;
 wire n_3364;
 wire n_3366;
 wire n_337;
 wire n_3374;
 wire n_3375;
 wire n_3376;
 wire n_338;
 wire n_339;
 wire n_3396;
 wire n_3398;
 wire n_34;
 wire n_3408;
 wire n_3409;
 wire n_341;
 wire n_343;
 wire n_3433;
 wire n_3436;
 wire n_344;
 wire n_3443;
 wire n_3445;
 wire n_3450;
 wire n_3454;
 wire n_3456;
 wire n_3457;
 wire n_3459;
 wire n_346;
 wire n_3461;
 wire n_3463;
 wire n_3468;
 wire n_3469;
 wire n_347;
 wire n_3474;
 wire n_3479;
 wire n_348;
 wire n_3491;
 wire n_3493;
 wire n_35;
 wire n_3504;
 wire n_351;
 wire n_3511;
 wire n_3516;
 wire n_3521;
 wire n_3522;
 wire n_3527;
 wire n_3528;
 wire n_353;
 wire n_354;
 wire n_3547;
 wire n_3548;
 wire n_355;
 wire n_3552;
 wire n_3553;
 wire n_3557;
 wire n_3558;
 wire n_3560;
 wire n_3562;
 wire n_358;
 wire n_359;
 wire n_3591;
 wire n_3592;
 wire n_3593;
 wire n_36;
 wire n_360;
 wire n_3611;
 wire n_3615;
 wire n_3619;
 wire n_3630;
 wire n_3633;
 wire n_364;
 wire n_3642;
 wire n_3644;
 wire n_3645;
 wire n_3647;
 wire n_3649;
 wire n_365;
 wire n_3650;
 wire n_3652;
 wire n_3654;
 wire n_3655;
 wire n_3657;
 wire n_3659;
 wire n_366;
 wire n_3661;
 wire n_3668;
 wire n_3669;
 wire n_3679;
 wire n_368;
 wire n_3681;
 wire n_3685;
 wire n_3686;
 wire n_3687;
 wire n_37;
 wire n_370;
 wire n_3706;
 wire n_3709;
 wire n_3711;
 wire n_3713;
 wire n_3714;
 wire n_372;
 wire n_3729;
 wire n_373;
 wire n_3736;
 wire n_3737;
 wire n_3738;
 wire n_374;
 wire n_3746;
 wire n_3759;
 wire n_376;
 wire n_3760;
 wire n_3761;
 wire n_3766;
 wire n_3770;
 wire n_3782;
 wire n_3795;
 wire n_3796;
 wire n_38;
 wire n_3806;
 wire n_381;
 wire n_3815;
 wire n_3817;
 wire n_3819;
 wire n_382;
 wire n_3823;
 wire n_3827;
 wire n_3833;
 wire n_385;
 wire n_3860;
 wire n_3868;
 wire n_3873;
 wire n_3877;
 wire n_3878;
 wire n_388;
 wire n_3880;
 wire n_3882;
 wire n_3893;
 wire n_39;
 wire n_3901;
 wire n_3905;
 wire n_3907;
 wire n_391;
 wire n_3915;
 wire n_3917;
 wire n_3918;
 wire n_3922;
 wire n_3923;
 wire n_3938;
 wire n_3942;
 wire n_3944;
 wire n_3946;
 wire n_395;
 wire n_3950;
 wire n_3953;
 wire n_3955;
 wire n_3957;
 wire n_3963;
 wire n_3965;
 wire n_397;
 wire n_3971;
 wire n_3973;
 wire n_3975;
 wire n_398;
 wire n_3983;
 wire n_3987;
 wire n_3988;
 wire n_3990;
 wire n_4;
 wire n_40;
 wire n_400;
 wire n_4012;
 wire n_4017;
 wire n_402;
 wire n_4022;
 wire n_4024;
 wire n_4026;
 wire n_4029;
 wire n_403;
 wire n_4031;
 wire n_4038;
 wire n_4041;
 wire n_4044;
 wire n_4048;
 wire n_405;
 wire n_406;
 wire n_4061;
 wire n_4062;
 wire n_4068;
 wire n_407;
 wire n_4070;
 wire n_4072;
 wire n_4074;
 wire n_4075;
 wire n_4079;
 wire n_4082;
 wire n_4084;
 wire n_4085;
 wire n_4087;
 wire n_4089;
 wire n_4095;
 wire n_41;
 wire n_4101;
 wire n_4102;
 wire n_4107;
 wire n_411;
 wire n_4123;
 wire n_4124;
 wire n_413;
 wire n_4138;
 wire n_414;
 wire n_4140;
 wire n_4151;
 wire n_416;
 wire n_417;
 wire n_418;
 wire n_4193;
 wire n_4197;
 wire n_4199;
 wire n_42;
 wire n_422;
 wire n_4224;
 wire n_423;
 wire n_4230;
 wire n_4231;
 wire n_4233;
 wire n_4234;
 wire n_4239;
 wire n_4245;
 wire n_4246;
 wire n_4248;
 wire n_425;
 wire n_4250;
 wire n_4251;
 wire n_4253;
 wire n_4262;
 wire n_4263;
 wire n_4268;
 wire n_4275;
 wire n_428;
 wire n_4286;
 wire n_4287;
 wire n_429;
 wire n_43;
 wire n_431;
 wire n_4314;
 wire n_4315;
 wire n_432;
 wire n_433;
 wire n_4331;
 wire n_434;
 wire n_4341;
 wire n_4349;
 wire n_4354;
 wire n_4365;
 wire n_4367;
 wire n_4377;
 wire n_4385;
 wire n_4386;
 wire n_44;
 wire n_440;
 wire n_4403;
 wire n_4404;
 wire n_4408;
 wire n_441;
 wire n_4410;
 wire n_4412;
 wire n_4413;
 wire n_4414;
 wire n_4415;
 wire n_4416;
 wire n_4417;
 wire n_4418;
 wire n_4419;
 wire n_4429;
 wire n_443;
 wire n_4430;
 wire n_4434;
 wire n_4435;
 wire n_4438;
 wire n_4439;
 wire n_444;
 wire n_4443;
 wire n_445;
 wire n_4451;
 wire n_446;
 wire n_4462;
 wire n_4463;
 wire n_4474;
 wire n_448;
 wire n_4480;
 wire n_4487;
 wire n_449;
 wire n_45;
 wire n_4515;
 wire n_4518;
 wire n_452;
 wire n_4521;
 wire n_4528;
 wire n_453;
 wire n_4539;
 wire n_4541;
 wire n_4549;
 wire n_4550;
 wire n_4553;
 wire n_4555;
 wire n_4565;
 wire n_457;
 wire n_46;
 wire n_460;
 wire n_463;
 wire n_464;
 wire n_4645;
 wire n_465;
 wire n_466;
 wire n_4665;
 wire n_467;
 wire n_4671;
 wire n_468;
 wire n_469;
 wire n_47;
 wire n_470;
 wire n_471;
 wire n_472;
 wire n_473;
 wire n_474;
 wire n_475;
 wire n_476;
 wire n_4762;
 wire n_4764;
 wire n_4767;
 wire n_4768;
 wire n_4769;
 wire n_477;
 wire n_4771;
 wire n_4772;
 wire n_4773;
 wire n_4777;
 wire n_4778;
 wire n_4779;
 wire n_478;
 wire n_4780;
 wire n_4782;
 wire n_4783;
 wire n_4784;
 wire n_4786;
 wire n_4787;
 wire n_4788;
 wire n_479;
 wire n_4790;
 wire n_4791;
 wire n_4793;
 wire n_4795;
 wire n_4796;
 wire n_48;
 wire n_480;
 wire n_4805;
 wire n_481;
 wire n_4810;
 wire n_482;
 wire n_4826;
 wire n_483;
 wire n_4831;
 wire n_4833;
 wire n_484;
 wire n_4842;
 wire n_4843;
 wire n_485;
 wire n_4856;
 wire n_486;
 wire n_4861;
 wire n_4864;
 wire n_4865;
 wire n_4866;
 wire n_487;
 wire n_488;
 wire n_489;
 wire n_49;
 wire n_490;
 wire n_4902;
 wire n_4903;
 wire n_4904;
 wire n_4906;
 wire n_4907;
 wire n_491;
 wire n_492;
 wire n_493;
 wire n_494;
 wire n_495;
 wire n_4951;
 wire n_4956;
 wire n_4957;
 wire n_496;
 wire n_4965;
 wire n_4967;
 wire n_4968;
 wire n_4969;
 wire n_497;
 wire n_4970;
 wire n_498;
 wire n_499;
 wire n_5;
 wire n_50;
 wire n_500;
 wire n_501;
 wire n_502;
 wire n_503;
 wire n_504;
 wire n_5045;
 wire n_5047;
 wire n_5048;
 wire n_505;
 wire n_506;
 wire n_5065;
 wire n_507;
 wire n_508;
 wire n_509;
 wire n_510;
 wire n_511;
 wire n_512;
 wire n_5126;
 wire n_5129;
 wire n_513;
 wire n_5131;
 wire n_5133;
 wire n_5137;
 wire n_515;
 wire n_516;
 wire n_517;
 wire n_518;
 wire n_519;
 wire n_520;
 wire n_521;
 wire n_522;
 wire n_523;
 wire n_524;
 wire n_525;
 wire n_526;
 wire n_527;
 wire n_5276;
 wire n_5277;
 wire n_528;
 wire n_529;
 wire n_53;
 wire n_530;
 wire n_5300;
 wire n_5301;
 wire n_531;
 wire n_532;
 wire n_5321;
 wire n_5322;
 wire n_5323;
 wire n_5324;
 wire n_5329;
 wire n_533;
 wire n_5330;
 wire n_5331;
 wire n_5332;
 wire n_5334;
 wire n_5339;
 wire n_534;
 wire n_5340;
 wire n_5342;
 wire n_5343;
 wire n_5344;
 wire n_5345;
 wire n_5346;
 wire n_5347;
 wire n_5348;
 wire n_5349;
 wire n_535;
 wire n_5351;
 wire n_536;
 wire n_5368;
 wire n_5369;
 wire n_537;
 wire n_5371;
 wire n_5372;
 wire n_5375;
 wire n_5376;
 wire n_5377;
 wire n_5378;
 wire n_5379;
 wire n_538;
 wire n_5380;
 wire n_5383;
 wire n_5385;
 wire n_539;
 wire n_5393;
 wire n_5398;
 wire n_5399;
 wire n_54;
 wire n_540;
 wire n_5400;
 wire n_5409;
 wire n_541;
 wire n_5410;
 wire n_5411;
 wire n_5412;
 wire n_5413;
 wire n_542;
 wire n_5420;
 wire n_5421;
 wire n_5422;
 wire n_5423;
 wire n_5426;
 wire n_5427;
 wire n_5428;
 wire n_5429;
 wire n_543;
 wire n_5430;
 wire n_5431;
 wire n_5432;
 wire n_5433;
 wire n_5438;
 wire n_5439;
 wire n_544;
 wire n_5440;
 wire n_5441;
 wire n_5442;
 wire n_5443;
 wire n_5444;
 wire n_5447;
 wire n_5448;
 wire n_5449;
 wire n_545;
 wire n_5450;
 wire n_5451;
 wire n_5453;
 wire n_5454;
 wire n_5456;
 wire n_5457;
 wire n_546;
 wire n_547;
 wire n_5471;
 wire n_5473;
 wire n_548;
 wire n_5487;
 wire n_549;
 wire n_5491;
 wire n_5492;
 wire n_5493;
 wire n_5494;
 wire n_55;
 wire n_550;
 wire n_5504;
 wire n_5505;
 wire n_5506;
 wire n_5507;
 wire n_5508;
 wire n_5509;
 wire n_551;
 wire n_5510;
 wire n_5511;
 wire n_5512;
 wire n_5513;
 wire n_5514;
 wire n_5515;
 wire n_5516;
 wire n_5517;
 wire n_552;
 wire n_5529;
 wire n_553;
 wire n_5536;
 wire n_554;
 wire n_5544;
 wire n_5548;
 wire n_5549;
 wire n_555;
 wire n_5553;
 wire n_556;
 wire n_5564;
 wire n_557;
 wire n_5570;
 wire n_5575;
 wire n_558;
 wire n_5582;
 wire n_5583;
 wire n_5584;
 wire n_5589;
 wire n_559;
 wire n_5593;
 wire n_56;
 wire n_560;
 wire n_5602;
 wire n_561;
 wire n_5616;
 wire n_5617;
 wire n_562;
 wire n_5627;
 wire n_563;
 wire n_5630;
 wire n_5637;
 wire n_5639;
 wire n_564;
 wire n_5640;
 wire n_5641;
 wire n_5643;
 wire n_5644;
 wire n_5645;
 wire n_5649;
 wire n_565;
 wire n_566;
 wire n_5660;
 wire n_5664;
 wire n_567;
 wire n_5679;
 wire n_568;
 wire n_5680;
 wire n_5681;
 wire n_5683;
 wire n_569;
 wire n_5697;
 wire n_57;
 wire n_570;
 wire n_571;
 wire n_5719;
 wire n_572;
 wire n_5724;
 wire n_573;
 wire n_5733;
 wire n_5737;
 wire n_5738;
 wire n_5739;
 wire n_574;
 wire n_5740;
 wire n_5741;
 wire n_5742;
 wire n_5743;
 wire n_5744;
 wire n_575;
 wire n_5751;
 wire n_576;
 wire n_577;
 wire n_578;
 wire n_5780;
 wire n_5781;
 wire n_5783;
 wire n_5784;
 wire n_5787;
 wire n_579;
 wire n_5792;
 wire n_5793;
 wire n_5794;
 wire n_5796;
 wire n_5798;
 wire n_5799;
 wire n_58;
 wire n_580;
 wire n_5800;
 wire n_5804;
 wire n_5806;
 wire n_581;
 wire n_5811;
 wire n_5815;
 wire n_5817;
 wire n_582;
 wire n_5826;
 wire n_583;
 wire n_584;
 wire n_5840;
 wire n_5841;
 wire n_5842;
 wire n_5849;
 wire n_585;
 wire n_586;
 wire n_5867;
 wire n_5869;
 wire n_587;
 wire n_5870;
 wire n_5872;
 wire n_5873;
 wire n_5874;
 wire n_588;
 wire n_5880;
 wire n_5881;
 wire n_5886;
 wire n_589;
 wire n_5890;
 wire n_5894;
 wire n_5895;
 wire n_5896;
 wire n_59;
 wire n_590;
 wire n_5903;
 wire n_5904;
 wire n_5909;
 wire n_591;
 wire n_5910;
 wire n_592;
 wire n_5929;
 wire n_593;
 wire n_5930;
 wire n_5935;
 wire n_5936;
 wire n_594;
 wire n_5941;
 wire n_5943;
 wire n_5944;
 wire n_5948;
 wire n_595;
 wire n_5951;
 wire n_5953;
 wire n_5954;
 wire n_5955;
 wire n_5959;
 wire n_596;
 wire n_5961;
 wire n_597;
 wire n_598;
 wire n_5980;
 wire n_5981;
 wire n_5982;
 wire n_5983;
 wire n_5985;
 wire n_5986;
 wire n_5988;
 wire n_599;
 wire n_5990;
 wire n_5991;
 wire n_5994;
 wire n_5996;
 wire n_6;
 wire n_60;
 wire n_600;
 wire n_6008;
 wire n_601;
 wire n_6016;
 wire n_6017;
 wire n_6019;
 wire n_602;
 wire n_6022;
 wire n_6024;
 wire n_6025;
 wire n_603;
 wire n_6030;
 wire n_6031;
 wire n_6032;
 wire n_6033;
 wire n_6034;
 wire n_6035;
 wire n_6037;
 wire n_6038;
 wire n_6039;
 wire n_604;
 wire n_6043;
 wire n_6044;
 wire n_6045;
 wire n_605;
 wire n_606;
 wire n_6062;
 wire n_6063;
 wire n_607;
 wire n_6076;
 wire n_6078;
 wire n_6079;
 wire n_608;
 wire n_6082;
 wire n_609;
 wire n_6094;
 wire n_6097;
 wire n_6098;
 wire n_6099;
 wire n_61;
 wire n_610;
 wire n_6100;
 wire n_6102;
 wire n_6107;
 wire n_6109;
 wire n_611;
 wire n_6113;
 wire n_6114;
 wire n_6115;
 wire n_6116;
 wire n_6117;
 wire n_6119;
 wire n_612;
 wire n_6125;
 wire n_6128;
 wire n_613;
 wire n_6131;
 wire n_614;
 wire n_6141;
 wire n_6144;
 wire n_6145;
 wire n_6147;
 wire n_6148;
 wire n_6149;
 wire n_615;
 wire n_6150;
 wire n_6151;
 wire n_6152;
 wire n_6153;
 wire n_6156;
 wire n_6157;
 wire n_616;
 wire n_617;
 wire n_6179;
 wire n_618;
 wire n_6186;
 wire n_6189;
 wire n_619;
 wire n_6190;
 wire n_6191;
 wire n_6194;
 wire n_6198;
 wire n_6199;
 wire n_62;
 wire n_620;
 wire n_6200;
 wire n_6201;
 wire n_6202;
 wire n_6203;
 wire n_6204;
 wire n_6205;
 wire n_6209;
 wire n_621;
 wire n_6210;
 wire n_6211;
 wire n_6218;
 wire n_6219;
 wire n_622;
 wire n_6220;
 wire n_6221;
 wire n_6222;
 wire n_6223;
 wire n_6224;
 wire n_6225;
 wire n_623;
 wire n_6230;
 wire n_6231;
 wire n_6232;
 wire n_6233;
 wire n_6234;
 wire n_6235;
 wire n_6237;
 wire n_6238;
 wire n_624;
 wire n_6240;
 wire n_6241;
 wire n_6242;
 wire n_6243;
 wire n_625;
 wire n_6251;
 wire n_6253;
 wire n_6254;
 wire n_6255;
 wire n_6256;
 wire n_6257;
 wire n_626;
 wire n_6264;
 wire n_6265;
 wire n_6266;
 wire n_627;
 wire n_6279;
 wire n_628;
 wire n_6280;
 wire n_6284;
 wire n_629;
 wire n_6295;
 wire n_6296;
 wire n_6298;
 wire n_63;
 wire n_630;
 wire n_6300;
 wire n_6301;
 wire n_6302;
 wire n_6303;
 wire n_6304;
 wire n_6305;
 wire n_631;
 wire n_6313;
 wire n_632;
 wire n_6323;
 wire n_6324;
 wire n_6325;
 wire n_6326;
 wire n_6327;
 wire n_6329;
 wire n_633;
 wire n_6331;
 wire n_6339;
 wire n_634;
 wire n_6341;
 wire n_6342;
 wire n_6343;
 wire n_6348;
 wire n_6349;
 wire n_635;
 wire n_6350;
 wire n_6351;
 wire n_6352;
 wire n_6353;
 wire n_6354;
 wire n_636;
 wire n_6360;
 wire n_6361;
 wire n_6365;
 wire n_6366;
 wire n_6368;
 wire n_6369;
 wire n_637;
 wire n_6370;
 wire n_6371;
 wire n_6372;
 wire n_6373;
 wire n_6377;
 wire n_638;
 wire n_6381;
 wire n_6382;
 wire n_6383;
 wire n_6384;
 wire n_6385;
 wire n_639;
 wire n_6391;
 wire n_6392;
 wire n_6394;
 wire n_6395;
 wire n_6396;
 wire n_6397;
 wire n_6399;
 wire n_64;
 wire n_640;
 wire n_6400;
 wire n_6401;
 wire n_6404;
 wire n_6406;
 wire n_6409;
 wire n_641;
 wire n_6410;
 wire n_6411;
 wire n_642;
 wire n_6420;
 wire n_6421;
 wire n_643;
 wire n_6430;
 wire n_6431;
 wire n_6437;
 wire n_6438;
 wire n_6439;
 wire n_644;
 wire n_6444;
 wire n_645;
 wire n_6452;
 wire n_6453;
 wire n_6456;
 wire n_646;
 wire n_6463;
 wire n_647;
 wire n_6471;
 wire n_6474;
 wire n_6476;
 wire n_6477;
 wire n_6478;
 wire n_6479;
 wire n_648;
 wire n_6480;
 wire n_6481;
 wire n_6483;
 wire n_649;
 wire n_650;
 wire n_651;
 wire n_6519;
 wire n_652;
 wire n_6523;
 wire n_6524;
 wire n_6527;
 wire n_6528;
 wire n_653;
 wire n_654;
 wire n_6546;
 wire n_655;
 wire n_656;
 wire n_6569;
 wire n_657;
 wire n_6576;
 wire n_6579;
 wire n_658;
 wire n_6585;
 wire n_6586;
 wire n_6588;
 wire n_6589;
 wire n_659;
 wire n_6591;
 wire n_6592;
 wire n_6593;
 wire n_6599;
 wire n_660;
 wire n_6601;
 wire n_6602;
 wire n_6603;
 wire n_6604;
 wire n_6605;
 wire n_6606;
 wire n_661;
 wire n_6610;
 wire n_6614;
 wire n_6615;
 wire n_6616;
 wire n_6617;
 wire n_6618;
 wire n_6619;
 wire n_662;
 wire n_6620;
 wire n_6635;
 wire n_6639;
 wire n_6646;
 wire n_6655;
 wire n_6656;
 wire n_6657;
 wire n_6658;
 wire n_6660;
 wire n_6661;
 wire n_6666;
 wire n_6667;
 wire n_6668;
 wire n_6669;
 wire n_6673;
 wire n_6675;
 wire n_6676;
 wire n_6687;
 wire n_669;
 wire n_67;
 wire n_670;
 wire n_6710;
 wire n_6724;
 wire n_6727;
 wire n_673;
 wire n_6730;
 wire n_6731;
 wire n_6733;
 wire n_6737;
 wire n_6738;
 wire n_6739;
 wire n_674;
 wire n_6740;
 wire n_6741;
 wire n_6742;
 wire n_6747;
 wire n_6748;
 wire n_6749;
 wire n_675;
 wire n_6751;
 wire n_6753;
 wire n_6754;
 wire n_6758;
 wire n_676;
 wire n_6766;
 wire n_6769;
 wire n_677;
 wire n_6771;
 wire n_6772;
 wire n_6773;
 wire n_6774;
 wire n_678;
 wire n_6783;
 wire n_6784;
 wire n_6787;
 wire n_6788;
 wire n_6789;
 wire n_679;
 wire n_6791;
 wire n_6792;
 wire n_6793;
 wire n_6794;
 wire n_6795;
 wire n_6796;
 wire n_6797;
 wire n_6798;
 wire n_6799;
 wire n_68;
 wire n_680;
 wire n_6806;
 wire n_681;
 wire n_682;
 wire n_6824;
 wire n_6825;
 wire n_683;
 wire n_6830;
 wire n_6832;
 wire n_6833;
 wire n_6836;
 wire n_684;
 wire n_685;
 wire n_6853;
 wire n_686;
 wire n_6861;
 wire n_6862;
 wire n_6866;
 wire n_6871;
 wire n_6872;
 wire n_6877;
 wire n_6878;
 wire n_6879;
 wire n_688;
 wire n_6880;
 wire n_6888;
 wire n_689;
 wire n_6890;
 wire n_6894;
 wire n_6895;
 wire n_6896;
 wire n_690;
 wire n_6902;
 wire n_6903;
 wire n_6904;
 wire n_6905;
 wire n_691;
 wire n_6910;
 wire n_6916;
 wire n_6917;
 wire n_692;
 wire n_6923;
 wire n_6924;
 wire n_6925;
 wire n_6926;
 wire n_6928;
 wire n_6929;
 wire n_693;
 wire n_6930;
 wire n_6932;
 wire n_6935;
 wire n_6936;
 wire n_6937;
 wire n_6938;
 wire n_6939;
 wire n_694;
 wire n_6940;
 wire n_6941;
 wire n_6942;
 wire n_6943;
 wire n_6949;
 wire n_695;
 wire n_6950;
 wire n_6954;
 wire n_6955;
 wire n_6957;
 wire n_6958;
 wire n_696;
 wire n_6960;
 wire n_6961;
 wire n_6962;
 wire n_6963;
 wire n_6964;
 wire n_6965;
 wire n_6967;
 wire n_6968;
 wire n_6969;
 wire n_697;
 wire n_6972;
 wire n_6973;
 wire n_6974;
 wire n_6975;
 wire n_6976;
 wire n_6978;
 wire n_6979;
 wire n_698;
 wire n_6984;
 wire n_6985;
 wire n_6986;
 wire n_6987;
 wire n_6988;
 wire n_6989;
 wire n_699;
 wire n_6991;
 wire n_6992;
 wire n_6993;
 wire n_6994;
 wire n_6995;
 wire n_6996;
 wire n_6997;
 wire n_6999;
 wire n_7;
 wire n_70;
 wire n_700;
 wire n_7000;
 wire n_7006;
 wire n_7007;
 wire n_7008;
 wire n_7009;
 wire n_701;
 wire n_7010;
 wire n_7011;
 wire n_7012;
 wire n_7013;
 wire n_7014;
 wire n_7015;
 wire n_7017;
 wire n_7018;
 wire n_7019;
 wire n_702;
 wire n_7020;
 wire n_7021;
 wire n_7025;
 wire n_7027;
 wire n_7028;
 wire n_7029;
 wire n_703;
 wire n_704;
 wire n_7040;
 wire n_7041;
 wire n_7049;
 wire n_705;
 wire n_7051;
 wire n_7052;
 wire n_7053;
 wire n_706;
 wire n_7060;
 wire n_7061;
 wire n_7062;
 wire n_7063;
 wire n_7064;
 wire n_707;
 wire n_7071;
 wire n_7072;
 wire n_7073;
 wire n_7075;
 wire n_7079;
 wire n_708;
 wire n_7080;
 wire n_7082;
 wire n_709;
 wire n_7096;
 wire n_7097;
 wire n_7098;
 wire n_7099;
 wire n_71;
 wire n_710;
 wire n_7100;
 wire n_7101;
 wire n_7102;
 wire n_7103;
 wire n_7104;
 wire n_7105;
 wire n_7106;
 wire n_7107;
 wire n_7109;
 wire n_711;
 wire n_7111;
 wire n_7116;
 wire n_7117;
 wire n_712;
 wire n_7121;
 wire n_7128;
 wire n_713;
 wire n_714;
 wire n_715;
 wire n_716;
 wire n_7162;
 wire n_7166;
 wire n_7167;
 wire n_7169;
 wire n_717;
 wire n_7170;
 wire n_7171;
 wire n_7172;
 wire n_7179;
 wire n_718;
 wire n_7188;
 wire n_7189;
 wire n_719;
 wire n_7190;
 wire n_7194;
 wire n_7195;
 wire n_7196;
 wire n_7197;
 wire n_7199;
 wire n_72;
 wire n_720;
 wire n_7200;
 wire n_721;
 wire n_7212;
 wire n_7213;
 wire n_7214;
 wire n_7215;
 wire n_722;
 wire n_7222;
 wire n_7223;
 wire n_7227;
 wire n_7228;
 wire n_723;
 wire n_7231;
 wire n_7232;
 wire n_7233;
 wire n_7234;
 wire n_7235;
 wire n_7236;
 wire n_7237;
 wire n_7239;
 wire n_724;
 wire n_7249;
 wire n_725;
 wire n_7250;
 wire n_7255;
 wire n_7256;
 wire n_7257;
 wire n_726;
 wire n_7263;
 wire n_7265;
 wire n_7269;
 wire n_727;
 wire n_728;
 wire n_7282;
 wire n_7283;
 wire n_7284;
 wire n_729;
 wire n_7296;
 wire n_7297;
 wire n_73;
 wire n_730;
 wire n_7307;
 wire n_7309;
 wire n_731;
 wire n_7311;
 wire n_7313;
 wire n_7314;
 wire n_7315;
 wire n_7316;
 wire n_7317;
 wire n_7318;
 wire n_732;
 wire n_7326;
 wire n_7327;
 wire n_7328;
 wire n_733;
 wire n_7330;
 wire n_7332;
 wire n_7333;
 wire n_7334;
 wire n_7335;
 wire n_7336;
 wire n_7338;
 wire n_734;
 wire n_7342;
 wire n_7343;
 wire n_735;
 wire n_7350;
 wire n_7351;
 wire n_7352;
 wire n_7353;
 wire n_7354;
 wire n_7356;
 wire n_736;
 wire n_7360;
 wire n_7361;
 wire n_7362;
 wire n_7363;
 wire n_7364;
 wire n_737;
 wire n_7370;
 wire n_7371;
 wire n_7378;
 wire n_7379;
 wire n_738;
 wire n_7381;
 wire n_7382;
 wire n_7383;
 wire n_7389;
 wire n_739;
 wire n_7390;
 wire n_7394;
 wire n_7397;
 wire n_7399;
 wire n_74;
 wire n_740;
 wire n_7402;
 wire n_7403;
 wire n_7404;
 wire n_7405;
 wire n_7406;
 wire n_7407;
 wire n_7408;
 wire n_7409;
 wire n_741;
 wire n_7410;
 wire n_742;
 wire n_743;
 wire n_7435;
 wire n_744;
 wire n_7447;
 wire n_745;
 wire n_7450;
 wire n_7451;
 wire n_7452;
 wire n_7453;
 wire n_7454;
 wire n_7455;
 wire n_7456;
 wire n_7457;
 wire n_7458;
 wire n_7459;
 wire n_746;
 wire n_7460;
 wire n_7462;
 wire n_7463;
 wire n_7464;
 wire n_7467;
 wire n_7468;
 wire n_7469;
 wire n_747;
 wire n_7470;
 wire n_7471;
 wire n_7473;
 wire n_7474;
 wire n_7476;
 wire n_7477;
 wire n_7478;
 wire n_7479;
 wire n_748;
 wire n_7480;
 wire n_7481;
 wire n_7482;
 wire n_7485;
 wire n_7487;
 wire n_7488;
 wire n_7489;
 wire n_749;
 wire n_7491;
 wire n_7492;
 wire n_7493;
 wire n_7494;
 wire n_7495;
 wire n_7496;
 wire n_7497;
 wire n_750;
 wire n_7502;
 wire n_7506;
 wire n_7507;
 wire n_7508;
 wire n_751;
 wire n_7514;
 wire n_7515;
 wire n_7516;
 wire n_7517;
 wire n_752;
 wire n_7520;
 wire n_7521;
 wire n_7523;
 wire n_7526;
 wire n_7527;
 wire n_753;
 wire n_7531;
 wire n_7534;
 wire n_7536;
 wire n_7537;
 wire n_7538;
 wire n_7539;
 wire n_754;
 wire n_7540;
 wire n_7542;
 wire n_7543;
 wire n_7544;
 wire n_7546;
 wire n_7547;
 wire n_7548;
 wire n_755;
 wire n_7553;
 wire n_7558;
 wire n_756;
 wire n_7565;
 wire n_7566;
 wire n_7568;
 wire n_7569;
 wire n_757;
 wire n_7570;
 wire n_7571;
 wire n_7572;
 wire n_7573;
 wire n_7575;
 wire n_7576;
 wire n_7577;
 wire n_7579;
 wire n_758;
 wire n_7581;
 wire n_7583;
 wire n_7584;
 wire n_7585;
 wire n_7586;
 wire n_7587;
 wire n_7588;
 wire n_7589;
 wire n_759;
 wire n_7590;
 wire n_7591;
 wire n_7592;
 wire n_7593;
 wire n_7595;
 wire n_7596;
 wire n_7597;
 wire n_7598;
 wire n_76;
 wire n_760;
 wire n_7601;
 wire n_7604;
 wire n_7608;
 wire n_7609;
 wire n_761;
 wire n_7610;
 wire n_7612;
 wire n_7615;
 wire n_7618;
 wire n_7619;
 wire n_762;
 wire n_7620;
 wire n_763;
 wire n_7637;
 wire n_7638;
 wire n_764;
 wire n_7644;
 wire n_765;
 wire n_7655;
 wire n_7656;
 wire n_7657;
 wire n_766;
 wire n_7661;
 wire n_7665;
 wire n_7669;
 wire n_767;
 wire n_7670;
 wire n_7675;
 wire n_7676;
 wire n_7677;
 wire n_768;
 wire n_7681;
 wire n_7682;
 wire n_7685;
 wire n_7686;
 wire n_769;
 wire n_7697;
 wire n_7698;
 wire n_77;
 wire n_770;
 wire n_7702;
 wire n_7703;
 wire n_7704;
 wire n_7705;
 wire n_7706;
 wire n_7707;
 wire n_7708;
 wire n_7709;
 wire n_771;
 wire n_7710;
 wire n_7716;
 wire n_7719;
 wire n_772;
 wire n_7720;
 wire n_7721;
 wire n_7724;
 wire n_7726;
 wire n_7727;
 wire n_773;
 wire n_774;
 wire n_7742;
 wire n_7746;
 wire n_7748;
 wire n_7749;
 wire n_775;
 wire n_7753;
 wire n_7754;
 wire n_776;
 wire n_777;
 wire n_7775;
 wire n_7776;
 wire n_7777;
 wire n_7778;
 wire n_7779;
 wire n_778;
 wire n_7780;
 wire n_7781;
 wire n_7782;
 wire n_7783;
 wire n_7784;
 wire n_7786;
 wire n_7787;
 wire n_7788;
 wire n_779;
 wire n_7798;
 wire n_7799;
 wire n_78;
 wire n_780;
 wire n_7800;
 wire n_7801;
 wire n_7803;
 wire n_7804;
 wire n_7805;
 wire n_781;
 wire n_7819;
 wire n_782;
 wire n_7820;
 wire n_7821;
 wire n_783;
 wire n_784;
 wire n_785;
 wire n_7854;
 wire n_7855;
 wire n_7858;
 wire n_7859;
 wire n_786;
 wire n_7862;
 wire n_7863;
 wire n_7868;
 wire n_7869;
 wire n_787;
 wire n_7871;
 wire n_7872;
 wire n_7873;
 wire n_7874;
 wire n_7876;
 wire n_7877;
 wire n_7879;
 wire n_788;
 wire n_7883;
 wire n_7884;
 wire n_7885;
 wire n_7886;
 wire n_789;
 wire n_7893;
 wire n_7894;
 wire n_7898;
 wire n_79;
 wire n_790;
 wire n_7903;
 wire n_7904;
 wire n_7905;
 wire n_7906;
 wire n_7907;
 wire n_7908;
 wire n_7909;
 wire n_791;
 wire n_792;
 wire n_7925;
 wire n_7926;
 wire n_7927;
 wire n_793;
 wire n_7932;
 wire n_7938;
 wire n_794;
 wire n_7947;
 wire n_795;
 wire n_796;
 wire n_7960;
 wire n_7963;
 wire n_7964;
 wire n_7965;
 wire n_797;
 wire n_7970;
 wire n_7971;
 wire n_7972;
 wire n_7973;
 wire n_7974;
 wire n_7979;
 wire n_798;
 wire n_7980;
 wire n_7981;
 wire n_799;
 wire n_7990;
 wire n_7991;
 wire n_7992;
 wire n_7994;
 wire n_7996;
 wire n_7997;
 wire n_7999;
 wire n_80;
 wire n_800;
 wire n_8000;
 wire n_8001;
 wire n_8002;
 wire n_8003;
 wire n_8005;
 wire n_8006;
 wire n_8007;
 wire n_801;
 wire n_8014;
 wire n_8016;
 wire n_8017;
 wire n_8018;
 wire n_8019;
 wire n_802;
 wire n_8022;
 wire n_8027;
 wire n_803;
 wire n_8030;
 wire n_8031;
 wire n_8032;
 wire n_8035;
 wire n_804;
 wire n_805;
 wire n_8053;
 wire n_8057;
 wire n_806;
 wire n_8066;
 wire n_8067;
 wire n_8068;
 wire n_8069;
 wire n_807;
 wire n_8071;
 wire n_8072;
 wire n_808;
 wire n_8088;
 wire n_8089;
 wire n_809;
 wire n_8090;
 wire n_8091;
 wire n_8092;
 wire n_810;
 wire n_8104;
 wire n_8105;
 wire n_8107;
 wire n_8108;
 wire n_8109;
 wire n_811;
 wire n_8115;
 wire n_812;
 wire n_8125;
 wire n_8129;
 wire n_813;
 wire n_8130;
 wire n_8131;
 wire n_8134;
 wire n_8135;
 wire n_8137;
 wire n_814;
 wire n_8140;
 wire n_8141;
 wire n_8144;
 wire n_8145;
 wire n_8146;
 wire n_8148;
 wire n_815;
 wire n_8150;
 wire n_8158;
 wire n_8159;
 wire n_816;
 wire n_8161;
 wire n_8166;
 wire n_8167;
 wire n_817;
 wire n_8170;
 wire n_8174;
 wire n_8175;
 wire n_8176;
 wire n_8178;
 wire n_8180;
 wire n_8185;
 wire n_8187;
 wire n_8188;
 wire n_819;
 wire n_8191;
 wire n_8194;
 wire n_8196;
 wire n_8197;
 wire n_82;
 wire n_820;
 wire n_821;
 wire n_8213;
 wire n_8214;
 wire n_822;
 wire n_8224;
 wire n_8225;
 wire n_8226;
 wire n_8227;
 wire n_8228;
 wire n_823;
 wire n_8232;
 wire n_8233;
 wire n_8235;
 wire n_8237;
 wire n_8238;
 wire n_8239;
 wire n_824;
 wire n_8240;
 wire n_8241;
 wire n_8244;
 wire n_8245;
 wire n_8248;
 wire n_8255;
 wire n_8256;
 wire n_8259;
 wire n_826;
 wire n_8260;
 wire n_8261;
 wire n_8265;
 wire n_827;
 wire n_828;
 wire n_8283;
 wire n_829;
 wire n_8290;
 wire n_8292;
 wire n_8295;
 wire n_8298;
 wire n_8299;
 wire n_83;
 wire n_830;
 wire n_8300;
 wire n_8302;
 wire n_8303;
 wire n_8304;
 wire n_8305;
 wire n_8306;
 wire n_8307;
 wire n_8308;
 wire n_8309;
 wire n_831;
 wire n_8310;
 wire n_8311;
 wire n_8312;
 wire n_8315;
 wire n_832;
 wire n_8320;
 wire n_8321;
 wire n_8322;
 wire n_8323;
 wire n_8324;
 wire n_8325;
 wire n_8326;
 wire n_8329;
 wire n_833;
 wire n_834;
 wire n_8344;
 wire n_8346;
 wire n_8347;
 wire n_8348;
 wire n_8349;
 wire n_835;
 wire n_8351;
 wire n_8352;
 wire n_836;
 wire n_8365;
 wire n_8367;
 wire n_8368;
 wire n_8369;
 wire n_837;
 wire n_8373;
 wire n_8374;
 wire n_8375;
 wire n_8376;
 wire n_8377;
 wire n_8378;
 wire n_838;
 wire n_8380;
 wire n_8387;
 wire n_8388;
 wire n_839;
 wire n_8390;
 wire n_8391;
 wire n_8392;
 wire n_84;
 wire n_840;
 wire n_8406;
 wire n_841;
 wire n_8412;
 wire n_8413;
 wire n_8414;
 wire n_8415;
 wire n_8416;
 wire n_8418;
 wire n_842;
 wire n_8421;
 wire n_8422;
 wire n_8428;
 wire n_843;
 wire n_8436;
 wire n_8437;
 wire n_8438;
 wire n_8439;
 wire n_844;
 wire n_8440;
 wire n_8441;
 wire n_8442;
 wire n_845;
 wire n_846;
 wire n_8461;
 wire n_847;
 wire n_8473;
 wire n_8474;
 wire n_8476;
 wire n_8478;
 wire n_848;
 wire n_8481;
 wire n_8482;
 wire n_8486;
 wire n_8488;
 wire n_8489;
 wire n_849;
 wire n_8490;
 wire n_8492;
 wire n_8494;
 wire n_8495;
 wire n_8496;
 wire n_8497;
 wire n_8498;
 wire n_8499;
 wire n_85;
 wire n_850;
 wire n_8500;
 wire n_8501;
 wire n_8505;
 wire n_8507;
 wire n_851;
 wire n_8512;
 wire n_8519;
 wire n_852;
 wire n_8520;
 wire n_8522;
 wire n_8525;
 wire n_8527;
 wire n_8528;
 wire n_853;
 wire n_8530;
 wire n_8531;
 wire n_8532;
 wire n_854;
 wire n_855;
 wire n_856;
 wire n_8563;
 wire n_8567;
 wire n_8568;
 wire n_857;
 wire n_8572;
 wire n_8573;
 wire n_8575;
 wire n_8576;
 wire n_858;
 wire n_8580;
 wire n_8581;
 wire n_8582;
 wire n_8585;
 wire n_8586;
 wire n_8587;
 wire n_8588;
 wire n_859;
 wire n_8594;
 wire n_8595;
 wire n_8596;
 wire n_860;
 wire n_8605;
 wire n_8606;
 wire n_861;
 wire n_8612;
 wire n_8613;
 wire n_8614;
 wire n_8615;
 wire n_862;
 wire n_8621;
 wire n_8623;
 wire n_8624;
 wire n_8625;
 wire n_8626;
 wire n_8628;
 wire n_8629;
 wire n_863;
 wire n_8631;
 wire n_8637;
 wire n_8638;
 wire n_8639;
 wire n_864;
 wire n_8640;
 wire n_8646;
 wire n_865;
 wire n_8652;
 wire n_8653;
 wire n_8657;
 wire n_8658;
 wire n_866;
 wire n_8660;
 wire n_8661;
 wire n_8662;
 wire n_8663;
 wire n_8665;
 wire n_8666;
 wire n_8667;
 wire n_867;
 wire n_8670;
 wire n_8671;
 wire n_8672;
 wire n_8673;
 wire n_8674;
 wire n_868;
 wire n_8688;
 wire n_8689;
 wire n_869;
 wire n_8690;
 wire n_8691;
 wire n_8694;
 wire n_8696;
 wire n_8697;
 wire n_87;
 wire n_870;
 wire n_8702;
 wire n_871;
 wire n_8719;
 wire n_872;
 wire n_8722;
 wire n_8725;
 wire n_873;
 wire n_8731;
 wire n_8732;
 wire n_8738;
 wire n_8739;
 wire n_874;
 wire n_8747;
 wire n_8748;
 wire n_875;
 wire n_8752;
 wire n_8756;
 wire n_8757;
 wire n_8758;
 wire n_8759;
 wire n_876;
 wire n_8760;
 wire n_8761;
 wire n_8766;
 wire n_8768;
 wire n_877;
 wire n_8770;
 wire n_8771;
 wire n_8772;
 wire n_8773;
 wire n_8776;
 wire n_8777;
 wire n_878;
 wire n_8781;
 wire n_8784;
 wire n_8787;
 wire n_879;
 wire n_8799;
 wire n_88;
 wire n_880;
 wire n_8800;
 wire n_8801;
 wire n_8802;
 wire n_8803;
 wire n_881;
 wire n_882;
 wire n_8821;
 wire n_8823;
 wire n_8826;
 wire n_883;
 wire n_8836;
 wire n_8837;
 wire n_8838;
 wire n_8839;
 wire n_884;
 wire n_8840;
 wire n_8841;
 wire n_8846;
 wire n_8847;
 wire n_8848;
 wire n_8849;
 wire n_885;
 wire n_8850;
 wire n_8851;
 wire n_8852;
 wire n_8853;
 wire n_8855;
 wire n_886;
 wire n_8861;
 wire n_8862;
 wire n_8864;
 wire n_8865;
 wire n_8866;
 wire n_887;
 wire n_8871;
 wire n_8872;
 wire n_8873;
 wire n_8878;
 wire n_888;
 wire n_8881;
 wire n_8882;
 wire n_8886;
 wire n_8888;
 wire n_889;
 wire n_8895;
 wire n_89;
 wire n_890;
 wire n_8901;
 wire n_8902;
 wire n_891;
 wire n_8919;
 wire n_892;
 wire n_8923;
 wire n_8924;
 wire n_8925;
 wire n_8926;
 wire n_8927;
 wire n_8928;
 wire n_8929;
 wire n_893;
 wire n_894;
 wire n_8943;
 wire n_8945;
 wire n_8947;
 wire n_8948;
 wire n_895;
 wire n_8951;
 wire n_8954;
 wire n_8955;
 wire n_8956;
 wire n_8957;
 wire n_8959;
 wire n_896;
 wire n_8962;
 wire n_897;
 wire n_8973;
 wire n_8974;
 wire n_8975;
 wire n_898;
 wire n_8980;
 wire n_8981;
 wire n_8983;
 wire n_8984;
 wire n_8985;
 wire n_8988;
 wire n_8989;
 wire n_899;
 wire n_8990;
 wire n_8991;
 wire n_8992;
 wire n_8993;
 wire n_90;
 wire n_900;
 wire n_9008;
 wire n_9009;
 wire n_901;
 wire n_902;
 wire n_903;
 wire n_9031;
 wire n_9032;
 wire n_9033;
 wire n_9034;
 wire n_9035;
 wire n_9036;
 wire n_9037;
 wire n_9038;
 wire n_904;
 wire n_9041;
 wire n_9042;
 wire n_9048;
 wire n_905;
 wire n_9053;
 wire n_9054;
 wire n_9058;
 wire n_9059;
 wire n_906;
 wire n_9060;
 wire n_9061;
 wire n_9065;
 wire n_9069;
 wire n_907;
 wire n_9070;
 wire n_9074;
 wire n_9076;
 wire n_9077;
 wire n_9078;
 wire n_9079;
 wire n_908;
 wire n_9080;
 wire n_9089;
 wire n_909;
 wire n_9091;
 wire n_9092;
 wire n_9094;
 wire n_91;
 wire n_910;
 wire n_9104;
 wire n_9105;
 wire n_9106;
 wire n_9107;
 wire n_911;
 wire n_9111;
 wire n_912;
 wire n_9120;
 wire n_9123;
 wire n_9124;
 wire n_9125;
 wire n_9126;
 wire n_913;
 wire n_9136;
 wire n_9138;
 wire n_914;
 wire n_9140;
 wire n_9141;
 wire n_9142;
 wire n_9143;
 wire n_915;
 wire n_9154;
 wire n_9155;
 wire n_9156;
 wire n_916;
 wire n_9160;
 wire n_9162;
 wire n_917;
 wire n_9172;
 wire n_9179;
 wire n_918;
 wire n_9180;
 wire n_9181;
 wire n_9182;
 wire n_9183;
 wire n_919;
 wire n_9198;
 wire n_9199;
 wire n_92;
 wire n_920;
 wire n_9200;
 wire n_9201;
 wire n_9202;
 wire n_9206;
 wire n_9209;
 wire n_921;
 wire n_9214;
 wire n_9215;
 wire n_9218;
 wire n_922;
 wire n_923;
 wire n_9231;
 wire n_9234;
 wire n_9235;
 wire n_9237;
 wire n_9238;
 wire n_924;
 wire n_9244;
 wire n_9246;
 wire n_925;
 wire n_9252;
 wire n_9253;
 wire n_9254;
 wire n_9255;
 wire n_9256;
 wire n_9258;
 wire n_9259;
 wire n_926;
 wire n_9261;
 wire n_9263;
 wire n_9267;
 wire n_9269;
 wire n_927;
 wire n_9270;
 wire n_9271;
 wire n_9273;
 wire n_9274;
 wire n_9279;
 wire n_928;
 wire n_9281;
 wire n_929;
 wire n_9292;
 wire n_9293;
 wire n_9295;
 wire n_9296;
 wire n_9297;
 wire n_9298;
 wire n_9299;
 wire n_93;
 wire n_930;
 wire n_9301;
 wire n_9305;
 wire n_931;
 wire n_9313;
 wire n_9316;
 wire n_9317;
 wire n_932;
 wire n_9321;
 wire n_9322;
 wire n_9323;
 wire n_9324;
 wire n_9325;
 wire n_9326;
 wire n_9327;
 wire n_933;
 wire n_9333;
 wire n_9334;
 wire n_9335;
 wire n_9336;
 wire n_9337;
 wire n_9338;
 wire n_9339;
 wire n_934;
 wire n_9340;
 wire n_9341;
 wire n_9342;
 wire n_9344;
 wire n_9349;
 wire n_935;
 wire n_9350;
 wire n_9354;
 wire n_9359;
 wire n_936;
 wire n_9367;
 wire n_9368;
 wire n_937;
 wire n_9370;
 wire n_9373;
 wire n_9375;
 wire n_9376;
 wire n_9379;
 wire n_938;
 wire n_9384;
 wire n_9385;
 wire n_9388;
 wire n_9389;
 wire n_939;
 wire n_9392;
 wire n_94;
 wire n_940;
 wire n_9402;
 wire n_9404;
 wire n_9405;
 wire n_9406;
 wire n_9407;
 wire n_9408;
 wire n_941;
 wire n_9410;
 wire n_9419;
 wire n_942;
 wire n_9420;
 wire n_943;
 wire n_9430;
 wire n_9432;
 wire n_9434;
 wire n_944;
 wire n_9441;
 wire n_9447;
 wire n_9449;
 wire n_945;
 wire n_9450;
 wire n_9451;
 wire n_9452;
 wire n_9453;
 wire n_9455;
 wire n_9456;
 wire n_946;
 wire n_9462;
 wire n_9463;
 wire n_9464;
 wire n_9467;
 wire n_947;
 wire n_9470;
 wire n_9471;
 wire n_9472;
 wire n_9479;
 wire n_948;
 wire n_9480;
 wire n_9481;
 wire n_9483;
 wire n_949;
 wire n_9494;
 wire n_9498;
 wire n_95;
 wire n_950;
 wire n_9501;
 wire n_9503;
 wire n_9506;
 wire n_9507;
 wire n_951;
 wire n_9510;
 wire n_9513;
 wire n_9514;
 wire n_9516;
 wire n_9518;
 wire n_952;
 wire n_9520;
 wire n_9525;
 wire n_953;
 wire n_9534;
 wire n_9535;
 wire n_9536;
 wire n_954;
 wire n_9541;
 wire n_9544;
 wire n_9545;
 wire n_9546;
 wire n_9548;
 wire n_9549;
 wire n_955;
 wire n_956;
 wire n_957;
 wire n_9570;
 wire n_9571;
 wire n_9573;
 wire n_9574;
 wire n_9575;
 wire n_9576;
 wire n_9577;
 wire n_958;
 wire n_9584;
 wire n_959;
 wire n_9591;
 wire n_96;
 wire n_960;
 wire n_9603;
 wire n_9604;
 wire n_9605;
 wire n_961;
 wire n_9614;
 wire n_9616;
 wire n_9617;
 wire n_9618;
 wire n_962;
 wire n_9624;
 wire n_9625;
 wire n_9627;
 wire n_9628;
 wire n_963;
 wire n_9631;
 wire n_9632;
 wire n_9633;
 wire n_9634;
 wire n_9635;
 wire n_9636;
 wire n_9637;
 wire n_9638;
 wire n_9639;
 wire n_964;
 wire n_9642;
 wire n_965;
 wire n_9650;
 wire n_9651;
 wire n_9652;
 wire n_9653;
 wire n_9657;
 wire n_9658;
 wire n_9659;
 wire n_966;
 wire n_9661;
 wire n_9662;
 wire n_9669;
 wire n_967;
 wire n_9671;
 wire n_9672;
 wire n_9675;
 wire n_9677;
 wire n_968;
 wire n_9682;
 wire n_9684;
 wire n_9685;
 wire n_9686;
 wire n_9687;
 wire n_969;
 wire n_9692;
 wire n_9693;
 wire n_9694;
 wire n_9695;
 wire n_9697;
 wire n_9698;
 wire n_970;
 wire n_9700;
 wire n_9704;
 wire n_9708;
 wire n_9709;
 wire n_971;
 wire n_9711;
 wire n_9712;
 wire n_9713;
 wire n_9714;
 wire n_972;
 wire n_9725;
 wire n_9726;
 wire n_9728;
 wire n_973;
 wire n_9735;
 wire n_9739;
 wire n_974;
 wire n_9740;
 wire n_9743;
 wire n_9744;
 wire n_9745;
 wire n_9746;
 wire n_9747;
 wire n_975;
 wire n_9750;
 wire n_9751;
 wire n_9752;
 wire n_9753;
 wire n_9754;
 wire n_9755;
 wire n_9756;
 wire n_9757;
 wire n_9759;
 wire n_976;
 wire n_9762;
 wire n_9763;
 wire n_977;
 wire n_9776;
 wire n_978;
 wire n_979;
 wire n_9792;
 wire n_9793;
 wire n_9794;
 wire n_9795;
 wire n_9797;
 wire n_9799;
 wire n_98;
 wire n_980;
 wire n_9801;
 wire n_9805;
 wire n_9806;
 wire n_9807;
 wire n_9808;
 wire n_981;
 wire n_9810;
 wire n_9811;
 wire n_9813;
 wire n_9818;
 wire n_9819;
 wire n_982;
 wire n_9820;
 wire n_9821;
 wire n_9827;
 wire n_9828;
 wire n_9829;
 wire n_983;
 wire n_9830;
 wire n_9831;
 wire n_9832;
 wire n_9833;
 wire n_984;
 wire n_9840;
 wire n_9841;
 wire n_9842;
 wire n_9848;
 wire n_9849;
 wire n_985;
 wire n_9859;
 wire n_986;
 wire n_9860;
 wire n_9862;
 wire n_9865;
 wire n_9866;
 wire n_987;
 wire n_9874;
 wire n_9879;
 wire n_988;
 wire n_9880;
 wire n_9881;
 wire n_9882;
 wire n_9883;
 wire n_9884;
 wire n_9885;
 wire n_989;
 wire n_9892;
 wire n_9893;
 wire n_9896;
 wire n_9897;
 wire n_9898;
 wire n_9899;
 wire n_99;
 wire n_990;
 wire n_9900;
 wire n_9902;
 wire n_9903;
 wire n_9904;
 wire n_9905;
 wire n_9908;
 wire n_991;
 wire n_9912;
 wire n_9917;
 wire n_992;
 wire n_9922;
 wire n_9923;
 wire n_9925;
 wire n_9926;
 wire n_9927;
 wire n_9928;
 wire n_9929;
 wire n_993;
 wire n_994;
 wire n_995;
 wire n_9950;
 wire n_9956;
 wire n_9957;
 wire n_9959;
 wire n_996;
 wire n_9960;
 wire n_9961;
 wire n_9963;
 wire n_9966;
 wire n_997;
 wire n_9971;
 wire n_9972;
 wire n_9973;
 wire n_9974;
 wire n_9977;
 wire n_9978;
 wire n_998;
 wire n_9985;
 wire n_9986;
 wire n_9987;
 wire n_9988;
 wire n_9989;
 wire n_999;
 wire n_9990;
 wire n_9991;
 wire n_9992;
 wire n_9997;
 wire u_NV_NVDLA_cmac_dp2reg_done;
 wire u_NV_NVDLA_cmac_u_core_in_dat_pvld;
 wire u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1;
 wire u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2;
 wire u_NV_NVDLA_cmac_u_core_in_dat_stripe_end;
 wire u_NV_NVDLA_cmac_u_core_in_dat_stripe_st;
 wire u_NV_NVDLA_cmac_u_core_in_wt_pvld;
 wire u_NV_NVDLA_cmac_u_core_u_active_dat_actv_stripe_end;
 wire u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521;
 wire u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_end_3520;
 wire u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_st_3519;
 wire u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_pvld_3195;
 wire u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_pvld_3196;
 wire u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_pvld_3197;
 wire u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_pvld_3198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_318;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_321;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_322;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_324;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_325;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_327;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_328;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_332;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_336;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_337;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_344;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_345;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_347;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_349;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_352;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_353;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_354;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_356;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_358;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_359;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_360;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_361;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_363;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_366;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_372;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_377;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_379;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_380;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_381;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_383;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_384;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_385;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_386;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_387;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_395;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_396;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_397;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_398;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_401;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_404;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_408;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_421;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_424;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_425;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_429;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_430;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_431;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_432;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_433;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_436;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_437;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_439;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_440;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_443;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_445;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_446;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_448;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_450;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_451;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_453;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_455;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_458;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_462;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_465;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_466;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_472;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_475;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_478;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_480;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_481;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_489;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_500;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_324;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_332;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_306;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_310;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_311;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_310;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_317;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_546;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_547;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_552;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_553;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_559;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_560;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_561;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_562;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_563;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_564;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_565;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_566;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_567;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_568;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_569;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_570;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_571;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_572;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_573;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_574;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_575;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_576;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_577;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_580;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_581;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_582;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_583;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_584;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_585;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_586;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_587;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_591;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_592;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_593;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_594;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_595;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_596;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_597;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_598;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_599;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_600;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_601;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_602;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_603;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_604;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_605;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_610;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_611;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_614;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_615;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_616;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_620;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_621;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_622;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_623;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_624;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_625;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_627;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_629;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_630;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_631;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_632;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_633;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_634;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_635;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_636;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_637;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_638;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_639;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_642;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_648;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_652;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_653;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_654;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_655;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_656;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_657;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_659;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_660;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_661;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_662;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_663;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_664;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_665;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_666;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_667;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_668;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_669;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_670;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_671;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_672;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_673;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_674;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_675;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_680;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_681;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_682;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_683;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_684;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_687;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_688;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_689;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_690;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_691;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_692;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_693;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_694;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_695;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_696;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_697;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_698;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_699;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_700;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_701;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_704;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_705;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_708;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_709;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_712;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_713;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_714;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_716;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_717;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_718;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_720;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_721;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_722;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_723;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_725;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_727;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_728;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_729;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_730;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_731;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_732;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_733;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_736;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_742;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_744;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_745;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_747;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_748;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_750;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_751;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_752;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_753;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_754;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_755;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_756;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_757;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_758;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_759;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_760;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_761;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_762;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_763;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_764;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_765;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_766;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_767;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_768;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_769;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_774;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_776;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_778;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_779;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_782;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_783;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_785;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_786;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_789;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_791;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_792;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_793;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_794;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_795;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_796;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_797;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_798;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_n_799;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_317;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_318;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_322;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_324;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_325;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_327;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_328;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_336;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_337;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_342;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_344;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_345;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_347;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_352;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_353;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_354;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_356;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_358;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_359;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_360;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_361;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_372;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_377;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_379;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_380;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_381;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_383;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_384;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_385;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_386;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_395;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_396;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_397;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_398;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_400;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_401;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_412;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_430;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_431;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_432;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_433;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_437;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_438;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_439;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_443;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_445;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_447;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_449;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_450;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_453;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_455;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_466;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_468;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_472;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_473;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_480;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_481;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_488;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_494;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_496;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_306;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_311;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_310;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_319;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_552;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_554;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_556;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_558;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_559;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_560;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_561;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_562;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_563;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_565;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_567;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_569;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_570;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_571;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_572;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_573;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_574;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_575;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_576;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_578;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_579;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_582;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_583;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_586;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_588;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_589;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_592;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_594;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_595;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_596;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_597;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_598;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_599;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_600;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_601;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_602;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_603;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_604;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_605;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_608;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_609;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_616;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_617;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_618;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_619;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_620;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_622;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_623;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_624;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_625;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_626;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_627;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_628;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_629;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_630;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_631;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_632;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_633;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_634;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_635;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_636;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_637;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_638;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_639;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_642;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_643;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_648;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_649;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_650;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_651;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_652;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_654;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_655;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_656;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_658;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_659;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_660;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_661;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_662;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_663;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_664;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_665;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_666;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_667;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_668;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_669;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_670;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_671;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_672;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_674;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_678;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_680;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_682;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_683;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_684;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_685;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_686;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_687;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_688;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_690;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_691;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_692;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_693;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_694;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_695;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_697;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_698;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_699;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_700;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_701;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_708;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_709;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_716;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_718;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_720;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_721;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_722;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_723;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_725;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_728;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_729;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_730;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_731;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_732;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_733;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_737;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_739;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_740;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_743;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_746;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_748;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_750;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_751;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_752;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_753;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_754;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_755;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_756;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_757;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_758;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_759;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_760;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_761;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_762;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_763;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_764;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_765;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_766;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_767;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_770;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_776;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_778;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_780;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_782;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_783;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_785;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_786;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_787;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_788;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_789;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_790;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_791;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_792;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_793;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_794;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_795;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_796;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_797;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_798;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_n_799;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_316;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_317;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_318;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_319;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_320;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_321;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_322;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_324;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_325;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_327;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_328;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_331;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_332;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_336;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_337;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_343;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_344;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_345;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_346;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_347;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_349;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_352;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_354;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_356;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_357;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_358;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_359;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_361;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_362;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_372;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_373;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_375;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_379;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_380;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_381;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_384;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_387;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_395;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_396;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_397;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_398;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_399;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_401;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_412;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_424;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_429;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_430;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_431;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_432;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_433;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_438;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_439;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_445;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_448;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_450;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_451;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_453;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_455;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_465;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_481;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_490;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_500;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_310;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_317;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_289;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_318;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_319;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_552;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_553;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_554;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_556;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_558;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_559;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_560;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_561;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_562;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_565;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_566;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_567;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_568;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_569;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_570;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_571;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_572;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_573;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_574;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_575;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_576;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_580;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_581;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_582;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_584;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_585;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_588;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_591;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_594;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_595;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_596;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_597;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_598;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_599;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_600;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_601;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_602;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_603;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_604;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_605;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_610;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_613;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_620;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_621;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_622;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_623;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_624;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_625;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_627;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_628;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_630;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_631;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_632;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_633;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_634;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_635;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_636;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_637;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_638;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_639;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_643;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_644;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_645;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_646;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_647;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_648;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_650;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_651;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_652;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_653;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_655;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_656;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_657;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_659;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_660;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_662;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_663;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_664;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_665;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_666;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_667;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_668;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_669;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_670;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_671;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_672;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_673;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_674;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_676;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_677;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_678;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_680;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_681;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_684;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_687;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_690;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_691;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_692;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_693;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_695;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_696;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_697;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_698;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_699;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_700;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_701;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_705;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_708;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_712;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_713;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_714;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_716;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_717;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_718;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_719;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_720;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_722;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_723;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_724;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_725;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_726;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_727;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_728;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_729;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_730;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_731;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_732;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_733;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_736;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_737;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_738;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_739;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_740;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_742;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_744;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_745;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_746;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_748;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_750;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_751;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_752;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_753;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_754;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_755;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_757;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_759;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_760;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_761;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_762;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_763;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_764;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_765;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_766;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_767;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_776;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_777;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_778;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_783;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_785;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_788;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_789;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_790;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_791;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_792;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_793;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_794;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_795;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_796;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_797;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_798;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_n_799;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_187;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_203;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_272;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_308;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_311;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_315;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_317;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_321;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_322;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_324;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_325;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_326;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_327;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_329;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_336;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_337;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_34;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_340;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_343;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_344;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_345;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_350;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_352;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_354;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_356;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_357;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_358;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_359;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_361;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_362;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_366;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_372;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_379;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_380;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_381;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_384;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_391;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_396;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_397;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_398;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_400;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_401;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_404;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_406;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_407;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_408;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_417;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_418;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_429;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_430;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_432;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_435;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_436;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_437;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_439;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_440;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_442;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_444;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_445;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_446;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_450;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_451;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_452;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_453;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_455;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_465;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_466;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_473;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_480;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_481;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_483;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_488;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_494;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_500;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_109;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_165;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_204;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_27;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_156;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_25;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_281;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_283;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_284;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_307;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_316;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_331;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_161;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_189;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_218;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_232;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_235;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_256;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_270;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_126;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_13;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_16;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_192;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_196;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_206;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_216;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_227;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_28;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_5;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_69;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_127;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_136;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_155;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_188;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_215;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_253;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_291;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_312;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_39;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_42;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_81;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_103;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_104;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_108;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_117;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_123;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_147;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_162;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_17;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_191;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_21;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_219;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_220;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_221;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_231;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_234;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_24;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_263;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_276;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_277;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_287;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_288;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_299;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_3;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_310;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_314;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_319;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_32;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_33;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_4;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_41;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_49;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_52;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_87;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_10;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_100;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_101;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_102;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_106;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_11;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_111;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_113;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_114;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_115;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_132;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_135;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_14;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_140;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_144;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_145;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_148;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_15;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_150;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_154;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_164;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_166;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_18;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_185;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_186;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_19;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_195;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_197;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_20;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_202;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_207;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_217;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_223;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_224;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_226;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_233;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_236;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_241;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_242;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_243;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_246;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_254;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_257;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_259;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_261;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_262;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_267;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_268;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_269;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_273;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_274;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_280;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_290;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_295;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_296;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_297;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_300;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_303;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_305;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_306;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_31;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_313;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_35;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_36;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_38;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_44;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_45;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_51;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_55;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_56;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_60;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_61;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_63;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_65;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_68;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_70;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_72;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_77;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_78;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_82;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_89;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_91;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_92;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_93;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_94;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_96;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_97;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_0;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_105;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_107;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_110;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_112;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_116;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_119;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_12;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_120;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_121;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_122;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_124;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_125;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_128;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_129;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_130;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_131;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_133;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_134;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_137;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_138;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_139;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_141;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_142;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_143;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_146;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_149;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_151;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_152;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_153;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_157;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_158;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_159;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_160;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_163;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_167;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_168;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_169;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_170;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_179;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_180;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_183;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_190;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_193;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_194;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_198;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_199;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_2;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_200;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_201;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_205;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_208;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_209;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_210;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_211;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_212;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_213;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_214;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_22;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_222;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_225;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_228;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_229;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_23;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_230;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_237;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_238;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_239;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_240;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_244;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_245;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_247;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_248;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_249;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_250;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_251;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_255;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_258;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_26;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_260;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_264;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_265;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_266;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_271;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_275;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_278;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_279;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_282;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_285;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_286;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_29;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_292;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_293;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_294;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_298;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_301;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_304;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_309;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_330;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_37;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_40;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_43;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_46;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_47;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_48;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_50;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_53;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_54;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_57;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_58;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_59;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_6;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_62;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_64;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_66;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_67;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_7;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_71;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_73;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_74;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_75;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_76;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_79;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_8;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_80;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_83;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_84;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_85;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_86;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_88;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_9;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_90;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_95;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_98;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_99;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_171;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_172;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_173;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_174;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_175;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_176;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_177;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_178;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_181;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_182;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_184;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_544;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_545;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_546;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_549;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_552;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_553;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_559;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_562;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_564;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_565;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_566;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_567;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_568;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_569;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_570;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_571;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_572;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_573;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_574;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_575;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_583;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_584;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_586;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_587;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_590;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_591;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_592;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_593;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_594;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_595;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_596;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_597;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_598;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_599;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_600;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_601;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_602;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_603;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_604;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_605;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_610;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_616;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_618;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_619;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_620;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_621;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_622;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_624;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_625;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_627;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_628;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_629;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_630;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_631;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_632;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_633;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_634;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_635;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_636;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_637;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_638;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_639;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_643;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_646;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_647;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_648;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_651;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_652;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_653;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_654;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_655;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_656;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_657;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_658;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_659;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_660;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_661;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_662;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_663;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_664;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_665;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_666;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_667;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_668;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_669;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_670;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_671;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_674;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_676;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_680;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_682;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_683;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_686;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_687;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_688;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_689;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_690;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_691;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_692;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_693;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_694;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_695;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_696;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_697;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_698;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_699;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_700;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_701;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_709;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_711;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_712;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_713;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_714;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_716;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_718;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_719;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_720;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_722;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_723;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_724;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_725;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_726;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_727;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_728;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_729;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_730;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_731;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_732;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_733;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_737;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_738;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_739;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_740;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_743;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_744;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_746;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_748;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_751;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_752;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_753;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_755;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_757;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_758;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_759;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_760;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_761;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_762;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_763;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_764;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_765;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_766;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_767;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_776;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_777;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_778;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_779;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_780;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_783;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_784;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_786;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_788;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_789;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_790;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_791;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_792;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_793;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_794;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_795;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_796;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_797;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_798;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_n_799;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1;
 wire u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2;
 wire u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1;
 wire u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1;
 wire u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d1;
 wire u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d2;
 wire u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1;
 wire u_NV_NVDLA_cmac_u_reg_dp2reg_consumer;
 wire u_NV_NVDLA_cmac_u_reg_n_1228_BAR;
 wire u_NV_NVDLA_cmac_u_reg_n_1258;
 wire u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en;
 wire u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en;
 wire u_NV_NVDLA_cmac_u_reg_reg2dp_producer;
 wire u_NV_NVDLA_cmac_u_reg_req_pvld;
 wire u_partition_m_reset_sync_reset_synced_rstn_NV_GENERIC_CELL_d0;
 wire u_partition_m_reset_sync_reset_synced_rstn_reset_;
 wire [63:0] u_NV_NVDLA_cmac_u_core_dat0_actv_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_dat0_actv_nz;
 wire [7:0] u_NV_NVDLA_cmac_u_core_dat0_actv_pvld;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data0;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data2;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data3;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data4;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data5;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data6;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_data7;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_dat_mask;
 wire [8:0] u_NV_NVDLA_cmac_u_core_in_dat_pd_d1;
 wire [8:0] u_NV_NVDLA_cmac_u_core_in_dat_pd_d2;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data0;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data2;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data3;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data4;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data5;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data6;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_data7;
 wire [7:0] u_NV_NVDLA_cmac_u_core_in_wt_mask;
 wire [3:0] u_NV_NVDLA_cmac_u_core_in_wt_sel;
 wire [18:0] u_NV_NVDLA_cmac_u_core_out_data0;
 wire [18:0] u_NV_NVDLA_cmac_u_core_out_data1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_out_data2;
 wire [18:0] u_NV_NVDLA_cmac_u_core_out_data3;
 wire [3:0] u_NV_NVDLA_cmac_u_core_out_mask;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz;
 wire [63:0] u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz;
 wire [3:0] u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1;
 wire [8:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1;
 wire [8:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1;
 wire [7:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1;
 wire [3:0] u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1;
 wire [18:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1;
 wire [3:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1;
 wire [8:0] u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1;
 wire [63:0] u_NV_NVDLA_cmac_u_core_wt0_actv_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt0_actv_nz;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt0_actv_pvld;
 wire [63:0] u_NV_NVDLA_cmac_u_core_wt1_actv_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt1_actv_nz;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt1_actv_pvld;
 wire [63:0] u_NV_NVDLA_cmac_u_core_wt2_actv_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt2_actv_nz;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt2_actv_pvld;
 wire [63:0] u_NV_NVDLA_cmac_u_core_wt3_actv_data;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt3_actv_nz;
 wire [7:0] u_NV_NVDLA_cmac_u_core_wt3_actv_pvld;
 wire [55:0] u_NV_NVDLA_cmac_u_reg_req_pd;
 wire [13:0] u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out;
 wire [13:0] u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out;

 HB1xp67_ASAP7_75t_SL fopt (.A(n_2588),
    .Y(n_26264));
 INVx1_ASAP7_75t_SL fopt1 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_152),
    .Y(n_12111));
 BUFx6f_ASAP7_75t_SL fopt10 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[2]),
    .Y(n_21183));
 INVxp67_ASAP7_75t_SL fopt101 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_0),
    .Y(n_10745));
 INVxp67_ASAP7_75t_SL fopt102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_74),
    .Y(n_22024));
 INVx1_ASAP7_75t_SL fopt103 (.A(n_22025),
    .Y(n_22026));
 INVx2_ASAP7_75t_SL fopt106 (.A(n_7710),
    .Y(n_23087));
 HB1xp67_ASAP7_75t_SL fopt1066 (.A(n_19495),
    .Y(n_12498));
 INVxp67_ASAP7_75t_SL fopt1067 (.A(n_21577),
    .Y(n_12513));
 HB1xp67_ASAP7_75t_SL fopt107 (.A(n_13123),
    .Y(n_13124));
 HB1xp67_ASAP7_75t_SL fopt109 (.A(n_14808),
    .Y(n_14810));
 INVx1_ASAP7_75t_SL fopt113 (.A(n_5894),
    .Y(n_5895));
 INVxp67_ASAP7_75t_SL fopt115 (.A(n_22519),
    .Y(n_11791));
 INVx2_ASAP7_75t_SL fopt116 (.A(n_22519),
    .Y(n_11787));
 INVx2_ASAP7_75t_SL fopt118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .Y(n_8053));
 INVx3_ASAP7_75t_SL fopt12 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[36]),
    .Y(n_22742));
 INVx1_ASAP7_75t_SL fopt125 (.A(n_19386),
    .Y(n_19387));
 INVx2_ASAP7_75t_SL fopt128 (.A(n_9138),
    .Y(n_11346));
 INVx1_ASAP7_75t_SL fopt1289 (.A(n_11583),
    .Y(n_11586));
 INVxp67_ASAP7_75t_SL fopt129 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_80),
    .Y(n_8895));
 INVxp67_ASAP7_75t_SL fopt1291 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_268),
    .Y(n_11568));
 INVx3_ASAP7_75t_SL fopt13 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[28]),
    .Y(n_14986));
 HB1xp67_ASAP7_75t_SL fopt13271 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_342),
    .Y(n_2271));
 HB1xp67_ASAP7_75t_SL fopt13273 (.A(n_13589),
    .Y(n_2275));
 HB1xp67_ASAP7_75t_SL fopt13274 (.A(n_21974),
    .Y(n_2277));
 HB1xp67_ASAP7_75t_SL fopt13277 (.A(n_8614),
    .Y(n_2283));
 HB1xp67_ASAP7_75t_SL fopt13282 (.A(n_22247),
    .Y(n_2312));
 INVxp67_ASAP7_75t_SL fopt13290 (.A(n_2325),
    .Y(n_2331));
 BUFx6f_ASAP7_75t_SL fopt13291 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[4]),
    .Y(n_2325));
 INVx2_ASAP7_75t_SL fopt13292 (.A(n_2339),
    .Y(n_2335));
 INVx2_ASAP7_75t_SL fopt13293 (.A(n_2339),
    .Y(n_2337));
 INVx2_ASAP7_75t_SL fopt13294 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[4]),
    .Y(n_2339));
 HB1xp67_ASAP7_75t_SL fopt133 (.A(n_20093),
    .Y(n_11071));
 INVxp67_ASAP7_75t_SL fopt13308 (.A(n_2364),
    .Y(n_2366));
 BUFx2_ASAP7_75t_L fopt13311 (.A(n_2359),
    .Y(n_2364));
 BUFx6f_ASAP7_75t_SL fopt13315 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(n_2359));
 BUFx3_ASAP7_75t_SL fopt13316 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(n_2377));
 INVxp67_ASAP7_75t_SL fopt13318 (.A(n_2381),
    .Y(n_2384));
 BUFx3_ASAP7_75t_SL fopt13322 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(n_2381));
 BUFx3_ASAP7_75t_SL fopt13323 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(n_2392));
 HB1xp67_ASAP7_75t_SL fopt13325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_37),
    .Y(n_2400));
 HB1xp67_ASAP7_75t_SL fopt13342 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_343),
    .Y(n_2429));
 HB1xp67_ASAP7_75t_SL fopt13343 (.A(n_21511),
    .Y(n_2431));
 HB1xp67_ASAP7_75t_SL fopt13345 (.A(n_22892),
    .Y(n_2435));
 HB1xp67_ASAP7_75t_SL fopt13347 (.A(n_24201),
    .Y(n_2439));
 INVx1_ASAP7_75t_SL fopt13348 (.A(n_2442),
    .Y(n_2441));
 INVx1_ASAP7_75t_SL fopt13350 (.A(n_2445),
    .Y(n_2444));
 INVxp67_ASAP7_75t_SL fopt13355 (.A(n_2466),
    .Y(n_2465));
 BUFx6f_ASAP7_75t_SL fopt13357 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(n_2466));
 INVxp67_ASAP7_75t_SL fopt13372 (.A(n_2499),
    .Y(n_2507));
 BUFx3_ASAP7_75t_SL fopt13373 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(n_2499));
 INVxp67_ASAP7_75t_SL fopt13375 (.A(n_2525),
    .Y(n_2524));
 HB1xp67_ASAP7_75t_SL fopt13380 (.A(n_5737),
    .Y(n_2525));
 INVxp67_ASAP7_75t_SL fopt13393 (.A(n_2544),
    .Y(n_2552));
 BUFx6f_ASAP7_75t_SL fopt13399 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(n_2544));
 INVxp67_ASAP7_75t_SL fopt13400 (.A(n_2564),
    .Y(n_2562));
 HB1xp67_ASAP7_75t_SL fopt13402 (.A(n_9494),
    .Y(n_2564));
 HB1xp67_ASAP7_75t_SL fopt13403 (.A(n_21646),
    .Y(n_2566));
 HB1xp67_ASAP7_75t_SL fopt13412 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .Y(n_2578));
 INVxp67_ASAP7_75t_SL fopt13417 (.A(n_2580),
    .Y(n_2582));
 INVx2_ASAP7_75t_SL fopt13419 (.A(n_26202),
    .Y(n_2580));
 INVxp67_ASAP7_75t_SL fopt13425 (.A(n_2591),
    .Y(n_2592));
 INVxp67_ASAP7_75t_SL fopt13427 (.A(n_8768),
    .Y(n_2591));
 HB1xp67_ASAP7_75t_SL fopt13437 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .Y(n_2620));
 HB1xp67_ASAP7_75t_SL fopt13451 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_37),
    .Y(n_2642));
 HB1xp67_ASAP7_75t_SL fopt13458 (.A(n_12959),
    .Y(n_2663));
 INVx1_ASAP7_75t_SL fopt13464 (.A(n_19342),
    .Y(n_2673));
 BUFx3_ASAP7_75t_SL fopt13468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_103),
    .Y(n_2685));
 HB1xp67_ASAP7_75t_SL fopt13469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_31),
    .Y(n_2686));
 HB1xp67_ASAP7_75t_SL fopt13471 (.A(n_17474),
    .Y(n_2689));
 HB1xp67_ASAP7_75t_SL fopt13474 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_31),
    .Y(n_2694));
 INVxp67_ASAP7_75t_SL fopt13476 (.A(n_2697),
    .Y(n_2700));
 BUFx3_ASAP7_75t_SL fopt13480 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(n_2697));
 BUFx3_ASAP7_75t_SL fopt13481 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(n_2711));
 BUFx3_ASAP7_75t_SL fopt13488 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_2728));
 HB1xp67_ASAP7_75t_SL fopt13492 (.A(n_12663),
    .Y(n_2735));
 INVx1_ASAP7_75t_SL fopt13496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .Y(n_2741));
 HB1xp67_ASAP7_75t_SL fopt13498 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_27),
    .Y(n_2744));
 INVx1_ASAP7_75t_SL fopt135 (.A(n_18842),
    .Y(n_8766));
 INVxp67_ASAP7_75t_SL fopt13501 (.A(n_2746),
    .Y(n_2747));
 BUFx3_ASAP7_75t_SL fopt13503 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(n_2746));
 HB1xp67_ASAP7_75t_SL fopt13504 (.A(n_20870),
    .Y(n_2764));
 INVxp67_ASAP7_75t_SL fopt13505 (.A(n_6965),
    .Y(n_2766));
 HB1xp67_ASAP7_75t_SL fopt13511 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_31),
    .Y(n_2781));
 HB1xp67_ASAP7_75t_SL fopt13513 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_31),
    .Y(n_2785));
 HB1xp67_ASAP7_75t_SL fopt13515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_31),
    .Y(n_2789));
 HB1xp67_ASAP7_75t_SL fopt13517 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_31),
    .Y(n_2793));
 HB1xp67_ASAP7_75t_SL fopt13521 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_31),
    .Y(n_2801));
 HB1xp67_ASAP7_75t_SL fopt13523 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_31),
    .Y(n_2805));
 INVxp33_ASAP7_75t_SRAM fopt13527 (.A(n_2820),
    .Y(n_2821));
 BUFx3_ASAP7_75t_SL fopt13528 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[60]),
    .Y(n_2820));
 BUFx6f_ASAP7_75t_SL fopt13529 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[60]),
    .Y(n_2825));
 INVx2_ASAP7_75t_SL fopt13535 (.A(n_2836),
    .Y(n_2831));
 INVxp67_ASAP7_75t_SL fopt13537 (.A(n_2827),
    .Y(n_2841));
 BUFx6f_ASAP7_75t_SL fopt13539 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(n_2827));
 HB1xp67_ASAP7_75t_SL fopt13540 (.A(n_24754),
    .Y(n_2848));
 INVxp67_ASAP7_75t_SL fopt13541 (.A(n_2852),
    .Y(n_2850));
 INVx5_ASAP7_75t_SL fopt13545 (.A(n_21185),
    .Y(n_2855));
 INVxp67_ASAP7_75t_SL fopt13548 (.A(n_2864),
    .Y(n_2865));
 INVx3_ASAP7_75t_SL fopt13549 (.A(n_21185),
    .Y(n_2864));
 HB1xp67_ASAP7_75t_SL fopt13554 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_177),
    .Y(n_2873));
 HB1xp67_ASAP7_75t_SL fopt13556 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_177),
    .Y(n_2877));
 HB1xp67_ASAP7_75t_SL fopt13559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_37),
    .Y(n_2883));
 HB1xp67_ASAP7_75t_SL fopt13561 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_37),
    .Y(n_2887));
 HB1xp67_ASAP7_75t_SL fopt13563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_177),
    .Y(n_2891));
 HB1xp67_ASAP7_75t_SL fopt13564 (.A(n_9252),
    .Y(n_2893));
 HB1xp67_ASAP7_75t_SL fopt13566 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_292),
    .Y(n_2897));
 HB1xp67_ASAP7_75t_SL fopt13568 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_292),
    .Y(n_2901));
 HB1xp67_ASAP7_75t_SL fopt13569 (.A(n_10501),
    .Y(n_2903));
 BUFx6f_ASAP7_75t_SL fopt13573 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[52]),
    .Y(n_2922));
 BUFx6f_ASAP7_75t_SL fopt13574 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[52]),
    .Y(n_2927));
 INVx1_ASAP7_75t_SL fopt13575 (.A(n_13423),
    .Y(n_2930));
 INVxp67_ASAP7_75t_SL fopt13577 (.A(n_2927),
    .Y(n_2934));
 INVxp33_ASAP7_75t_SL fopt13580 (.A(n_22463),
    .Y(n_2939));
 INVx1_ASAP7_75t_SL fopt13581 (.A(n_22463),
    .Y(n_2940));
 INVx1_ASAP7_75t_SL fopt13585 (.A(n_2943),
    .Y(n_2945));
 INVxp67_ASAP7_75t_SL fopt13586 (.A(n_2944),
    .Y(n_2943));
 BUFx3_ASAP7_75t_SL fopt13588 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(n_2944));
 HB1xp67_ASAP7_75t_SL fopt13589 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(n_2958));
 INVxp67_ASAP7_75t_SL fopt13590 (.A(n_22735),
    .Y(n_2962));
 INVxp67_ASAP7_75t_SL fopt13592 (.A(n_9682),
    .Y(n_2965));
 INVx1_ASAP7_75t_SL fopt13593 (.A(n_9682),
    .Y(n_2966));
 INVx2_ASAP7_75t_SL fopt13600 (.A(n_22615),
    .Y(n_2985));
 INVx2_ASAP7_75t_SL fopt13602 (.A(n_22615),
    .Y(n_2990));
 HB1xp67_ASAP7_75t_SL fopt13613 (.A(n_10159),
    .Y(n_3011));
 HB1xp67_ASAP7_75t_SL fopt13620 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_36),
    .Y(n_3030));
 HB1xp67_ASAP7_75t_SL fopt13621 (.A(n_21340),
    .Y(n_3032));
 BUFx3_ASAP7_75t_SL fopt13640 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_103),
    .Y(n_3090));
 INVx4_ASAP7_75t_SL fopt13644 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(n_3107));
 INVxp67_ASAP7_75t_SL fopt13660 (.A(n_3150),
    .Y(n_3149));
 HB1xp67_ASAP7_75t_SL fopt13662 (.A(n_3148),
    .Y(n_3150));
 BUFx6f_ASAP7_75t_SL fopt13672 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(n_3148));
 INVxp67_ASAP7_75t_SL fopt13674 (.A(n_3168),
    .Y(n_3170));
 BUFx3_ASAP7_75t_SL fopt13677 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(n_3168));
 BUFx3_ASAP7_75t_SL fopt13678 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(n_3181));
 INVxp67_ASAP7_75t_SL fopt13681 (.A(n_22879),
    .Y(n_3190));
 HB1xp67_ASAP7_75t_SL fopt13687 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_27),
    .Y(n_3204));
 HB1xp67_ASAP7_75t_SL fopt13689 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .Y(n_3208));
 INVxp67_ASAP7_75t_SL fopt13690 (.A(n_19041),
    .Y(n_3210));
 HB1xp67_ASAP7_75t_SL fopt13691 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .Y(n_3212));
 BUFx6f_ASAP7_75t_SL fopt13692 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[34]),
    .Y(n_3214));
 INVxp67_ASAP7_75t_SL fopt13693 (.A(n_3218),
    .Y(n_3224));
 BUFx6f_ASAP7_75t_SL fopt13694 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[34]),
    .Y(n_3218));
 INVxp67_ASAP7_75t_SL fopt13695 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_131),
    .Y(n_3229));
 HB1xp67_ASAP7_75t_SL fopt13696 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .Y(n_3231));
 INVxp67_ASAP7_75t_SL fopt13697 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_131),
    .Y(n_3233));
 HB1xp67_ASAP7_75t_SL fopt13699 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .Y(n_3237));
 INVxp67_ASAP7_75t_SL fopt13700 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_131),
    .Y(n_3239));
 INVxp67_ASAP7_75t_SL fopt13702 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_226),
    .Y(n_3243));
 INVxp67_ASAP7_75t_SL fopt13704 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_275),
    .Y(n_3246));
 BUFx3_ASAP7_75t_SL fopt13711 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(n_3260));
 INVxp67_ASAP7_75t_SL fopt13712 (.A(n_3266),
    .Y(n_3265));
 BUFx3_ASAP7_75t_SL fopt13718 (.A(n_3275),
    .Y(n_3266));
 BUFx6f_ASAP7_75t_SL fopt13719 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(n_3275));
 INVxp67_ASAP7_75t_SL fopt13733 (.A(n_3309),
    .Y(n_3314));
 BUFx6f_ASAP7_75t_SL fopt13734 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[42]),
    .Y(n_3309));
 BUFx6f_ASAP7_75t_SL fopt13735 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[42]),
    .Y(n_3317));
 INVxp67_ASAP7_75t_SL fopt13736 (.A(n_3331),
    .Y(n_3332));
 BUFx3_ASAP7_75t_SL fopt13737 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(n_3331));
 HB1xp67_ASAP7_75t_SL fopt13750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_9),
    .Y(n_3358));
 HB1xp67_ASAP7_75t_SL fopt13751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_9),
    .Y(n_3360));
 HB1xp67_ASAP7_75t_SL fopt13753 (.A(n_9677),
    .Y(n_3364));
 INVxp67_ASAP7_75t_SL fopt13754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_129),
    .Y(n_3366));
 INVxp67_ASAP7_75t_SL fopt13756 (.A(n_3375),
    .Y(n_3376));
 BUFx3_ASAP7_75t_SL fopt13757 (.A(n_3374),
    .Y(n_3375));
 BUFx3_ASAP7_75t_SL fopt13758 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(n_3374));
 INVxp67_ASAP7_75t_SL fopt13761 (.A(n_3396),
    .Y(n_3398));
 BUFx3_ASAP7_75t_SL fopt13764 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(n_3396));
 INVxp67_ASAP7_75t_SL fopt13765 (.A(n_3408),
    .Y(n_3409));
 BUFx3_ASAP7_75t_SL fopt13766 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(n_3408));
 INVxp67_ASAP7_75t_SL fopt13769 (.A(n_12800),
    .Y(n_3433));
 HB1xp67_ASAP7_75t_SL fopt13771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_31),
    .Y(n_3436));
 HB1xp67_ASAP7_75t_SL fopt13775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_142),
    .Y(n_3443));
 HB1xp67_ASAP7_75t_SL fopt13776 (.A(n_22172),
    .Y(n_3445));
 HB1xp67_ASAP7_75t_SL fopt13781 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_31),
    .Y(n_3454));
 HB1xp67_ASAP7_75t_SL fopt13782 (.A(n_3457),
    .Y(n_3456));
 INVx1_ASAP7_75t_SL fopt13783 (.A(n_26077),
    .Y(n_3457));
 HB1xp67_ASAP7_75t_SL fopt13784 (.A(n_8582),
    .Y(n_3459));
 HB1xp67_ASAP7_75t_SL fopt13786 (.A(n_19820),
    .Y(n_3463));
 INVxp67_ASAP7_75t_SRAM fopt13789 (.A(n_3468),
    .Y(n_3469));
 BUFx3_ASAP7_75t_SL fopt13790 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[51]),
    .Y(n_3468));
 BUFx6f_ASAP7_75t_SL fopt13792 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[51]),
    .Y(n_3474));
 BUFx6f_ASAP7_75t_SL fopt13794 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[51]),
    .Y(n_3479));
 INVxp67_ASAP7_75t_SL fopt13798 (.A(n_3491),
    .Y(n_3493));
 HB1xp67_ASAP7_75t_SL fopt138 (.A(n_20716),
    .Y(n_20721));
 BUFx3_ASAP7_75t_SL fopt13800 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(n_3491));
 BUFx3_ASAP7_75t_SL fopt13801 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(n_3504));
 INVx2_ASAP7_75t_SL fopt13803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_226),
    .Y(n_3511));
 INVx2_ASAP7_75t_SL fopt13806 (.A(n_26167),
    .Y(n_3516));
 INVxp67_ASAP7_75t_SL fopt13809 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_226),
    .Y(n_3521));
 INVx1_ASAP7_75t_SL fopt13810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_226),
    .Y(n_3522));
 INVxp67_ASAP7_75t_SL fopt13813 (.A(n_3528),
    .Y(n_3527));
 BUFx6f_ASAP7_75t_SL fopt13814 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .Y(n_3528));
 HB1xp67_ASAP7_75t_SL fopt13821 (.A(n_3548),
    .Y(n_3547));
 INVx1_ASAP7_75t_SL fopt13822 (.A(n_9042),
    .Y(n_3548));
 BUFx2_ASAP7_75t_SL fopt13824 (.A(n_3553),
    .Y(n_3552));
 INVx1_ASAP7_75t_SL fopt13825 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_222),
    .Y(n_3553));
 HB1xp67_ASAP7_75t_SL fopt13827 (.A(n_3558),
    .Y(n_3557));
 INVx1_ASAP7_75t_SL fopt13828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_222),
    .Y(n_3558));
 HB1xp67_ASAP7_75t_SL fopt13829 (.A(n_11384),
    .Y(n_3560));
 HB1xp67_ASAP7_75t_SL fopt13830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_150),
    .Y(n_3562));
 INVxp67_ASAP7_75t_SL fopt13844 (.A(n_3592),
    .Y(n_3593));
 BUFx3_ASAP7_75t_SL fopt13845 (.A(n_3591),
    .Y(n_3592));
 BUFx6f_ASAP7_75t_SL fopt13846 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(n_3591));
 HB1xp67_ASAP7_75t_SL fopt13853 (.A(n_15176),
    .Y(n_3619));
 INVxp67_ASAP7_75t_SL fopt13858 (.A(n_3630),
    .Y(n_3633));
 BUFx3_ASAP7_75t_SL fopt13864 (.A(n_19411),
    .Y(n_3630));
 HB1xp67_ASAP7_75t_SL fopt13866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_29),
    .Y(n_3642));
 INVx1_ASAP7_75t_SL fopt13867 (.A(n_3645),
    .Y(n_3644));
 HB1xp67_ASAP7_75t_SL fopt13868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .Y(n_3645));
 HB1xp67_ASAP7_75t_SL fopt13869 (.A(n_23069),
    .Y(n_3647));
 INVx1_ASAP7_75t_SL fopt13870 (.A(n_3650),
    .Y(n_3649));
 HB1xp67_ASAP7_75t_SL fopt13871 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .Y(n_3650));
 HB1xp67_ASAP7_75t_SL fopt13872 (.A(n_12033),
    .Y(n_3652));
 INVx1_ASAP7_75t_SL fopt13873 (.A(n_3655),
    .Y(n_3654));
 HB1xp67_ASAP7_75t_SL fopt13874 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .Y(n_3655));
 HB1xp67_ASAP7_75t_SL fopt13876 (.A(n_23426),
    .Y(n_3659));
 HB1xp67_ASAP7_75t_SL fopt13877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_44),
    .Y(n_3661));
 INVx1_ASAP7_75t_SL fopt13881 (.A(n_3669),
    .Y(n_3668));
 HB1xp67_ASAP7_75t_SL fopt13882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .Y(n_3669));
 INVxp67_ASAP7_75t_SL fopt13888 (.A(n_3681),
    .Y(n_3679));
 INVxp67_ASAP7_75t_SL fopt13892 (.A(n_3687),
    .Y(n_3685));
 INVxp67_ASAP7_75t_SL fopt13893 (.A(n_3687),
    .Y(n_3686));
 HB1xp67_ASAP7_75t_SL fopt13894 (.A(n_9627),
    .Y(n_3687));
 BUFx3_ASAP7_75t_SL fopt13905 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(n_3706));
 INVxp67_ASAP7_75t_SL fopt13907 (.A(n_3711),
    .Y(n_3709));
 INVxp67_ASAP7_75t_SL fopt13908 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(n_3711));
 INVxp67_ASAP7_75t_SL fopt13909 (.A(n_3713),
    .Y(n_3714));
 BUFx6f_ASAP7_75t_SL fopt13912 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(n_3713));
 INVxp67_ASAP7_75t_SL fopt13920 (.A(n_3738),
    .Y(n_3736));
 INVxp67_ASAP7_75t_SL fopt13921 (.A(n_3738),
    .Y(n_3737));
 HB1xp67_ASAP7_75t_SL fopt13922 (.A(n_9513),
    .Y(n_3738));
 INVxp67_ASAP7_75t_SL fopt13926 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_205),
    .Y(n_3746));
 INVx1_ASAP7_75t_SL fopt13929 (.A(n_3759),
    .Y(n_3761));
 INVxp67_ASAP7_75t_SL fopt13930 (.A(n_3760),
    .Y(n_3759));
 BUFx3_ASAP7_75t_SL fopt13931 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(n_3760));
 HB1xp67_ASAP7_75t_SL fopt13932 (.A(n_10236),
    .Y(n_3766));
 INVxp67_ASAP7_75t_SL fopt13934 (.A(n_9271),
    .Y(n_3770));
 HB1xp67_ASAP7_75t_SL fopt13940 (.A(n_17491),
    .Y(n_3782));
 INVx1_ASAP7_75t_SL fopt13947 (.A(n_3796),
    .Y(n_3795));
 HB1xp67_ASAP7_75t_SL fopt13948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_23),
    .Y(n_3796));
 HB1xp67_ASAP7_75t_SL fopt13959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_32),
    .Y(n_3815));
 HB1xp67_ASAP7_75t_SL fopt13960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_32),
    .Y(n_3817));
 HB1xp67_ASAP7_75t_SL fopt13961 (.A(n_17830),
    .Y(n_3819));
 HB1xp67_ASAP7_75t_SL fopt13963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_32),
    .Y(n_3823));
 HB1xp67_ASAP7_75t_SL fopt13965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_107),
    .Y(n_3827));
 HB1xp67_ASAP7_75t_SL fopt13968 (.A(n_10294),
    .Y(n_3833));
 HB1xp67_ASAP7_75t_SL fopt13978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_32),
    .Y(n_3860));
 BUFx12f_ASAP7_75t_SL fopt13982 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(n_3868));
 HB1xp67_ASAP7_75t_SL fopt13983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_29),
    .Y(n_3877));
 INVx1_ASAP7_75t_SL fopt13984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_29),
    .Y(n_3878));
 HB1xp67_ASAP7_75t_SL fopt13985 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_32),
    .Y(n_3880));
 INVxp67_ASAP7_75t_SL fopt13986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_131),
    .Y(n_3882));
 HB1xp67_ASAP7_75t_SL fopt13993 (.A(n_22567),
    .Y(n_3893));
 HB1xp67_ASAP7_75t_SL fopt13998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_32),
    .Y(n_3901));
 BUFx3_ASAP7_75t_SL fopt14 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(n_3112));
 INVx1_ASAP7_75t_SL fopt140 (.A(n_10640),
    .Y(n_10641));
 HB1xp67_ASAP7_75t_SL fopt14000 (.A(n_8841),
    .Y(n_3905));
 HB1xp67_ASAP7_75t_SL fopt14001 (.A(n_23113),
    .Y(n_3907));
 HB1xp67_ASAP7_75t_SL fopt14005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_25),
    .Y(n_3915));
 HB1xp67_ASAP7_75t_SL fopt14006 (.A(n_3918),
    .Y(n_3917));
 INVx1_ASAP7_75t_SL fopt14007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_222),
    .Y(n_3918));
 HB1xp67_ASAP7_75t_SL fopt14009 (.A(n_3923),
    .Y(n_3922));
 INVx1_ASAP7_75t_SL fopt14010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_222),
    .Y(n_3923));
 HB1xp67_ASAP7_75t_SL fopt14018 (.A(n_12780),
    .Y(n_3938));
 HB1xp67_ASAP7_75t_SL fopt14020 (.A(n_21479),
    .Y(n_3942));
 HB1xp67_ASAP7_75t_SL fopt14021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_153),
    .Y(n_3944));
 HB1xp67_ASAP7_75t_SL fopt14022 (.A(n_10327),
    .Y(n_3946));
 INVxp67_ASAP7_75t_SL fopt14024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_69),
    .Y(n_3950));
 HB1xp67_ASAP7_75t_SL fopt14026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_36),
    .Y(n_3953));
 HB1xp67_ASAP7_75t_SL fopt14027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_130),
    .Y(n_3955));
 INVxp67_ASAP7_75t_SL fopt14028 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .Y(n_3957));
 HB1xp67_ASAP7_75t_SL fopt14032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_36),
    .Y(n_3963));
 INVxp67_ASAP7_75t_SL fopt14033 (.A(n_18692),
    .Y(n_3965));
 HB1xp67_ASAP7_75t_SL fopt14037 (.A(n_7462),
    .Y(n_3971));
 HB1xp67_ASAP7_75t_SL fopt14038 (.A(n_25313),
    .Y(n_3973));
 INVxp67_ASAP7_75t_SL fopt14039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .Y(n_3975));
 HB1xp67_ASAP7_75t_SL fopt14044 (.A(n_10014),
    .Y(n_3983));
 HB1xp67_ASAP7_75t_SL fopt14046 (.A(n_10291),
    .Y(n_3987));
 INVx1_ASAP7_75t_SL fopt14047 (.A(n_10291),
    .Y(n_3988));
 HB1xp67_ASAP7_75t_SL fopt14048 (.A(n_6377),
    .Y(n_3990));
 HB1xp67_ASAP7_75t_SL fopt14052 (.A(n_14394),
    .Y(n_4012));
 INVx1_ASAP7_75t_SL fopt14056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_134),
    .Y(n_4017));
 HB1xp67_ASAP7_75t_SL fopt14058 (.A(n_22011),
    .Y(n_4022));
 HB1xp67_ASAP7_75t_SL fopt14059 (.A(n_22786),
    .Y(n_4024));
 INVxp67_ASAP7_75t_SL fopt14060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_69),
    .Y(n_4026));
 HB1xp67_ASAP7_75t_SL fopt14062 (.A(n_19282),
    .Y(n_4029));
 INVx1_ASAP7_75t_SL fopt14064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_69),
    .Y(n_4031));
 INVx1_ASAP7_75t_SL fopt14068 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_69),
    .Y(n_4038));
 HB1xp67_ASAP7_75t_SL fopt14069 (.A(n_21976),
    .Y(n_4041));
 INVxp67_ASAP7_75t_SL fopt14073 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .Y(n_4048));
 INVxp67_ASAP7_75t_SL fopt14081 (.A(n_4062),
    .Y(n_4061));
 INVxp67_ASAP7_75t_SL fopt14082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_285),
    .Y(n_4062));
 HB1xp67_ASAP7_75t_SL fopt14085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_42),
    .Y(n_4068));
 HB1xp67_ASAP7_75t_SL fopt14086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_42),
    .Y(n_4070));
 INVx1_ASAP7_75t_SL fopt14088 (.A(n_4075),
    .Y(n_4074));
 HB1xp67_ASAP7_75t_SL fopt14089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_23),
    .Y(n_4075));
 INVx1_ASAP7_75t_SL fopt14093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_446),
    .Y(n_4082));
 INVx1_ASAP7_75t_SL fopt14094 (.A(n_4085),
    .Y(n_4084));
 HB1xp67_ASAP7_75t_SL fopt14095 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_23),
    .Y(n_4085));
 INVx1_ASAP7_75t_SL fopt14096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_446),
    .Y(n_4087));
 HB1xp67_ASAP7_75t_SL fopt14097 (.A(n_12634),
    .Y(n_4089));
 HB1xp67_ASAP7_75t_SL fopt14101 (.A(n_20101),
    .Y(n_4095));
 HB1xp67_ASAP7_75t_SL fopt14105 (.A(n_4102),
    .Y(n_4101));
 INVx2_ASAP7_75t_SL fopt14106 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_329),
    .Y(n_4102));
 INVxp67_ASAP7_75t_SL fopt14109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_215),
    .Y(n_4107));
 INVx1_ASAP7_75t_SL fopt1411 (.A(n_18752),
    .Y(n_9202));
 INVx1_ASAP7_75t_SL fopt14121 (.A(n_4123),
    .Y(n_4124));
 BUFx3_ASAP7_75t_SL fopt14126 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(n_4123));
 INVxp67_ASAP7_75t_SL fopt14127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_205),
    .Y(n_4138));
 INVxp67_ASAP7_75t_SL fopt14128 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .Y(n_4140));
 INVx1_ASAP7_75t_SL fopt14148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_275),
    .Y(n_4193));
 INVx1_ASAP7_75t_SL fopt14150 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_275),
    .Y(n_4197));
 INVx1_ASAP7_75t_SL fopt14151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_275),
    .Y(n_4199));
 INVx1_ASAP7_75t_SL fopt14163 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_190),
    .Y(n_4224));
 INVxp67_ASAP7_75t_SL fopt14166 (.A(n_4231),
    .Y(n_4230));
 INVxp67_ASAP7_75t_SL fopt14168 (.A(n_4234),
    .Y(n_4233));
 INVxp67_ASAP7_75t_SL fopt14169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_285),
    .Y(n_4234));
 INVxp67_ASAP7_75t_SL fopt14172 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .Y(n_4239));
 HB1xp67_ASAP7_75t_SL fopt14176 (.A(n_4246),
    .Y(n_4245));
 INVx2_ASAP7_75t_SL fopt14177 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .Y(n_4246));
 HB1xp67_ASAP7_75t_SL fopt14178 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_22),
    .Y(n_4248));
 INVxp67_ASAP7_75t_SL fopt14179 (.A(n_4251),
    .Y(n_4250));
 INVxp67_ASAP7_75t_SL fopt14180 (.A(n_15813),
    .Y(n_4251));
 INVxp67_ASAP7_75t_SL fopt14181 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .Y(n_4253));
 INVxp67_ASAP7_75t_SL fopt14187 (.A(n_4263),
    .Y(n_4262));
 HB1xp67_ASAP7_75t_SL fopt14189 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .Y(n_4263));
 INVxp67_ASAP7_75t_SL fopt14191 (.A(n_6576),
    .Y(n_4268));
 BUFx6f_ASAP7_75t_SL fopt14195 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[12]),
    .Y(n_4275));
 INVxp67_ASAP7_75t_SL fopt14197 (.A(n_4286),
    .Y(n_4287));
 INVxp67_ASAP7_75t_SL fopt14207 (.A(n_4314),
    .Y(n_4315));
 BUFx6f_ASAP7_75t_SL fopt14208 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(n_4314));
 HB1xp67_ASAP7_75t_SL fopt14212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_153),
    .Y(n_4331));
 HB1xp67_ASAP7_75t_SL fopt14217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_22),
    .Y(n_4341));
 INVxp67_ASAP7_75t_SL fopt14226 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .Y(n_4354));
 HB1xp67_ASAP7_75t_SL fopt14233 (.A(n_8197),
    .Y(n_4365));
 INVxp67_ASAP7_75t_SL fopt14234 (.A(n_11833),
    .Y(n_4367));
 INVxp67_ASAP7_75t_SL fopt14241 (.A(n_14732),
    .Y(n_4377));
 INVxp67_ASAP7_75t_SL fopt14246 (.A(n_4386),
    .Y(n_4385));
 BUFx3_ASAP7_75t_SL fopt14247 (.A(n_22156),
    .Y(n_4386));
 HB1xp67_ASAP7_75t_SL fopt14250 (.A(n_8376),
    .Y(n_4403));
 INVx1_ASAP7_75t_SL fopt14251 (.A(n_8376),
    .Y(n_4404));
 HB1xp67_ASAP7_75t_SL fopt14253 (.A(n_10902),
    .Y(n_4408));
 HB1xp67_ASAP7_75t_SL fopt14254 (.A(n_13011),
    .Y(n_4410));
 INVx2_ASAP7_75t_SL fopt14297 (.A(n_6097),
    .Y(n_4451));
 INVxp67_ASAP7_75t_SL fopt14301 (.A(n_4462),
    .Y(n_4463));
 INVxp67_ASAP7_75t_SL fopt14302 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(n_4462));
 INVx1_ASAP7_75t_SL fopt14306 (.A(n_8134),
    .Y(n_4474));
 HB1xp67_ASAP7_75t_SL fopt14309 (.A(n_24405),
    .Y(n_4480));
 INVx1_ASAP7_75t_SL fopt14331 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_161),
    .Y(n_4518));
 INVxp67_ASAP7_75t_SL fopt14335 (.A(n_4521),
    .Y(n_4528));
 BUFx6f_ASAP7_75t_SL fopt14337 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(n_4521));
 HB1xp67_ASAP7_75t_SL fopt14338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_56),
    .Y(n_4539));
 HB1xp67_ASAP7_75t_SL fopt14339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_19),
    .Y(n_4541));
 INVx2_ASAP7_75t_SL fopt14341 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(n_4549));
 INVx3_ASAP7_75t_SL fopt14342 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(n_4550));
 INVx3_ASAP7_75t_SL fopt14348 (.A(n_4553),
    .Y(n_4555));
 BUFx3_ASAP7_75t_SL fopt14350 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(n_4553));
 HB1xp67_ASAP7_75t_SL fopt14351 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_239),
    .Y(n_4565));
 INVxp67_ASAP7_75t_SL fopt14443 (.A(n_12624),
    .Y(n_4665));
 INVx1_ASAP7_75t_SL fopt14448 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_33),
    .Y(n_4671));
 INVx2_ASAP7_75t_SL fopt14544 (.A(n_4768),
    .Y(n_4769));
 HB1xp67_ASAP7_75t_SL fopt14574 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_194),
    .Y(n_4805));
 INVxp67_ASAP7_75t_SL fopt14577 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_215),
    .Y(n_4810));
 INVx4_ASAP7_75t_SL fopt14586 (.A(n_4833),
    .Y(n_4826));
 INVx2_ASAP7_75t_SL fopt14587 (.A(n_4833),
    .Y(n_4831));
 INVx3_ASAP7_75t_SL fopt14589 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[36]),
    .Y(n_4833));
 HB1xp67_ASAP7_75t_SL fopt14594 (.A(n_10628),
    .Y(n_4842));
 INVx1_ASAP7_75t_SL fopt14595 (.A(n_10628),
    .Y(n_4843));
 INVx1_ASAP7_75t_SL fopt146 (.A(n_19354),
    .Y(n_19355));
 INVx2_ASAP7_75t_SL fopt14609 (.A(n_20976),
    .Y(n_4864));
 INVx1_ASAP7_75t_L fopt14615 (.A(n_4864),
    .Y(n_4865));
 INVxp67_ASAP7_75t_SL fopt14656 (.A(n_13477),
    .Y(n_4903));
 HB1xp67_ASAP7_75t_SL fopt14705 (.A(n_8091),
    .Y(n_4956));
 HB1xp67_ASAP7_75t_SL fopt14792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_32),
    .Y(n_5045));
 INVxp67_ASAP7_75t_SL fopt14793 (.A(n_5048),
    .Y(n_5047));
 HB1xp67_ASAP7_75t_SL fopt14794 (.A(n_6190),
    .Y(n_5048));
 INVxp67_ASAP7_75t_SL fopt14804 (.A(n_7960),
    .Y(n_5065));
 HB1xp67_ASAP7_75t_SL fopt14869 (.A(n_23683),
    .Y(n_5131));
 HB1xp67_ASAP7_75t_SL fopt14870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_22),
    .Y(n_5133));
 INVx1_ASAP7_75t_L fopt14872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_97),
    .Y(n_5137));
 HB1xp67_ASAP7_75t_SL fopt14990 (.A(n_12720),
    .Y(n_5301));
 HB1xp67_ASAP7_75t_SL fopt15036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_147),
    .Y(n_5385));
 HB1xp67_ASAP7_75t_SL fopt15051 (.A(n_5412),
    .Y(n_5413));
 INVxp67_ASAP7_75t_SL fopt15052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_151),
    .Y(n_5410));
 HB1xp67_ASAP7_75t_SL fopt15060 (.A(n_16058),
    .Y(n_5433));
 INVxp67_ASAP7_75t_SL fopt15072 (.A(n_23580),
    .Y(n_5450));
 HB1xp67_ASAP7_75t_SL fopt15083 (.A(n_20346),
    .Y(n_5473));
 HB1xp67_ASAP7_75t_SL fopt15154 (.A(n_9957),
    .Y(n_5589));
 HB1xp67_ASAP7_75t_SL fopt15158 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_27),
    .Y(n_5593));
 HB1xp67_ASAP7_75t_SL fopt15206 (.A(n_19900),
    .Y(n_5660));
 BUFx3_ASAP7_75t_SL fopt15257 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(n_5737));
 INVxp67_ASAP7_75t_SL fopt15324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_53),
    .Y(n_5811));
 HB1xp67_ASAP7_75t_SL fopt15378 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_24),
    .Y(n_5903));
 INVx2_ASAP7_75t_SL fopt15380 (.A(n_19827),
    .Y(n_5909));
 INVxp67_ASAP7_75t_SL fopt15426 (.A(n_5981),
    .Y(n_5982));
 INVx1_ASAP7_75t_SL fopt15460 (.A(n_18856),
    .Y(n_6076));
 HB1xp67_ASAP7_75t_SL fopt15462 (.A(n_18856),
    .Y(n_6078));
 HB1xp67_ASAP7_75t_SL fopt15596 (.A(n_19554),
    .Y(n_6326));
 BUFx3_ASAP7_75t_SL fopt15750 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[12]),
    .Y(n_6576));
 HB1xp67_ASAP7_75t_SL fopt15885 (.A(n_6730),
    .Y(n_6731));
 INVx1_ASAP7_75t_SL fopt15973 (.A(n_13295),
    .Y(n_6825));
 INVxp67_ASAP7_75t_SL fopt160 (.A(n_19787),
    .Y(n_8473));
 INVx3_ASAP7_75t_SL fopt16005 (.A(n_22742),
    .Y(n_6861));
 HB1xp67_ASAP7_75t_SL fopt16088 (.A(n_10481),
    .Y(n_6960));
 HB1xp67_ASAP7_75t_SL fopt16467 (.A(n_22055),
    .Y(n_7409));
 HB1xp67_ASAP7_75t_SL fopt16493 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_262),
    .Y(n_7435));
 HB1xp67_ASAP7_75t_SL fopt16606 (.A(n_7570),
    .Y(n_7571));
 HB1xp67_ASAP7_75t_SL fopt16628 (.A(n_7588),
    .Y(n_7589));
 HB1xp67_ASAP7_75t_SL fopt16652 (.A(n_18891),
    .Y(n_7612));
 HB1xp67_ASAP7_75t_SL fopt16904 (.A(n_20098),
    .Y(n_7883));
 HB1xp67_ASAP7_75t_SL fopt16927 (.A(n_9904),
    .Y(n_7907));
 HB1xp67_ASAP7_75t_SL fopt16978 (.A(n_14024),
    .Y(n_7960));
 HB1xp67_ASAP7_75t_SL fopt17 (.A(n_19395),
    .Y(n_19396));
 HB1xp67_ASAP7_75t_SL fopt17083 (.A(n_8067),
    .Y(n_8071));
 HB1xp67_ASAP7_75t_SL fopt17084 (.A(n_8068),
    .Y(n_8072));
 INVxp67_ASAP7_75t_SL fopt17189 (.A(n_19597),
    .Y(n_8191));
 INVx1_ASAP7_75t_SL fopt172 (.A(n_19898),
    .Y(n_19899));
 INVxp67_ASAP7_75t_SL fopt17273 (.A(n_19551),
    .Y(n_8283));
 HB1xp67_ASAP7_75t_SL fopt17307 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_26),
    .Y(n_8320));
 INVxp67_ASAP7_75t_SL fopt17313 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_26),
    .Y(n_8326));
 HB1xp67_ASAP7_75t_SL fopt17333 (.A(n_16325),
    .Y(n_8351));
 INVxp67_ASAP7_75t_SL fopt17418 (.A(n_23430),
    .Y(n_8441));
 INVx1_ASAP7_75t_SL fopt17481 (.A(n_8505),
    .Y(n_8507));
 INVxp33_ASAP7_75t_SL fopt17551 (.A(n_8585),
    .Y(n_2791));
 INVxp33_ASAP7_75t_SL fopt17581 (.A(n_22819),
    .Y(n_8637));
 HB1xp67_ASAP7_75t_SL fopt17606 (.A(n_8666),
    .Y(n_8667));
 INVxp33_ASAP7_75t_SL fopt17611 (.A(n_8672),
    .Y(n_5399));
 INVxp67_ASAP7_75t_SL fopt17622 (.A(n_8690),
    .Y(n_8691));
 HB1xp67_ASAP7_75t_SL fopt17675 (.A(n_18915),
    .Y(n_8747));
 HB1xp67_ASAP7_75t_SL fopt17676 (.A(n_8760),
    .Y(n_8761));
 HB1xp67_ASAP7_75t_SL fopt17697 (.A(n_8771),
    .Y(n_8772));
 INVx1_ASAP7_75t_SL fopt17698 (.A(n_18842),
    .Y(n_8771));
 HB1xp67_ASAP7_75t_SL fopt17699 (.A(n_18842),
    .Y(n_8773));
 HB1xp67_ASAP7_75t_SL fopt177 (.A(n_15590),
    .Y(n_19623));
 BUFx6f_ASAP7_75t_SL fopt17708 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[3]),
    .Y(n_6972));
 HB1xp67_ASAP7_75t_SL fopt17709 (.A(n_12287),
    .Y(n_8784));
 INVx1_ASAP7_75t_SL fopt17712 (.A(n_8799),
    .Y(n_8800));
 HB1xp67_ASAP7_75t_SL fopt17749 (.A(n_23036),
    .Y(n_8846));
 INVx2_ASAP7_75t_SL fopt178 (.A(n_20898),
    .Y(n_20899));
 HB1xp67_ASAP7_75t_SL fopt17864 (.A(n_8991),
    .Y(n_8992));
 INVxp67_ASAP7_75t_SL fopt17932 (.A(n_18751),
    .Y(n_9058));
 INVx1_ASAP7_75t_SL fopt18 (.A(n_19394),
    .Y(n_19395));
 HB1xp67_ASAP7_75t_SL fopt18078 (.A(n_22260),
    .Y(n_9231));
 INVx1_ASAP7_75t_SL fopt18082 (.A(n_12565),
    .Y(n_9235));
 INVxp33_ASAP7_75t_SL fopt181 (.A(n_14877),
    .Y(n_7926));
 HB1xp67_ASAP7_75t_SL fopt18100 (.A(n_9255),
    .Y(n_9256));
 INVx2_ASAP7_75t_SL fopt18115 (.A(n_9267),
    .Y(n_9269));
 HB1xp67_ASAP7_75t_SL fopt18164 (.A(n_9317),
    .Y(n_9322));
 BUFx6f_ASAP7_75t_SL fopt18191 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[12]),
    .Y(n_9349));
 INVxp33_ASAP7_75t_SL fopt18212 (.A(n_9368),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_76));
 INVxp67_ASAP7_75t_SL fopt18225 (.A(n_12374),
    .Y(n_9384));
 HB1xp67_ASAP7_75t_SL fopt18284 (.A(n_9450),
    .Y(n_9452));
 INVx1_ASAP7_75t_SL fopt18301 (.A(n_18754),
    .Y(n_9472));
 HB1xp67_ASAP7_75t_SL fopt18341 (.A(n_21961),
    .Y(n_9520));
 HB1xp67_ASAP7_75t_SL fopt18356 (.A(n_9534),
    .Y(n_9535));
 HB1xp67_ASAP7_75t_SL fopt18439 (.A(n_8613),
    .Y(n_9624));
 INVx1_ASAP7_75t_SL fopt18464 (.A(n_9650),
    .Y(n_9651));
 HB1xp67_ASAP7_75t_SL fopt18498 (.A(n_9686),
    .Y(n_9687));
 HB1xp67_ASAP7_75t_SL fopt18522 (.A(n_13148),
    .Y(n_9712));
 HB1xp67_ASAP7_75t_SL fopt18526 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_30),
    .Y(n_9714));
 HB1xp67_ASAP7_75t_SL fopt18544 (.A(n_12985),
    .Y(n_9735));
 INVx1_ASAP7_75t_SL fopt186 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_89),
    .Y(n_7315));
 INVxp33_ASAP7_75t_SL fopt18601 (.A(n_9792),
    .Y(n_9795));
 INVxp33_ASAP7_75t_SL fopt18631 (.A(n_19430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_76));
 HB1xp67_ASAP7_75t_SL fopt18682 (.A(n_13081),
    .Y(n_9879));
 HB1xp67_ASAP7_75t_SL fopt18688 (.A(n_9884),
    .Y(n_9885));
 INVxp33_ASAP7_75t_SL fopt18697 (.A(n_20164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_72));
 INVxp33_ASAP7_75t_R fopt187 (.A(n_12593),
    .Y(n_12595));
 INVxp67_ASAP7_75t_SL fopt18755 (.A(n_22429),
    .Y(n_9956));
 HB1xp67_ASAP7_75t_SL fopt18757 (.A(n_9959),
    .Y(n_9960));
 HB1xp67_ASAP7_75t_SL fopt18994 (.A(n_10200),
    .Y(n_10201));
 INVxp67_ASAP7_75t_SL fopt19 (.A(n_19393),
    .Y(n_19394));
 HB1xp67_ASAP7_75t_SL fopt19039 (.A(n_16327),
    .Y(n_10247));
 HB1xp67_ASAP7_75t_SL fopt19041 (.A(n_6968),
    .Y(n_10249));
 INVx1_ASAP7_75t_SL fopt19091 (.A(n_9389),
    .Y(n_10302));
 INVxp67_ASAP7_75t_SL fopt19168 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_127),
    .Y(n_10387));
 HB1xp67_ASAP7_75t_SL fopt19268 (.A(n_19827),
    .Y(n_10490));
 INVxp33_ASAP7_75t_SL fopt19269 (.A(n_11871),
    .Y(n_10492));
 INVx2_ASAP7_75t_SL fopt19345 (.A(n_7721),
    .Y(n_7724));
 INVx1_ASAP7_75t_L fopt19346 (.A(n_3461),
    .Y(n_10567));
 HB1xp67_ASAP7_75t_SL fopt19359 (.A(n_13929),
    .Y(n_10582));
 INVx1_ASAP7_75t_SL fopt19380 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_108),
    .Y(n_10601));
 HB1xp67_ASAP7_75t_SL fopt19392 (.A(n_26134),
    .Y(n_10617));
 INVxp67_ASAP7_75t_SL fopt19394 (.A(n_26000),
    .Y(n_10618));
 HB1xp67_ASAP7_75t_SL fopt19418 (.A(n_10641),
    .Y(n_10643));
 HB1xp67_ASAP7_75t_SL fopt19422 (.A(n_10645),
    .Y(n_10647));
 HB1xp67_ASAP7_75t_SL fopt19463 (.A(n_10693),
    .Y(n_10694));
 HB1xp67_ASAP7_75t_SL fopt19486 (.A(n_14698),
    .Y(n_10713));
 HB1xp67_ASAP7_75t_SL fopt19526 (.A(n_10757),
    .Y(n_10758));
 INVx1_ASAP7_75t_SL fopt19531 (.A(n_10757),
    .Y(n_10759));
 HB1xp67_ASAP7_75t_SL fopt19568 (.A(n_10796),
    .Y(n_10797));
 HB1xp67_ASAP7_75t_SL fopt19726 (.A(n_10964),
    .Y(n_10965));
 HB1xp67_ASAP7_75t_SL fopt19804 (.A(n_22968),
    .Y(n_11036));
 INVx1_ASAP7_75t_SL fopt19836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_28),
    .Y(n_11066));
 INVx3_ASAP7_75t_SL fopt2 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(n_12120));
 INVxp67_ASAP7_75t_SL fopt20010 (.A(n_11243),
    .Y(n_11248));
 HB1xp67_ASAP7_75t_SL fopt20023 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_251),
    .Y(n_11264));
 INVxp67_ASAP7_75t_SL fopt20191 (.A(n_18781),
    .Y(n_11444));
 HB1xp67_ASAP7_75t_SL fopt20277 (.A(n_20128),
    .Y(n_11610));
 BUFx6f_ASAP7_75t_SL fopt20409 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[60]),
    .Y(n_11770));
 INVx2_ASAP7_75t_SL fopt20421 (.A(n_11788),
    .Y(n_11789));
 HB1xp67_ASAP7_75t_SL fopt20466 (.A(n_11830),
    .Y(n_11833));
 INVx1_ASAP7_75t_SL fopt20512 (.A(n_10144),
    .Y(n_11887));
 INVx2_ASAP7_75t_SL fopt20536 (.A(n_11913),
    .Y(n_11914));
 HB1xp67_ASAP7_75t_SL fopt20605 (.A(n_20288),
    .Y(n_11984));
 INVx2_ASAP7_75t_SL fopt20682 (.A(n_23408),
    .Y(n_12114));
 INVx1_ASAP7_75t_SL fopt20688 (.A(n_12120),
    .Y(n_12124));
 INVx1_ASAP7_75t_SL fopt20691 (.A(n_12129),
    .Y(n_12134));
 BUFx6f_ASAP7_75t_SL fopt20692 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(n_12129));
 HB1xp67_ASAP7_75t_SL fopt20698 (.A(n_20759),
    .Y(n_12152));
 INVxp67_ASAP7_75t_SL fopt20699 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_102),
    .Y(n_12154));
 INVxp67_ASAP7_75t_SL fopt20896 (.A(n_10427),
    .Y(n_12392));
 INVxp67_ASAP7_75t_SL fopt20942 (.A(n_12498),
    .Y(n_12499));
 HB1xp67_ASAP7_75t_SL fopt21 (.A(n_19391),
    .Y(n_19393));
 INVx1_ASAP7_75t_SL fopt21037 (.A(n_12603),
    .Y(n_12604));
 HB1xp67_ASAP7_75t_SL fopt21344 (.A(n_13012),
    .Y(n_13013));
 INVxp67_ASAP7_75t_SL fopt21486 (.A(n_13173),
    .Y(n_13172));
 HB1xp67_ASAP7_75t_SL fopt21487 (.A(n_22487),
    .Y(n_13173));
 HB1xp67_ASAP7_75t_SL fopt21488 (.A(n_13176),
    .Y(n_13175));
 INVx1_ASAP7_75t_SL fopt21489 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_290),
    .Y(n_13176));
 INVx1_ASAP7_75t_SL fopt21490 (.A(n_10913),
    .Y(n_13178));
 INVxp67_ASAP7_75t_SRAM fopt21492 (.A(n_20936),
    .Y(n_13181));
 HB1xp67_ASAP7_75t_SL fopt21494 (.A(n_13186),
    .Y(n_13185));
 INVx1_ASAP7_75t_SL fopt21495 (.A(n_19882),
    .Y(n_13186));
 INVxp67_ASAP7_75t_SL fopt21496 (.A(n_23387),
    .Y(n_13188));
 HB1xp67_ASAP7_75t_SL fopt21497 (.A(n_13191),
    .Y(n_13190));
 INVx1_ASAP7_75t_SL fopt21498 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_159),
    .Y(n_13191));
 INVxp67_ASAP7_75t_SL fopt21499 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_151),
    .Y(n_13193));
 INVx1_ASAP7_75t_SL fopt21503 (.A(n_15939),
    .Y(n_13201));
 INVx1_ASAP7_75t_SL fopt21505 (.A(n_9350),
    .Y(n_13203));
 HB1xp67_ASAP7_75t_SL fopt21506 (.A(n_9350),
    .Y(n_13204));
 BUFx6f_ASAP7_75t_SL fopt21529 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[57]),
    .Y(n_13228));
 INVxp67_ASAP7_75t_SL fopt21530 (.A(n_2657),
    .Y(n_13230));
 BUFx3_ASAP7_75t_SL fopt21531 (.A(n_13228),
    .Y(n_2657));
 BUFx8_ASAP7_75t_SL fopt21533 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[57]),
    .Y(n_13231));
 HB1xp67_ASAP7_75t_SL fopt21660 (.A(n_13362),
    .Y(n_13364));
 HB1xp67_ASAP7_75t_SL fopt21700 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_273),
    .Y(n_13406));
 INVxp67_ASAP7_75t_SL fopt21714 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[52]),
    .Y(n_13423));
 INVx1_ASAP7_75t_SL fopt21732 (.A(n_9763),
    .Y(n_13440));
 INVxp67_ASAP7_75t_SL fopt21737 (.A(n_14368),
    .Y(n_13449));
 HB1xp67_ASAP7_75t_SL fopt21785 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_75),
    .Y(n_13504));
 HB1xp67_ASAP7_75t_SL fopt21800 (.A(n_13522),
    .Y(n_13523));
 HB1xp67_ASAP7_75t_SL fopt21816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_675),
    .Y(n_13539));
 INVx2_ASAP7_75t_SL fopt21873 (.A(n_13599),
    .Y(n_13600));
 INVx1_ASAP7_75t_SL fopt21930 (.A(n_6673),
    .Y(n_13667));
 HB1xp67_ASAP7_75t_SL fopt21932 (.A(n_21372),
    .Y(n_13674));
 INVxp67_ASAP7_75t_SL fopt21933 (.A(n_8847),
    .Y(n_13676));
 INVxp67_ASAP7_75t_SL fopt21934 (.A(n_18009),
    .Y(n_13678));
 INVx1_ASAP7_75t_SL fopt21936 (.A(n_14675),
    .Y(n_13681));
 HB1xp67_ASAP7_75t_SL fopt21938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_36),
    .Y(n_13685));
 HB1xp67_ASAP7_75t_SL fopt21939 (.A(n_17655),
    .Y(n_13687));
 INVx1_ASAP7_75t_SL fopt21940 (.A(n_17655),
    .Y(n_13688));
 HB1xp67_ASAP7_75t_SL fopt21944 (.A(n_21830),
    .Y(n_13694));
 INVx2_ASAP7_75t_SL fopt21946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_95),
    .Y(n_13697));
 INVx2_ASAP7_75t_SL fopt21947 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_53),
    .Y(n_13699));
 HB1xp67_ASAP7_75t_SL fopt21948 (.A(n_10235),
    .Y(n_13701));
 INVx1_ASAP7_75t_SL fopt21949 (.A(n_10235),
    .Y(n_13702));
 BUFx12f_ASAP7_75t_SL fopt21952 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .Y(n_13707));
 INVx1_ASAP7_75t_SL fopt22122 (.A(n_13880),
    .Y(n_13877));
 INVx2_ASAP7_75t_SL fopt22260 (.A(n_3112),
    .Y(n_3113));
 INVx1_ASAP7_75t_SL fopt22393 (.A(n_21931),
    .Y(n_14172));
 HB1xp67_ASAP7_75t_SL fopt22394 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_185),
    .Y(n_14174));
 INVxp67_ASAP7_75t_SL fopt22395 (.A(n_14177),
    .Y(n_14176));
 INVx1_ASAP7_75t_SL fopt22396 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_272),
    .Y(n_14177));
 INVx2_ASAP7_75t_SL fopt22398 (.A(n_14181),
    .Y(n_14179));
 INVx1_ASAP7_75t_SL fopt22402 (.A(n_14181),
    .Y(n_14186));
 INVx4_ASAP7_75t_SL fopt22405 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(n_14181));
 INVx3_ASAP7_75t_SL fopt22407 (.A(n_14181),
    .Y(n_14183));
 HB1xp67_ASAP7_75t_SL fopt22409 (.A(n_13056),
    .Y(n_14203));
 INVx1_ASAP7_75t_SL fopt22410 (.A(n_13056),
    .Y(n_14204));
 INVx1_ASAP7_75t_SL fopt22413 (.A(n_23685),
    .Y(n_14208));
 INVxp67_ASAP7_75t_SL fopt22414 (.A(n_14213),
    .Y(n_14211));
 INVx2_ASAP7_75t_SL fopt22416 (.A(n_7255),
    .Y(n_14213));
 INVx1_ASAP7_75t_SL fopt22571 (.A(n_14373),
    .Y(n_2718));
 INVx2_ASAP7_75t_SL fopt22572 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_14372));
 HB1xp67_ASAP7_75t_SL fopt22583 (.A(n_22626),
    .Y(n_14388));
 INVxp67_ASAP7_75t_SL fopt22624 (.A(n_14425),
    .Y(n_14429));
 BUFx6f_ASAP7_75t_SL fopt22704 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_14523));
 HB1xp67_ASAP7_75t_SL fopt22708 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_14537));
 BUFx3_ASAP7_75t_SL fopt22821 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[43]),
    .Y(n_14674));
 INVx2_ASAP7_75t_SL fopt22938 (.A(n_14798),
    .Y(n_14800));
 INVxp67_ASAP7_75t_SL fopt22947 (.A(n_14810),
    .Y(n_14811));
 INVx1_ASAP7_75t_SL fopt23 (.A(n_16253),
    .Y(n_20156));
 INVxp67_ASAP7_75t_SL fopt23066 (.A(n_14938),
    .Y(n_14947));
 HB1xp67_ASAP7_75t_SL fopt23068 (.A(n_10648),
    .Y(n_14951));
 INVxp67_ASAP7_75t_SL fopt23083 (.A(n_14978),
    .Y(n_14977));
 BUFx3_ASAP7_75t_SL fopt23084 (.A(n_14975),
    .Y(n_14978));
 INVx2_ASAP7_75t_SL fopt23085 (.A(n_21989),
    .Y(n_14975));
 BUFx3_ASAP7_75t_SL fopt23087 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[28]),
    .Y(n_14981));
 INVx2_ASAP7_75t_SL fopt23088 (.A(n_14986),
    .Y(n_14984));
 INVx2_ASAP7_75t_SL fopt23089 (.A(n_14986),
    .Y(n_14985));
 INVx5_ASAP7_75t_SL fopt23093 (.A(n_14986),
    .Y(n_14987));
 INVxp67_ASAP7_75t_SL fopt23096 (.A(n_14457),
    .Y(n_14998));
 INVxp67_ASAP7_75t_SL fopt23097 (.A(n_15001),
    .Y(n_15000));
 INVx1_ASAP7_75t_SL fopt23098 (.A(n_21437),
    .Y(n_15001));
 INVxp67_ASAP7_75t_SL fopt23104 (.A(n_15014),
    .Y(n_15013));
 INVxp67_ASAP7_75t_SL fopt23122 (.A(n_15045),
    .Y(n_15046));
 BUFx6f_ASAP7_75t_SL fopt23127 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(n_15045));
 HB1xp67_ASAP7_75t_SL fopt23128 (.A(n_11515),
    .Y(n_15060));
 HB1xp67_ASAP7_75t_SL fopt23131 (.A(n_15068),
    .Y(n_15067));
 INVxp67_ASAP7_75t_SL fopt23132 (.A(n_17420),
    .Y(n_15068));
 INVxp67_ASAP7_75t_SL fopt23133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_145),
    .Y(n_15070));
 INVx1_ASAP7_75t_SL fopt23134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_145),
    .Y(n_15071));
 INVx1_ASAP7_75t_SL fopt23137 (.A(n_9327),
    .Y(n_15077));
 HB1xp67_ASAP7_75t_SL fopt23138 (.A(n_13082),
    .Y(n_15079));
 INVxp67_ASAP7_75t_SL fopt23139 (.A(n_14671),
    .Y(n_15081));
 HB1xp67_ASAP7_75t_SL fopt23208 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .Y(n_15149));
 HB1xp67_ASAP7_75t_SL fopt23209 (.A(n_8505),
    .Y(n_15150));
 HB1xp67_ASAP7_75t_SL fopt23210 (.A(n_13968),
    .Y(n_15151));
 BUFx6f_ASAP7_75t_SL fopt23220 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(n_15192));
 INVxp67_ASAP7_75t_SL fopt23223 (.A(n_15201),
    .Y(n_15200));
 BUFx3_ASAP7_75t_SL fopt23226 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(n_15201));
 INVx2_ASAP7_75t_SL fopt23227 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_145),
    .Y(n_15210));
 INVx2_ASAP7_75t_SL fopt23229 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_204),
    .Y(n_15213));
 INVx1_ASAP7_75t_SL fopt23230 (.A(n_15584),
    .Y(n_15215));
 HB1xp67_ASAP7_75t_SL fopt23231 (.A(n_15218),
    .Y(n_15217));
 INVx2_ASAP7_75t_SL fopt23232 (.A(n_19783),
    .Y(n_15218));
 INVx1_ASAP7_75t_SL fopt23236 (.A(n_11084),
    .Y(n_15223));
 HB1xp67_ASAP7_75t_SL fopt23237 (.A(n_15227),
    .Y(n_15226));
 INVx1_ASAP7_75t_SL fopt23238 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_316),
    .Y(n_15227));
 INVxp67_ASAP7_75t_SL fopt23240 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_155),
    .Y(n_15231));
 HB1xp67_ASAP7_75t_SL fopt23241 (.A(n_9671),
    .Y(n_15233));
 HB1xp67_ASAP7_75t_SL fopt23242 (.A(n_14025),
    .Y(n_15235));
 INVxp67_ASAP7_75t_SL fopt23244 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_91),
    .Y(n_15239));
 INVx1_ASAP7_75t_SL fopt23245 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_91),
    .Y(n_15240));
 HB1xp67_ASAP7_75t_SL fopt23326 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_104),
    .Y(n_15324));
 INVx1_ASAP7_75t_SL fopt23327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_104),
    .Y(n_15325));
 INVxp67_ASAP7_75t_SL fopt23331 (.A(n_18798),
    .Y(n_15332));
 INVxp67_ASAP7_75t_SL fopt23333 (.A(n_19432),
    .Y(n_15334));
 HB1xp67_ASAP7_75t_SL fopt23341 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_21),
    .Y(n_15355));
 INVx1_ASAP7_75t_SL fopt23343 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_253),
    .Y(n_15358));
 INVxp67_ASAP7_75t_SL fopt23345 (.A(n_11456),
    .Y(n_15361));
 HB1xp67_ASAP7_75t_SL fopt23356 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_263),
    .Y(n_15380));
 BUFx2_ASAP7_75t_SL fopt23358 (.A(n_22622),
    .Y(n_15384));
 INVxp67_ASAP7_75t_SL fopt23359 (.A(n_23416),
    .Y(n_15386));
 INVx1_ASAP7_75t_SL fopt23432 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_143),
    .Y(n_15462));
 INVxp67_ASAP7_75t_SL fopt23433 (.A(n_11085),
    .Y(n_15464));
 INVx1_ASAP7_75t_SL fopt23701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .Y(n_15740));
 INVxp67_ASAP7_75t_SL fopt24 (.A(n_22079),
    .Y(n_22080));
 INVxp33_ASAP7_75t_SRAM fopt241 (.A(n_8770),
    .Y(n_6255));
 INVxp67_ASAP7_75t_SL fopt24184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .Y(n_16247));
 INVxp67_ASAP7_75t_SL fopt24191 (.A(n_16253),
    .Y(n_16256));
 INVxp67_ASAP7_75t_SL fopt24283 (.A(n_16349),
    .Y(n_16352));
 INVxp67_ASAP7_75t_SL fopt24328 (.A(n_12494),
    .Y(n_16397));
 INVx1_ASAP7_75t_SL fopt244 (.A(n_11359),
    .Y(n_11356));
 INVxp67_ASAP7_75t_SL fopt24602 (.A(n_16684),
    .Y(n_16685));
 INVx1_ASAP7_75t_SL fopt24604 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .Y(n_16684));
 INVxp67_ASAP7_75t_SL fopt24660 (.A(n_16749),
    .Y(n_16751));
 BUFx6f_ASAP7_75t_SL fopt24661 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[20]),
    .Y(n_16749));
 BUFx6f_ASAP7_75t_SL fopt24662 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[20]),
    .Y(n_16753));
 BUFx6f_ASAP7_75t_SL fopt24664 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[20]),
    .Y(n_16757));
 INVxp67_ASAP7_75t_SL fopt24665 (.A(n_16763),
    .Y(n_16764));
 BUFx6f_ASAP7_75t_SL fopt24666 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[44]),
    .Y(n_16763));
 BUFx6f_ASAP7_75t_SL fopt24667 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[44]),
    .Y(n_16769));
 BUFx6f_ASAP7_75t_SL fopt24668 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[44]),
    .Y(n_16772));
 HB1xp67_ASAP7_75t_SL fopt24961 (.A(n_17075),
    .Y(n_17076));
 HB1xp67_ASAP7_75t_SL fopt251 (.A(n_20856),
    .Y(n_20767));
 INVxp67_ASAP7_75t_SL fopt25313 (.A(n_18828),
    .Y(n_17438));
 INVxp67_ASAP7_75t_SRAM fopt25453 (.A(n_11932),
    .Y(n_17587));
 INVxp67_ASAP7_75t_SL fopt25622 (.A(n_9892),
    .Y(n_17754));
 HB1xp67_ASAP7_75t_SL fopt25775 (.A(n_5456),
    .Y(n_17908));
 INVxp67_ASAP7_75t_SL fopt25882 (.A(n_18031),
    .Y(n_18034));
 BUFx6f_ASAP7_75t_SL fopt25884 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[35]),
    .Y(n_18031));
 HB1xp67_ASAP7_75t_SL fopt25885 (.A(n_18039),
    .Y(n_18041));
 BUFx6f_ASAP7_75t_SL fopt25886 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[35]),
    .Y(n_18039));
 INVxp67_ASAP7_75t_SL fopt25888 (.A(n_18049),
    .Y(n_18050));
 BUFx3_ASAP7_75t_SL fopt25891 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(n_18049));
 INVxp67_ASAP7_75t_SL fopt25911 (.A(n_18085),
    .Y(n_18084));
 INVxp67_ASAP7_75t_SL fopt25912 (.A(n_16158),
    .Y(n_18085));
 INVxp67_ASAP7_75t_SL fopt25979 (.A(n_18155),
    .Y(n_18154));
 HB1xp67_ASAP7_75t_SL fopt25980 (.A(n_9246),
    .Y(n_18155));
 INVx2_ASAP7_75t_SL fopt25982 (.A(n_9246),
    .Y(n_18157));
 INVxp67_ASAP7_75t_SL fopt26386 (.A(n_9432),
    .Y(n_18597));
 INVxp67_ASAP7_75t_SL fopt26393 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_421),
    .Y(n_18605));
 INVx2_ASAP7_75t_SL fopt26432 (.A(n_21146),
    .Y(n_18648));
 INVxp67_ASAP7_75t_SL fopt27032 (.A(n_24670),
    .Y(n_19263));
 HB1xp67_ASAP7_75t_SL fopt27041 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_250),
    .Y(n_19274));
 HB1xp67_ASAP7_75t_SL fopt27042 (.A(n_19278),
    .Y(n_19289));
 BUFx6f_ASAP7_75t_SL fopt27082 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(n_19340));
 BUFx3_ASAP7_75t_SL fopt27083 (.A(n_19340),
    .Y(n_19342));
 HB1xp67_ASAP7_75t_SL fopt27096 (.A(n_7682),
    .Y(n_19357));
 INVxp67_ASAP7_75t_SL fopt27124 (.A(n_19387),
    .Y(n_19390));
 BUFx12f_ASAP7_75t_SL fopt27126 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[47]),
    .Y(n_19391));
 INVx1_ASAP7_75t_L fopt27140 (.A(n_19410),
    .Y(n_19411));
 HB1xp67_ASAP7_75t_SL fopt27168 (.A(n_19441),
    .Y(n_19442));
 INVxp33_ASAP7_75t_SRAM fopt27200 (.A(n_26009),
    .Y(n_19484));
 INVxp67_ASAP7_75t_SL fopt27293 (.A(n_19598),
    .Y(n_19600));
 HB1xp67_ASAP7_75t_SL fopt273 (.A(n_13014),
    .Y(n_13015));
 INVxp67_ASAP7_75t_SRAM fopt27309 (.A(n_21159),
    .Y(n_19621));
 INVxp33_ASAP7_75t_SL fopt27312 (.A(n_19622),
    .Y(n_10032));
 INVxp67_ASAP7_75t_SL fopt27326 (.A(n_24679),
    .Y(n_19644));
 BUFx12f_ASAP7_75t_SL fopt27328 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[27]),
    .Y(n_19645));
 HB1xp67_ASAP7_75t_SL fopt27330 (.A(n_18939),
    .Y(n_19648));
 HB1xp67_ASAP7_75t_SL fopt27386 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_20),
    .Y(n_19714));
 HB1xp67_ASAP7_75t_SL fopt27438 (.A(n_10972),
    .Y(n_19777));
 INVxp67_ASAP7_75t_SL fopt27449 (.A(n_19792),
    .Y(n_19789));
 HB1xp67_ASAP7_75t_SL fopt27463 (.A(n_19802),
    .Y(n_19803));
 HB1xp67_ASAP7_75t_SL fopt27470 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_177),
    .Y(n_19810));
 HB1xp67_ASAP7_75t_SL fopt27531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_111),
    .Y(n_19877));
 INVx2_ASAP7_75t_SL fopt27539 (.A(n_10225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_193));
 HB1xp67_ASAP7_75t_SL fopt27653 (.A(n_19407),
    .Y(n_20006));
 INVx1_ASAP7_75t_SL fopt27657 (.A(n_19407),
    .Y(n_20008));
 INVx1_ASAP7_75t_SL fopt27661 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_171),
    .Y(n_20013));
 HB1xp67_ASAP7_75t_SL fopt27687 (.A(n_20044),
    .Y(n_20045));
 INVx1_ASAP7_75t_SL fopt27786 (.A(n_26120),
    .Y(n_20151));
 HB1xp67_ASAP7_75t_SL fopt27847 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_21),
    .Y(n_20223));
 HB1xp67_ASAP7_75t_SL fopt27855 (.A(n_20231),
    .Y(n_20232));
 BUFx3_ASAP7_75t_SL fopt28 (.A(n_2307),
    .Y(n_2293));
 HB1xp67_ASAP7_75t_SL fopt28007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_237),
    .Y(n_20401));
 INVxp67_ASAP7_75t_SL fopt28009 (.A(n_23166),
    .Y(n_20405));
 INVxp67_ASAP7_75t_SL fopt28014 (.A(n_26017),
    .Y(n_20413));
 HB1xp67_ASAP7_75t_SL fopt28020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_23),
    .Y(n_20421));
 INVx1_ASAP7_75t_SL fopt28021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_23),
    .Y(n_20422));
 INVxp67_ASAP7_75t_SL fopt28035 (.A(n_20464),
    .Y(n_20463));
 HB1xp67_ASAP7_75t_SL fopt28039 (.A(n_20459),
    .Y(n_20464));
 BUFx6f_ASAP7_75t_SL fopt28040 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(n_20459));
 HB1xp67_ASAP7_75t_SL fopt28041 (.A(n_20376),
    .Y(n_20478));
 HB1xp67_ASAP7_75t_SL fopt28042 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_17),
    .Y(n_20480));
 INVx1_ASAP7_75t_SL fopt28043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_17),
    .Y(n_20481));
 HB1xp67_ASAP7_75t_SL fopt28047 (.A(n_12213),
    .Y(n_20488));
 INVxp67_ASAP7_75t_SL fopt28050 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_106),
    .Y(n_20494));
 INVxp67_ASAP7_75t_SL fopt28051 (.A(n_20296),
    .Y(n_20496));
 INVxp67_ASAP7_75t_SL fopt28053 (.A(n_20501),
    .Y(n_20500));
 INVxp67_ASAP7_75t_SL fopt28054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_285),
    .Y(n_20501));
 INVxp67_ASAP7_75t_SL fopt28055 (.A(n_20504),
    .Y(n_20503));
 HB1xp67_ASAP7_75t_SL fopt28057 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .Y(n_20504));
 INVxp67_ASAP7_75t_SL fopt28060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_83),
    .Y(n_20510));
 INVx2_ASAP7_75t_SL fopt28061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_102),
    .Y(n_20512));
 INVx1_ASAP7_75t_L fopt28065 (.A(n_23138),
    .Y(n_20519));
 INVx2_ASAP7_75t_SL fopt28066 (.A(n_23138),
    .Y(n_20520));
 HB1xp67_ASAP7_75t_SL fopt28169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_18),
    .Y(n_20674));
 HB1xp67_ASAP7_75t_SL fopt28214 (.A(n_20717),
    .Y(n_20720));
 HB1xp67_ASAP7_75t_SL fopt28252 (.A(n_25311),
    .Y(n_20764));
 HB1xp67_ASAP7_75t_SL fopt283 (.A(n_21880),
    .Y(n_21881));
 INVxp67_ASAP7_75t_SL fopt28373 (.A(n_20899),
    .Y(n_20901));
 HB1xp67_ASAP7_75t_SL fopt28427 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_21),
    .Y(n_20967));
 INVxp67_ASAP7_75t_SL fopt28432 (.A(n_20972),
    .Y(n_20975));
 HB1xp67_ASAP7_75t_SL fopt28522 (.A(n_21083),
    .Y(n_21084));
 INVxp67_ASAP7_75t_SL fopt28529 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120),
    .Y(n_21075));
 INVx1_ASAP7_75t_L fopt28546 (.A(n_9342),
    .Y(n_21092));
 INVx4_ASAP7_75t_SL fopt28627 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[2]),
    .Y(n_21185));
 HB1xp67_ASAP7_75t_SL fopt28648 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_139),
    .Y(n_21206));
 INVxp67_ASAP7_75t_SL fopt28652 (.A(n_25921),
    .Y(n_21211));
 INVx1_ASAP7_75t_SL fopt28714 (.A(n_21276),
    .Y(n_21277));
 INVx1_ASAP7_75t_SL fopt28716 (.A(n_26135),
    .Y(n_21282));
 INVx1_ASAP7_75t_SL fopt28723 (.A(n_21285),
    .Y(n_21286));
 HB1xp67_ASAP7_75t_SL fopt28725 (.A(n_21286),
    .Y(n_21288));
 INVx1_ASAP7_75t_SL fopt28790 (.A(n_22456),
    .Y(n_21359));
 INVxp67_ASAP7_75t_SL fopt28793 (.A(n_22456),
    .Y(n_21361));
 HB1xp67_ASAP7_75t_SL fopt28794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_22),
    .Y(n_21362));
 INVxp67_ASAP7_75t_SRAM fopt28799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255),
    .Y(n_21367));
 HB1xp67_ASAP7_75t_SL fopt28820 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_234),
    .Y(n_21387));
 HB1xp67_ASAP7_75t_SL fopt28827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_22),
    .Y(n_21397));
 HB1xp67_ASAP7_75t_SL fopt28839 (.A(n_21410),
    .Y(n_21411));
 INVxp67_ASAP7_75t_SL fopt28856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_250),
    .Y(n_21427));
 HB1xp67_ASAP7_75t_SL fopt28858 (.A(n_21429),
    .Y(n_21430));
 HB1xp67_ASAP7_75t_SL fopt28865 (.A(n_26252),
    .Y(n_21435));
 HB1xp67_ASAP7_75t_SL fopt28920 (.A(n_21489),
    .Y(n_21492));
 HB1xp67_ASAP7_75t_SL fopt28948 (.A(n_9156),
    .Y(n_21520));
 INVx2_ASAP7_75t_SL fopt28972 (.A(n_21543),
    .Y(n_21544));
 HB1xp67_ASAP7_75t_SL fopt28974 (.A(n_21544),
    .Y(n_21546));
 HB1xp67_ASAP7_75t_SL fopt28981 (.A(n_21552),
    .Y(n_21553));
 HB1xp67_ASAP7_75t_SL fopt29004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_290),
    .Y(n_21576));
 HB1xp67_ASAP7_75t_SL fopt29042 (.A(n_21617),
    .Y(n_21618));
 HB1xp67_ASAP7_75t_SL fopt29050 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_251),
    .Y(n_21622));
 HB1xp67_ASAP7_75t_SL fopt29066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_683),
    .Y(n_21638));
 HB1xp67_ASAP7_75t_SL fopt29067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_587),
    .Y(n_21639));
 INVx1_ASAP7_75t_SL fopt29081 (.A(n_18843),
    .Y(n_21649));
 INVx1_ASAP7_75t_SL fopt29092 (.A(n_21675),
    .Y(n_21676));
 HB1xp67_ASAP7_75t_SL fopt29095 (.A(n_21676),
    .Y(n_21679));
 HB1xp67_ASAP7_75t_SL fopt29103 (.A(n_21686),
    .Y(n_21687));
 INVxp67_ASAP7_75t_SL fopt29253 (.A(n_23365),
    .Y(n_21848));
 HB1xp67_ASAP7_75t_SL fopt29319 (.A(n_21927),
    .Y(n_21928));
 HB1xp67_ASAP7_75t_SL fopt29344 (.A(n_26212),
    .Y(n_21951));
 INVx2_ASAP7_75t_SL fopt29381 (.A(n_21989),
    .Y(n_21990));
 INVx2_ASAP7_75t_SL fopt29382 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[28]),
    .Y(n_21989));
 HB1xp67_ASAP7_75t_SL fopt29385 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_24),
    .Y(n_21994));
 INVxp67_ASAP7_75t_SL fopt29391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_621),
    .Y(n_21999));
 BUFx12f_ASAP7_75t_SL fopt29410 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[63]),
    .Y(n_22019));
 HB1xp67_ASAP7_75t_SL fopt29413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_74),
    .Y(n_22023));
 HB1xp67_ASAP7_75t_SL fopt29455 (.A(n_22073),
    .Y(n_22074));
 INVxp67_ASAP7_75t_SL fopt29457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_101),
    .Y(n_22069));
 INVxp67_ASAP7_75t_SL fopt29466 (.A(n_22080),
    .Y(n_22082));
 HB1xp67_ASAP7_75t_SL fopt29491 (.A(n_22112),
    .Y(n_22113));
 INVx1_ASAP7_75t_SL fopt29525 (.A(n_23228),
    .Y(n_22141));
 HB1xp67_ASAP7_75t_SL fopt29539 (.A(n_22157),
    .Y(n_22158));
 INVxp33_ASAP7_75t_SL fopt29543 (.A(n_22156),
    .Y(n_22161));
 BUFx3_ASAP7_75t_SL fopt29597 (.A(n_17487),
    .Y(n_22214));
 INVx2_ASAP7_75t_SL fopt29607 (.A(n_22230),
    .Y(n_22231));
 INVxp33_ASAP7_75t_SL fopt29628 (.A(n_22244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_72));
 INVxp67_ASAP7_75t_SL fopt29634 (.A(n_26153),
    .Y(n_22256));
 INVx2_ASAP7_75t_SL fopt29779 (.A(n_15003),
    .Y(n_22416));
 HB1xp67_ASAP7_75t_SL fopt29781 (.A(n_22427),
    .Y(n_22428));
 INVxp67_ASAP7_75t_SL fopt29788 (.A(n_19007),
    .Y(n_22423));
 HB1xp67_ASAP7_75t_SL fopt29946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_22),
    .Y(n_22594));
 INVx1_ASAP7_75t_SL fopt29948 (.A(n_21593),
    .Y(n_22596));
 INVx1_ASAP7_75t_SL fopt29953 (.A(n_8105),
    .Y(n_22604));
 INVxp67_ASAP7_75t_SL fopt29954 (.A(n_22794),
    .Y(n_22606));
 INVx5_ASAP7_75t_SL fopt29962 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[43]),
    .Y(n_22615));
 INVx5_ASAP7_75t_SL fopt29964 (.A(n_22615),
    .Y(n_22616));
 INVxp67_ASAP7_75t_SL fopt29984 (.A(n_22637),
    .Y(n_22638));
 INVxp67_ASAP7_75t_SL fopt3 (.A(n_22019),
    .Y(n_19410));
 BUFx6f_ASAP7_75t_SL fopt30 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(n_2307));
 INVx3_ASAP7_75t_SL fopt30088 (.A(n_22742),
    .Y(n_22743));
 HB1xp67_ASAP7_75t_SL fopt30089 (.A(n_22744),
    .Y(n_22745));
 INVxp67_ASAP7_75t_SL fopt30144 (.A(n_22834),
    .Y(n_22836));
 BUFx3_ASAP7_75t_SL fopt30146 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_22834));
 INVxp67_ASAP7_75t_SL fopt30176 (.A(n_22865),
    .Y(n_22866));
 BUFx3_ASAP7_75t_SL fopt30177 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22865));
 BUFx6f_ASAP7_75t_SL fopt30196 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22886));
 INVxp67_ASAP7_75t_SL fopt30197 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22879));
 HB1xp67_ASAP7_75t_SL fopt30284 (.A(n_22973),
    .Y(n_22974));
 HB1xp67_ASAP7_75t_SL fopt30305 (.A(n_22994),
    .Y(n_22995));
 HB1xp67_ASAP7_75t_SL fopt30307 (.A(n_7893),
    .Y(n_22997));
 BUFx6f_ASAP7_75t_SL fopt30325 (.A(n_23016),
    .Y(n_15014));
 BUFx3_ASAP7_75t_SL fopt30326 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(n_23016));
 INVxp67_ASAP7_75t_SL fopt30346 (.A(n_25983),
    .Y(n_23068));
 HB1xp67_ASAP7_75t_SL fopt30526 (.A(n_24169),
    .Y(n_23266));
 HB1xp67_ASAP7_75t_SL fopt30527 (.A(n_18711),
    .Y(n_23268));
 HB1xp67_ASAP7_75t_SL fopt30529 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(n_23272));
 HB1xp67_ASAP7_75t_SL fopt30530 (.A(n_23278),
    .Y(n_23276));
 INVxp67_ASAP7_75t_SL fopt30531 (.A(n_23278),
    .Y(n_23277));
 HB1xp67_ASAP7_75t_SL fopt30533 (.A(n_23280),
    .Y(n_23278));
 HB1xp67_ASAP7_75t_SL fopt30534 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(n_23280));
 INVxp67_ASAP7_75t_SL fopt30535 (.A(n_23291),
    .Y(n_23289));
 INVx1_ASAP7_75t_SL fopt30536 (.A(n_23291),
    .Y(n_23290));
 HB1xp67_ASAP7_75t_SL fopt30537 (.A(n_13566),
    .Y(n_23291));
 INVx2_ASAP7_75t_SL fopt30539 (.A(n_23037),
    .Y(n_23296));
 INVx1_ASAP7_75t_SL fopt30615 (.A(n_23373),
    .Y(n_23374));
 HB1xp67_ASAP7_75t_SL fopt30616 (.A(n_23374),
    .Y(n_23376));
 INVx2_ASAP7_75t_SL fopt30626 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_91),
    .Y(n_21801));
 HB1xp67_ASAP7_75t_SL fopt30643 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .Y(n_23399));
 HB1xp67_ASAP7_75t_SL fopt30705 (.A(n_23463),
    .Y(n_23466));
 INVx2_ASAP7_75t_SL fopt30729 (.A(n_12956),
    .Y(n_23493));
 HB1xp67_ASAP7_75t_SL fopt30730 (.A(n_22610),
    .Y(n_23495));
 HB1xp67_ASAP7_75t_SL fopt30731 (.A(n_20095),
    .Y(n_23497));
 HB1xp67_ASAP7_75t_SL fopt308 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_37),
    .Y(n_7584));
 INVxp67_ASAP7_75t_SL fopt30982 (.A(n_15886),
    .Y(n_23753));
 INVx1_ASAP7_75t_SL fopt31016 (.A(n_23790),
    .Y(n_23789));
 HB1xp67_ASAP7_75t_SL fopt31017 (.A(n_8803),
    .Y(n_23790));
 HB1xp67_ASAP7_75t_SL fopt31245 (.A(n_21949),
    .Y(n_24021));
 INVx1_ASAP7_75t_SL fopt31246 (.A(n_21949),
    .Y(n_24022));
 INVx1_ASAP7_75t_SL fopt31248 (.A(n_24024),
    .Y(n_24025));
 INVxp67_ASAP7_75t_SL fopt313 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120),
    .Y(n_21079));
 INVxp67_ASAP7_75t_SL fopt314 (.A(n_26021),
    .Y(n_20886));
 BUFx6f_ASAP7_75t_SL fopt31526 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_24402));
 INVxp67_ASAP7_75t_SL fopt321 (.A(n_21860),
    .Y(n_21861));
 INVxp67_ASAP7_75t_SL fopt322 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .Y(n_21860));
 INVxp67_ASAP7_75t_SL fopt32221 (.A(n_25132),
    .Y(n_25131));
 HB1xp67_ASAP7_75t_SL fopt32222 (.A(n_19730),
    .Y(n_25132));
 HB1xp67_ASAP7_75t_SL fopt32387 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_154),
    .Y(n_25300));
 INVx1_ASAP7_75t_SL fopt32523 (.A(n_25446),
    .Y(n_25447));
 INVx1_ASAP7_75t_L fopt32662 (.A(n_25604),
    .Y(n_25606));
 INVx1_ASAP7_75t_SL fopt3294 (.A(n_17559),
    .Y(n_12023));
 INVx1_ASAP7_75t_SL fopt3296 (.A(n_12017),
    .Y(n_12035));
 INVxp67_ASAP7_75t_SL fopt33273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_143),
    .Y(n_26266));
 INVx1_ASAP7_75t_SL fopt33274 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_143),
    .Y(n_26267));
 INVx2_ASAP7_75t_SL fopt35 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(n_2836));
 INVxp67_ASAP7_75t_SL fopt357 (.A(n_21841),
    .Y(n_21842));
 INVx1_ASAP7_75t_SL fopt39 (.A(n_14372),
    .Y(n_14373));
 INVxp67_ASAP7_75t_SL fopt4 (.A(n_2293),
    .Y(n_2298));
 INVxp67_ASAP7_75t_SL fopt40 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_29),
    .Y(n_5724));
 BUFx12f_ASAP7_75t_SL fopt41 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[19]),
    .Y(n_22156));
 INVx1_ASAP7_75t_SL fopt42 (.A(n_26258),
    .Y(n_5733));
 INVxp67_ASAP7_75t_SL fopt423 (.A(n_6984),
    .Y(n_6992));
 HB1xp67_ASAP7_75t_SL fopt424 (.A(n_6975),
    .Y(n_6984));
 INVx1_ASAP7_75t_SL fopt4264 (.A(n_23046),
    .Y(n_23060));
 INVx1_ASAP7_75t_SL fopt447 (.A(n_19675),
    .Y(n_19676));
 INVxp67_ASAP7_75t_SL fopt477 (.A(n_19381),
    .Y(n_13606));
 INVxp67_ASAP7_75t_SL fopt49 (.A(n_13464),
    .Y(n_13467));
 INVx2_ASAP7_75t_SL fopt572 (.A(n_14749),
    .Y(n_7297));
 INVx1_ASAP7_75t_SL fopt576 (.A(n_18795),
    .Y(n_14933));
 INVx1_ASAP7_75t_SL fopt579 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_201),
    .Y(n_14931));
 INVx1_ASAP7_75t_L fopt580 (.A(n_12394),
    .Y(n_10318));
 BUFx12f_ASAP7_75t_SL fopt60 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[27]),
    .Y(n_12800));
 INVxp67_ASAP7_75t_SRAM fopt64 (.A(n_20841),
    .Y(n_19989));
 HB1xp67_ASAP7_75t_SL fopt71 (.A(n_21359),
    .Y(n_21276));
 BUFx3_ASAP7_75t_SL fopt77 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_21),
    .Y(n_15003));
 INVxp33_ASAP7_75t_SL fopt86 (.A(n_19429),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_75));
 INVx1_ASAP7_75t_SL fopt916 (.A(n_17979),
    .Y(n_11474));
 INVx1_ASAP7_75t_SL fopt917 (.A(n_21503),
    .Y(n_11473));
 INVx1_ASAP7_75t_SL fopt918 (.A(n_11492),
    .Y(n_11493));
 HB1xp67_ASAP7_75t_SL fopt919 (.A(n_21503),
    .Y(n_11492));
 INVx1_ASAP7_75t_SL fopt92 (.A(n_10173),
    .Y(n_10174));
 HB1xp67_ASAP7_75t_SL fopt94 (.A(n_21389),
    .Y(n_21390));
 HB1xp67_ASAP7_75t_SL g1 (.A(n_7362),
    .Y(n_16070));
 NAND2xp5_ASAP7_75t_SL g10 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .Y(n_12643));
 INVx1_ASAP7_75t_SL g10022 (.A(n_2085),
    .Y(n_2084));
 NAND2xp5_ASAP7_75t_SL g101 (.A(n_5321),
    .B(n_5322),
    .Y(n_5323));
 INVx1_ASAP7_75t_SL g10129 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d2),
    .Y(n_2196));
 INVx1_ASAP7_75t_SL g10139 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d1),
    .Y(n_2191));
 AND2x2_ASAP7_75t_SL g10145__2398 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_797));
 AND2x2_ASAP7_75t_SL g10146__5107 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_582),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_583));
 AND2x2_ASAP7_75t_SL g10148__4319 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_794),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_795));
 AND2x2_ASAP7_75t_SL g10149__8428 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_718),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_719));
 AND2x2_ASAP7_75t_SL g10150__5526 (.A(n_2154),
    .B(n_11587),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_743));
 AND2x2_ASAP7_75t_SL g10151__6783 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_602),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_603));
 AND2x2_ASAP7_75t_SL g10153__1617 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_595));
 AND2x2_ASAP7_75t_SL g10154__2802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_596),
    .B(n_22164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_597));
 AND2x2_ASAP7_75t_SL g10155__1705 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_598),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_599));
 AND2x2_ASAP7_75t_SL g10156__5122 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_600),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_601));
 AND2x2_ASAP7_75t_SL g10157__8246 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_604),
    .B(n_12748),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_605));
 AND2x2_ASAP7_75t_SL g10159__6131 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_602),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_603));
 AND2x2_ASAP7_75t_SL g10160__1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_604),
    .B(n_22164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_605));
 AND2x2_ASAP7_75t_SL g10161__28137 (.A(n_2182),
    .B(n_21595),
    .Y(n_20589));
 AND2x2_ASAP7_75t_SL g10164__30060 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_744),
    .Y(n_22712));
 AND2x2_ASAP7_75t_SL g10166__9945 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_552),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_553));
 AND2x2_ASAP7_75t_SL g10174__5107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_558),
    .B(n_2182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_559));
 AND2x2_ASAP7_75t_SL g10176__4319 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_652),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_653));
 AND2x2_ASAP7_75t_SL g10179__6783 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_560),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_561));
 AND2x2_ASAP7_75t_SL g10180__3680 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_654),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_655));
 AND2x2_ASAP7_75t_SL g10181__1617 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_656),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_657));
 AND2x2_ASAP7_75t_SL g10183__1705 (.A(n_2180),
    .B(n_17672),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_659));
 AND2x2_ASAP7_75t_SL g10184__5122 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_660),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_661));
 AND2x2_ASAP7_75t_SL g10185__8246 (.A(n_2182),
    .B(n_10543),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_565));
 AND2x2_ASAP7_75t_SL g10186__7098 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_663));
 AND2x2_ASAP7_75t_SL g10187__6131 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_664),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_665));
 AND2x2_ASAP7_75t_SL g10188__1881 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_566),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_567));
 AND2x2_ASAP7_75t_SL g10189__5115 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_667));
 AND2x2_ASAP7_75t_SL g10190__7482 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_668),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_669));
 AND2x2_ASAP7_75t_SL g10193__9315 (.A(n_2154),
    .B(n_7179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_757));
 AND2x2_ASAP7_75t_SL g10194__9945 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_568),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_569));
 AND2x2_ASAP7_75t_SL g10195__2883 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_634),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_635));
 AND2x2_ASAP7_75t_SL g10196__2346 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_670),
    .B(n_2180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_671));
 AND2x2_ASAP7_75t_SL g10198__7410 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_570),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_571));
 AND2x2_ASAP7_75t_SL g10199__6417 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_546),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_547));
 NAND2xp5_ASAP7_75t_SL g102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[18]),
    .B(n_17870),
    .Y(n_5322));
 AND2x2_ASAP7_75t_SL g10201__2398 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_572),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_573));
 AND2x2_ASAP7_75t_SL g10204__4319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_574),
    .B(n_2182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_575));
 AND2x2_ASAP7_75t_SL g10205__8428 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_552),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_553));
 AND2x2_ASAP7_75t_SL g10207__6783 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_722),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_723));
 AND2x2_ASAP7_75t_SL g10208__3680 (.A(n_2154),
    .B(n_18825),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_751));
 AND2x2_ASAP7_75t_SL g10211__26368 (.A(n_18578),
    .B(n_18577),
    .Y(n_18579));
 AND2x2_ASAP7_75t_SL g10212__5122 (.A(n_18577),
    .B(n_18896),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_559));
 AND2x2_ASAP7_75t_SL g10213__8246 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_560),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_561));
 AND2x2_ASAP7_75t_SL g10214__7098 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_562),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_563));
 AND2x2_ASAP7_75t_SL g10216__1881 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_564),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_565));
 AND2x2_ASAP7_75t_SL g10217__5115 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_566),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_567));
 AND2x2_ASAP7_75t_SL g10219__4733 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_568),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_569));
 AND2x2_ASAP7_75t_SL g10220__6161 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_570),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_571));
 AND2x2_ASAP7_75t_SL g10221__9315 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_752),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_753));
 AND2x2_ASAP7_75t_SL g10222__9945 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_618),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_619));
 AND2x2_ASAP7_75t_SL g10223__2883 (.A(n_9661),
    .B(n_7903),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_613));
 AND2x2_ASAP7_75t_SL g10224__2346 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_572),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_573));
 AND2x2_ASAP7_75t_SL g10225__1666 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_574),
    .B(n_18577),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_575));
 AND2x2_ASAP7_75t_SL g10228__5477 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_620),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_621));
 AND2x2_ASAP7_75t_SL g10230__5107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_610),
    .B(n_2176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_611));
 AND2x2_ASAP7_75t_SL g10233__8428 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_614),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_615));
 AND2x2_ASAP7_75t_SL g10234__5526 (.A(n_2154),
    .B(n_7172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_755));
 AND2x2_ASAP7_75t_SL g10236__3680 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_620),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_621));
 AND2x2_ASAP7_75t_SL g10239__1705 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_622),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_623));
 AND2x2_ASAP7_75t_SL g10240__5122 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_620),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_621));
 AND2x2_ASAP7_75t_SL g10241__8246 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_622),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_623));
 AND2x2_ASAP7_75t_SL g10242__7098 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_625));
 AND2x2_ASAP7_75t_SL g10243__6131 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_625));
 AND2x2_ASAP7_75t_SL g10244__1881 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_625));
 AND2x2_ASAP7_75t_SL g10245__5115 (.A(n_2176),
    .B(n_14946),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_627));
 AND2x2_ASAP7_75t_SL g10246__7482 (.A(n_9661),
    .B(n_7062),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_627));
 AND2x2_ASAP7_75t_SL g10247__4733 (.A(n_2176),
    .B(n_14950),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_629));
 AND2x2_ASAP7_75t_SL g10248__6161 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_631));
 AND2x2_ASAP7_75t_SL g10250__9945 (.A(n_2179),
    .B(n_6035),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_627));
 AND2x2_ASAP7_75t_SL g10251__30066 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_628),
    .Y(n_22719));
 AND2x2_ASAP7_75t_SL g10252__2346 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_633));
 AND2x2_ASAP7_75t_SL g10253__1666 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_634),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_635));
 AND2x2_ASAP7_75t_SL g10254__7410 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_631));
 AND2x2_ASAP7_75t_SL g10255__6417 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_636),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_637));
 AND2x2_ASAP7_75t_SL g10256__5477 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_638),
    .B(n_2176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_639));
 AND2x2_ASAP7_75t_SL g10258__5107 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_633));
 AND2x2_ASAP7_75t_SL g10259__6260 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_564),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_565));
 AND2x2_ASAP7_75t_SL g10260__4319 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_628),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_629));
 AND2x2_ASAP7_75t_SL g10261__8428 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_724),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_725));
 AND2x2_ASAP7_75t_SL g10262__5526 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_566),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_567));
 AND2x2_ASAP7_75t_SL g10263__6783 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_631));
 AND2x2_ASAP7_75t_SL g10264__3680 (.A(n_9661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_636),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_637));
 AND2x2_ASAP7_75t_SL g10265__1617 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_726),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_727));
 AND2x2_ASAP7_75t_SL g10266__2802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_638),
    .B(n_9661),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_639));
 AND2x2_ASAP7_75t_SL g10267__1705 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_758),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_759));
 AND2x2_ASAP7_75t_SL g10268__5122 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_633));
 AND2x2_ASAP7_75t_SL g10269__8246 (.A(n_6879),
    .B(n_10322),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_737));
 AND2x2_ASAP7_75t_SL g10270__7098 (.A(n_2181),
    .B(n_20656),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_549));
 AND2x2_ASAP7_75t_SL g10271__6131 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_761));
 AND2x2_ASAP7_75t_SL g10272__1881 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_634),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_635));
 AND2x2_ASAP7_75t_SL g10273__5115 (.A(n_6879),
    .B(n_12391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_739));
 AND2x2_ASAP7_75t_SL g10274__7482 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_636),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_637));
 AND2x2_ASAP7_75t_SL g10276__6161 (.A(n_6879),
    .B(n_10319),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_743));
 AND2x2_ASAP7_75t_SL g10277__9315 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_763));
 AND2x2_ASAP7_75t_SL g10278__9945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_638),
    .B(n_2179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_639));
 AND2x2_ASAP7_75t_SL g10281__1666 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_736),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_737));
 AND2x2_ASAP7_75t_SL g10283__6417 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_750),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_751));
 AND2x2_ASAP7_75t_SL g10284__5477 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_752),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_753));
 AND2x2_ASAP7_75t_SL g10285__2398 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_754),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_755));
 AND2x2_ASAP7_75t_SL g10286__5107 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_729));
 AND2x2_ASAP7_75t_SL g10287__6260 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_764),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_765));
 AND2x2_ASAP7_75t_SL g10288__4319 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_756),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_757));
 AND2x2_ASAP7_75t_SL g10289__8428 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_758),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_759));
 AND2x2_ASAP7_75t_SL g10290__5526 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_568),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_569));
 AND2x2_ASAP7_75t_SL g10291__6783 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_730),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_731));
 AND2x2_ASAP7_75t_SL g10292__3680 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_766),
    .B(n_2154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_767));
 AND2x2_ASAP7_75t_SL g10293__1617 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_738),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_739));
 AND2x2_ASAP7_75t_SL g10294__2802 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_761));
 AND2x2_ASAP7_75t_SL g10295__1705 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_763));
 AND2x2_ASAP7_75t_SL g10297__8246 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_764),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_765));
 AND2x2_ASAP7_75t_SL g10298__7098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_766),
    .B(n_6879),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_767));
 INVx1_ASAP7_75t_SL g103 (.A(n_17869),
    .Y(n_5324));
 AND2x2_ASAP7_75t_SL g10302__7482 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_744),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_745));
 AND2x2_ASAP7_75t_SL g10304__6161 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_732),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_733));
 AND2x2_ASAP7_75t_SL g10311__6417 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_750),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_751));
 AND2x2_ASAP7_75t_SL g10313__2398 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_782),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_783));
 AND2x2_ASAP7_75t_SL g10314__5107 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_752),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_753));
 AND2x2_ASAP7_75t_SL g10315__6260 (.A(n_2173),
    .B(n_10369),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_785));
 AND2x2_ASAP7_75t_SL g10316__4319 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_786),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_787));
 AND2x2_ASAP7_75t_SL g10318__5526 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_570),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_571));
 AND2x2_ASAP7_75t_SL g10321__1617 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_754),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_755));
 AND2x2_ASAP7_75t_SL g10322__2802 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_788),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_789));
 AND2x2_ASAP7_75t_SL g10323__1705 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_790),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_791));
 AND2x2_ASAP7_75t_SL g10324__5122 (.A(n_2174),
    .B(n_6962),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_757));
 AND2x2_ASAP7_75t_SL g10325__8246 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_792),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_793));
 AND2x2_ASAP7_75t_SL g10326__7098 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_794),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_795));
 AND2x2_ASAP7_75t_SL g10328__1881 (.A(n_2174),
    .B(n_6964),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_759));
 AND2x2_ASAP7_75t_SL g10329__5115 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_797));
 AND2x2_ASAP7_75t_SL g10330__7482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_798),
    .B(n_2173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_799));
 AND2x2_ASAP7_75t_SL g10331__4733 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_761));
 AND2x2_ASAP7_75t_SL g10335__2883 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_763));
 AND2x2_ASAP7_75t_SL g10337__1666 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_708),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_709));
 AND2x2_ASAP7_75t_SL g10338__7410 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_764),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_765));
 AND2x2_ASAP7_75t_SL g10341__2398 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_776),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_777));
 AND2x2_ASAP7_75t_SL g10342__5107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_766),
    .B(n_2174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_767));
 AND2x2_ASAP7_75t_SL g10347__6783 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_720),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_721));
 AND2x2_ASAP7_75t_SL g10348__3680 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_572),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_573));
 AND2x2_ASAP7_75t_SL g10349__1617 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_778),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_779));
 AND2x2_ASAP7_75t_SL g10350__2802 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_722),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_723));
 AND2x2_ASAP7_75t_SL g10351__1705 (.A(n_20825),
    .B(n_21486),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_725));
 AND2x2_ASAP7_75t_SL g10353__8246 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_729));
 AND2x2_ASAP7_75t_SL g10356__1881 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_730),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_731));
 AND2x2_ASAP7_75t_SL g10357__5115 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_732),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_733));
 AND2x2_ASAP7_75t_SL g10361__9315 (.A(n_21789),
    .B(n_13625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_783));
 AND2x2_ASAP7_75t_SL g10363__2883 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_776),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_777));
 AND2x2_ASAP7_75t_SL g10371__6260 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_682),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_683));
 AND2x2_ASAP7_75t_SL g10372__4319 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_684),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_685));
 AND2x2_ASAP7_75t_SL g10373__8428 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_552),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_553));
 AND2x2_ASAP7_75t_SL g10374__5526 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_574),
    .B(n_2181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_575));
 AND2x2_ASAP7_75t_SL g10375__6783 (.A(n_2169),
    .B(n_20786),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_643));
 AND2x2_ASAP7_75t_SL g10377__1617 (.A(n_14804),
    .B(n_24102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_783));
 AND2x2_ASAP7_75t_SL g10378__2802 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_686),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_687));
 AND2x2_ASAP7_75t_SL g10380__5122 (.A(n_24102),
    .B(n_14806),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_785));
 AND2x2_ASAP7_75t_SL g10381__8246 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_690),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_691));
 AND2x2_ASAP7_75t_SL g10382__7098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_692),
    .B(n_2160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_693));
 AND2x2_ASAP7_75t_SL g10383__6131 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_788),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_789));
 AND2x2_ASAP7_75t_SL g10385__5115 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_695));
 AND2x2_ASAP7_75t_SL g10386__7482 (.A(n_2160),
    .B(n_21413),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_697));
 AND2x2_ASAP7_75t_SL g10387__4733 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_788),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_789));
 AND2x2_ASAP7_75t_SL g10388__6161 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_698),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_699));
 AND2x2_ASAP7_75t_SL g10389__9315 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_700),
    .B(n_2160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_701));
 XNOR2xp5_ASAP7_75t_SL g1039 (.A(n_12492),
    .B(n_12510),
    .Y(n_12511));
 AND2x2_ASAP7_75t_SL g10391__2883 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_790),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_791));
 AND2x2_ASAP7_75t_SL g10392__2346 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_790),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_791));
 AND2x2_ASAP7_75t_SL g10395__6417 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_792),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_793));
 AND2x2_ASAP7_75t_SL g10396__5477 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_578),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_579));
 AND2x2_ASAP7_75t_SL g10397__2398 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_792),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_793));
 INVxp67_ASAP7_75t_SL g104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_5321));
 XNOR2xp5_ASAP7_75t_SL g1040 (.A(n_12091),
    .B(n_24671),
    .Y(n_12101));
 AND2x2_ASAP7_75t_SL g10402__5107 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_593));
 AND2x2_ASAP7_75t_SL g10405__8428 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_646),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_647));
 AND2x2_ASAP7_75t_SL g10406__5526 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_794),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_795));
 AND2x2_ASAP7_75t_SL g10407__6783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_798),
    .B(n_24102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_799));
 AND2x2_ASAP7_75t_SL g10408__3680 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_588),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_589));
 AND2x2_ASAP7_75t_SL g10410__2802 (.A(n_19370),
    .B(n_10139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_705));
 AND2x2_ASAP7_75t_SL g10412__5122 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_595));
 AND2x2_ASAP7_75t_SL g10413__8246 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_797));
 AND2x2_ASAP7_75t_SL g10414__7098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_596),
    .B(n_2168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_597));
 AND2x2_ASAP7_75t_SL g10415__6131 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_598),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_599));
 AND2x2_ASAP7_75t_SL g10417__5115 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_600),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_601));
 AND2x2_ASAP7_75t_SL g10418__7482 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_602),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_603));
 AND2x2_ASAP7_75t_SL g10420__6161 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_798),
    .B(n_21789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_799));
 AND2x2_ASAP7_75t_SL g10422__9945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_604),
    .B(n_2168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_605));
 AND2x2_ASAP7_75t_SL g10427__6417 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_712),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_713));
 AND2x2_ASAP7_75t_SL g10428__5477 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_642),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_643));
 AND2x2_ASAP7_75t_SL g10433__8428 (.A(n_2169),
    .B(n_10044),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_651));
 AND2x2_ASAP7_75t_SL g10434__5526 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_652),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_653));
 AND2x2_ASAP7_75t_SL g10435__6783 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_716),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_717));
 AND2x2_ASAP7_75t_SL g10436__3680 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_718),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_719));
 AND2x2_ASAP7_75t_SL g10437__1617 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_648),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_649));
 AND2x2_ASAP7_75t_SL g10438__2802 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_650),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_651));
 AND2x2_ASAP7_75t_SL g10440__5122 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_654),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_655));
 AND2x2_ASAP7_75t_SL g10443__6131 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_658),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_659));
 AND2x2_ASAP7_75t_SL g10444__1881 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_722),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_723));
 AND2x2_ASAP7_75t_SL g10445__5115 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_660),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_661));
 AND2x2_ASAP7_75t_SL g10446__7482 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_663));
 AND2x2_ASAP7_75t_SL g10448__6161 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_724),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_725));
 AND2x2_ASAP7_75t_SL g10449__9315 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_664),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_665));
 OAI21xp5_ASAP7_75t_SL g1045 (.A1(n_21829),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_285),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_292),
    .Y(n_12110));
 AND2x2_ASAP7_75t_SL g10450__9945 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_667));
 AND2x2_ASAP7_75t_SL g10451__2883 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_726),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_727));
 AND2x2_ASAP7_75t_SL g10452__2346 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_668),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_669));
 AND2x2_ASAP7_75t_SL g10453__1666 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_670),
    .B(n_7595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_671));
 AND2x2_ASAP7_75t_SL g10454__14426 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_676),
    .Y(n_4645));
 AND2x2_ASAP7_75t_SL g10455__6417 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_729));
 AND2x2_ASAP7_75t_SL g10457__2398 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_730),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_731));
 AND2x2_ASAP7_75t_SL g10460__4319 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_654),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_655));
 AND2x2_ASAP7_75t_SL g10462__5526 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_732),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_733));
 AND2x2_ASAP7_75t_SL g10468__30062 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_680),
    .Y(n_22714));
 AND2x2_ASAP7_75t_SL g10469__8246 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_672),
    .B(n_2162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_673));
 OAI21xp5_ASAP7_75t_SL g1047 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_263),
    .A2(n_12975),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_267),
    .Y(n_12108));
 AND2x2_ASAP7_75t_SL g10470__7098 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_558),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_559));
 AND2x2_ASAP7_75t_SL g10471__6131 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_560),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_561));
 AND2x2_ASAP7_75t_SL g10472__1881 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_562),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_563));
 AND2x2_ASAP7_75t_SL g10473__5115 (.A(n_2163),
    .B(n_8306),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_565));
 AND2x2_ASAP7_75t_SL g10474__7482 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_656),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_657));
 AND2x2_ASAP7_75t_SL g10475__4733 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_682),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_683));
 AND2x2_ASAP7_75t_SL g10476__6161 (.A(n_2163),
    .B(n_8311),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_567));
 AND2x2_ASAP7_75t_SL g10477__9315 (.A(n_2163),
    .B(n_10799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_569));
 AND2x2_ASAP7_75t_SL g10478__14706 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_674),
    .Y(n_4957));
 AND2x2_ASAP7_75t_SL g10479__2883 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_570),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_571));
 NOR2xp33_ASAP7_75t_SL g1048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_263),
    .B(n_24669),
    .Y(n_12107));
 AND2x2_ASAP7_75t_SL g10480__2346 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_572),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_573));
 AND2x2_ASAP7_75t_SL g10482__7410 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_676),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_677));
 AND2x2_ASAP7_75t_SL g10483__6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_574),
    .B(n_2163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_575));
 AND2x2_ASAP7_75t_SL g10484__5477 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_608),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_609));
 AND2x2_ASAP7_75t_SL g10488__4319 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_658),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_659));
 AND2x2_ASAP7_75t_SL g10489__8428 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_686),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_687));
 AOI21xp5_ASAP7_75t_SRAM g1049 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266),
    .B(n_19505),
    .Y(n_12492));
 AND2x2_ASAP7_75t_SL g10490__5526 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_680),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_681));
 AND2x2_ASAP7_75t_SL g10495__1705 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_616),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_617));
 AND2x2_ASAP7_75t_SL g10496__5122 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_688),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_689));
 AND2x2_ASAP7_75t_SL g10498__7098 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_618),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_619));
 AND2x2_ASAP7_75t_SL g10500__1881 (.A(n_2162),
    .B(n_19017),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_687));
 AND2x2_ASAP7_75t_SL g10501__5115 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_622),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_623));
 AND2x2_ASAP7_75t_SL g10502__7482 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_625));
 AND2x2_ASAP7_75t_SL g10503__4733 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_660),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_661));
 AND2x2_ASAP7_75t_SL g10504__6161 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_690),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_691));
 AND2x2_ASAP7_75t_SL g10506__9945 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_626),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_627));
 AND2x2_ASAP7_75t_SL g10507__2883 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_628),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_629));
 AND2x2_ASAP7_75t_SL g10508__2346 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_690),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_691));
 AND2x2_ASAP7_75t_SL g10509__1666 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_631));
 AND2x2_ASAP7_75t_SL g10510__7410 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_633));
 AND2x2_ASAP7_75t_SL g10511__6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_692),
    .B(n_2165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_693));
 AND2x2_ASAP7_75t_SL g10512__5477 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_692),
    .B(n_2162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_693));
 AND2x2_ASAP7_75t_SL g10513__2398 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_634),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_635));
 AND2x2_ASAP7_75t_SL g10514__5107 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_636),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_637));
 AND2x2_ASAP7_75t_SL g10515__6260 (.A(n_2162),
    .B(n_17475),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_695));
 AND2x2_ASAP7_75t_SL g10516__4319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_638),
    .B(n_2161),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_639));
 AND2x2_ASAP7_75t_SL g10518__5526 (.A(n_13030),
    .B(n_20238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_709));
 AND2x2_ASAP7_75t_SL g10519__6783 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_663));
 AND2x2_ASAP7_75t_SL g10520__3680 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_695));
 AND2x2_ASAP7_75t_SL g10521__1617 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_696),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_697));
 AND2x2_ASAP7_75t_SL g10522__2802 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_698),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_699));
 AND2x2_ASAP7_75t_SL g10525__8246 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_696),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_697));
 AND2x2_ASAP7_75t_SL g10526__7098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_700),
    .B(n_2162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_701));
 AND2x2_ASAP7_75t_SL g10528__1881 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_744),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_745));
 AND2x2_ASAP7_75t_SL g10530__7482 (.A(n_2151),
    .B(n_10057),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_747));
 AND2x2_ASAP7_75t_SL g10532__6161 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_664),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_665));
 AND2x2_ASAP7_75t_SL g10533__9315 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_698),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_699));
 AND2x2_ASAP7_75t_SL g10535__2883 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_750),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_751));
 AND2x2_ASAP7_75t_SL g10536__2346 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_752),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_753));
 AND2x2_ASAP7_75t_SL g10537__1666 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_754),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_755));
 AND2x2_ASAP7_75t_SL g10538__7410 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_756),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_757));
 AND2x2_ASAP7_75t_SL g10539__6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_700),
    .B(n_2165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_701));
 AND2x2_ASAP7_75t_SL g10541__2398 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_758),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_759));
 AND2x2_ASAP7_75t_SL g10542__5107 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_761));
 AND2x2_ASAP7_75t_SL g10543__6260 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_580),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_581));
 AND2x2_ASAP7_75t_SL g10544__4319 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_763));
 AND2x2_ASAP7_75t_SL g10545__8428 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_764),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_765));
 AND2x2_ASAP7_75t_SL g10546__5526 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_545));
 AND2x2_ASAP7_75t_SL g10547__6783 (.A(n_2181),
    .B(n_23127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_559));
 AND2x2_ASAP7_75t_SL g10548__3680 (.A(n_26221),
    .B(n_13030),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_711));
 AND2x2_ASAP7_75t_SL g10549__1617 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_667));
 AND2x2_ASAP7_75t_SL g10552__5122 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_766),
    .B(n_2151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_767));
 AND2x2_ASAP7_75t_SL g10553__8246 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_768),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_769));
 AND2x2_ASAP7_75t_SL g10554__7098 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_584),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_585));
 AND2x2_ASAP7_75t_SL g10562__9945 (.A(n_2169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_668),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_669));
 AND2x2_ASAP7_75t_SL g10563__2883 (.A(n_2159),
    .B(n_18973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_591));
 AND2x2_ASAP7_75t_SL g10564__2346 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_778),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_779));
 AND2x2_ASAP7_75t_SL g10567__6417 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_782),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_783));
 AND2x2_ASAP7_75t_SL g10568__5477 (.A(n_2158),
    .B(n_7788),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_785));
 AND2x2_ASAP7_75t_SL g10569__2398 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_595));
 AND2x2_ASAP7_75t_SL g10571__6260 (.A(n_2158),
    .B(n_6661),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_789));
 AND2x2_ASAP7_75t_SL g10572__4319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_596),
    .B(n_2159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_597));
 AND2x2_ASAP7_75t_SL g10573__8428 (.A(n_2158),
    .B(n_6666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_791));
 AND2x2_ASAP7_75t_SL g10574__5526 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_792),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_793));
 AND2x2_ASAP7_75t_SL g10575__6783 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_712),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_713));
 AND2x2_ASAP7_75t_SL g10576__3680 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_670),
    .B(n_2169),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_671));
 AND2x2_ASAP7_75t_SL g10578__2802 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_598),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_599));
 AND2x2_ASAP7_75t_SL g10579__1705 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_794),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_795));
 INVx1_ASAP7_75t_SL g1058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_280),
    .Y(n_12091));
 AND2x2_ASAP7_75t_SL g10580__5122 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_797));
 AND2x2_ASAP7_75t_SL g10581__8246 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_600),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_601));
 AND2x2_ASAP7_75t_SL g10582__7098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_798),
    .B(n_2158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_799));
 AND2x2_ASAP7_75t_SL g10583__6131 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_704),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_705));
 AND2x2_ASAP7_75t_SL g10585__5115 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_602),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_603));
 AND2x2_ASAP7_75t_SL g10587__4733 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_604),
    .B(n_2159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_605));
 AND2x2_ASAP7_75t_SL g10588__6161 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_708),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_709));
 AND2x2_ASAP7_75t_SL g10590__9945 (.A(n_2154),
    .B(n_11590),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_737));
 AND2x2_ASAP7_75t_SL g10591__2883 (.A(n_12748),
    .B(n_19145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_583));
 AND2x2_ASAP7_75t_SL g10593__1666 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_712),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_713));
 AND2x2_ASAP7_75t_SL g10596__5477 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_716),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_717));
 AND2x2_ASAP7_75t_SL g10599__6260 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_720),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_721));
 INVx1_ASAP7_75t_SL g106 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_237),
    .Y(n_5582));
 NOR2x1_ASAP7_75t_SL g1060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_283),
    .B(n_19696),
    .Y(n_12494));
 AND2x2_ASAP7_75t_SL g10600__4319 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_722),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_723));
 AND2x2_ASAP7_75t_SL g10601__8428 (.A(n_12781),
    .B(n_7591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_725));
 AND2x2_ASAP7_75t_SL g10602__5526 (.A(n_12781),
    .B(n_7593),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_727));
 AND2x2_ASAP7_75t_SL g10605__1617 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_586),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_587));
 AND2x2_ASAP7_75t_SL g10606__2802 (.A(n_9662),
    .B(n_20328),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_643));
 AND2x2_ASAP7_75t_SL g10607__1705 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_729));
 AND2x2_ASAP7_75t_SL g10608__5122 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_730),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_731));
 AND2x2_ASAP7_75t_SL g10609__8246 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_644),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_645));
 AND2x2_ASAP7_75t_SL g10610__7098 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_732),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_733));
 AND2x2_ASAP7_75t_SL g10613__5115 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_646),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_647));
 AND2x2_ASAP7_75t_SL g10614__7482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_672),
    .B(n_19838),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_673));
 AND2x2_ASAP7_75t_SL g10616__6161 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_674),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_675));
 AND2x2_ASAP7_75t_SL g10617__9315 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_590),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_591));
 AND2x2_ASAP7_75t_SL g10618__9945 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_650),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_651));
 AND2x2_ASAP7_75t_SL g10621__1666 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_652),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_653));
 AND2x2_ASAP7_75t_SL g10622__7410 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_680),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_681));
 AND2x2_ASAP7_75t_SL g10623__6417 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_682),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_683));
 AND2x2_ASAP7_75t_SL g10624__5477 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_593));
 AND2x2_ASAP7_75t_SL g10625__2398 (.A(n_9662),
    .B(n_10039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_655));
 AND2x2_ASAP7_75t_SL g10627__6260 (.A(n_19838),
    .B(n_4779),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_687));
 AND2x2_ASAP7_75t_SL g10628__4319 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_656),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_657));
 AND2x2_ASAP7_75t_SL g10629__8428 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_688),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_689));
 AND2x2_ASAP7_75t_SL g10630__5526 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_690),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_691));
 AND2x2_ASAP7_75t_SL g10632__3680 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_738),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_739));
 AND2x2_ASAP7_75t_SL g10633__1617 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_595));
 AND2x2_ASAP7_75t_SL g10634__2802 (.A(n_9662),
    .B(n_6233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_659));
 AND2x2_ASAP7_75t_SL g10635__1705 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_692),
    .B(n_19838),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_693));
 AND2x2_ASAP7_75t_SL g10636__5122 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_695));
 AND2x2_ASAP7_75t_SL g10637__30067 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_660),
    .Y(n_22720));
 AND2x2_ASAP7_75t_SL g10638__7098 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_696),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_697));
 AND2x2_ASAP7_75t_SL g10639__6131 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_698),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_699));
 AND2x2_ASAP7_75t_SL g10640__1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_596),
    .B(n_12748),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_597));
 AND2x2_ASAP7_75t_SL g10641__5115 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_663));
 AND2x2_ASAP7_75t_SL g10642__7482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_700),
    .B(n_19838),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_701));
 AND2x2_ASAP7_75t_SL g10644__6161 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_664),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_665));
 AND2x2_ASAP7_75t_SL g10645__9315 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_576),
    .B(n_22164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_577));
 AND2x2_ASAP7_75t_SL g10647__2883 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_598),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_599));
 AND2x2_ASAP7_75t_SL g10648__2346 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_667));
 AND2x2_ASAP7_75t_SL g10650__7410 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_580),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_581));
 AND2x2_ASAP7_75t_SL g10651__6417 (.A(n_9662),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_668),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_669));
 AND2x2_ASAP7_75t_SL g10652__5477 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_582),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_583));
 AND2x2_ASAP7_75t_SL g10653__2398 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_584),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_585));
 AND2x2_ASAP7_75t_SL g10654__5107 (.A(n_12748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_600),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_601));
 AND2x2_ASAP7_75t_SL g10655__6260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_670),
    .B(n_9662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_671));
 AND2x2_ASAP7_75t_SL g10656__4319 (.A(n_22164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_586),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_587));
 AND2x2_ASAP7_75t_SL g10659__6783 (.A(n_22164),
    .B(n_4788),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_591));
 AND3x4_ASAP7_75t_SL g10670__1617 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[7]),
    .Y(n_2182));
 AND3x4_ASAP7_75t_SL g10671__2802 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[7]),
    .Y(n_2181));
 AND3x2_ASAP7_75t_SL g10672__1705 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[4]),
    .Y(n_2180));
 AND3x4_ASAP7_75t_L g10673__5122 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[5]),
    .Y(n_2179));
 AND3x2_ASAP7_75t_SL g10674__26366 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[7]),
    .Y(n_18577));
 AND3x1_ASAP7_75t_SL g10675__7098 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[5]),
    .Y(n_2177));
 AND3x4_ASAP7_75t_L g10676__6131 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[5]),
    .Y(n_2176));
 AND3x2_ASAP7_75t_SL g10678__5115 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[0]),
    .Y(n_2174));
 AND3x4_ASAP7_75t_L g10679__7482 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[1]),
    .Y(n_2173));
 AND3x2_ASAP7_75t_SL g10683__9945 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[4]),
    .Y(n_2169));
 NAND3xp33_ASAP7_75t_SL g10684__2883 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[6]),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[8]),
    .C(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .Y(n_2150));
 AND3x2_ASAP7_75t_SL g10685__2346 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[6]),
    .Y(n_2168));
 AND3x2_ASAP7_75t_SL g10688__6417 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[3]),
    .Y(n_2165));
 AND3x4_ASAP7_75t_L g10690__2398 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[7]),
    .Y(n_2163));
 AND3x4_ASAP7_75t_L g10691__5107 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[3]),
    .Y(n_2162));
 AND3x4_ASAP7_75t_SL g10692__6260 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[5]),
    .Y(n_2161));
 AND3x2_ASAP7_75t_SL g10693__4319 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[3]),
    .Y(n_2160));
 AND3x4_ASAP7_75t_L g10694__8428 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[6]),
    .Y(n_2159));
 AND3x4_ASAP7_75t_L g10695__5526 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[1]),
    .Y(n_2158));
 AND3x1_ASAP7_75t_SL g10698__1617 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[4]),
    .Y(n_2155));
 AND3x4_ASAP7_75t_SL g10699__2802 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[0]),
    .Y(n_2154));
 OAI21x1_ASAP7_75t_SL g107 (.A1(n_5512),
    .A2(n_5515),
    .B(n_5516),
    .Y(n_5517));
 AND3x2_ASAP7_75t_L g10702__8246 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[0]),
    .Y(n_2151));
 AND2x2_ASAP7_75t_SL g10712__1881 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_pvld[7]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_pvld[7]),
    .Y(n_2146));
 INVx1_ASAP7_75t_SL g10718 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_end_3520),
    .Y(n_2144));
 NAND2xp5_ASAP7_75t_SL g10727__7482 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_sel[0]),
    .Y(n_2140));
 NAND2xp5_ASAP7_75t_SL g10730__4733 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_stripe_st),
    .Y(n_2139));
 NAND2xp5_ASAP7_75t_SL g10731__6161 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_sel[3]),
    .Y(n_2138));
 NAND2xp5_ASAP7_75t_SL g10732__9315 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_stripe_end),
    .Y(n_2137));
 NAND2xp5_ASAP7_75t_SL g10733__9945 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_sel[1]),
    .Y(n_2136));
 NAND2xp5_ASAP7_75t_SL g10734__2883 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_sel[2]),
    .Y(n_2135));
 OAI21xp5_ASAP7_75t_SL g10738__2346 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[55]),
    .A2(n_335),
    .B(u_NV_NVDLA_cmac_u_reg_req_pvld),
    .Y(u_NV_NVDLA_cmac_u_reg_n_1258));
 INVxp67_ASAP7_75t_SL g10740 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1),
    .Y(n_2133));
 INVxp67_ASAP7_75t_SL g10742 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1),
    .Y(n_2132));
 OA21x2_ASAP7_75t_SRAM g10745__1666 (.A1(test_mode),
    .A2(u_partition_m_reset_sync_reset_synced_rstn_reset_),
    .B(n_2129),
    .Y(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 INVx1_ASAP7_75t_SL g10747 (.A(u_partition_m_reset_sync_reset_synced_rstn_NV_GENERIC_CELL_d0),
    .Y(n_2131));
 OA21x2_ASAP7_75t_SRAM g10749__7410 (.A1(test_mode),
    .A2(dla_reset_rstn),
    .B(n_2129),
    .Y(n_2130));
 NAND2xp33_ASAP7_75t_SL g10750__6417 (.A(test_mode),
    .B(n_2128),
    .Y(n_2129));
 INVxp67_ASAP7_75t_SL g10751 (.A(direct_reset_),
    .Y(n_2128));
 INVx1_ASAP7_75t_SL g10752 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .Y(n_335));
 INVx1_ASAP7_75t_SL g10753 (.A(sc2mac_dat_pvld),
    .Y(n_2126));
 INVx1_ASAP7_75t_SL g10754 (.A(sc2mac_wt_pvld),
    .Y(n_2125));
 INVx1_ASAP7_75t_SL g10756 (.A(dla_reset_rstn),
    .Y(n_2123));
 NOR5xp2_ASAP7_75t_SL g10757__5477 (.A(n_2083),
    .B(u_NV_NVDLA_cmac_u_reg_req_pd[3]),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[6]),
    .D(u_NV_NVDLA_cmac_u_reg_req_pd[5]),
    .E(u_NV_NVDLA_cmac_u_reg_req_pd[4]),
    .Y(n_2085));
 XOR2xp5_ASAP7_75t_SL g108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_114),
    .B(n_5511),
    .Y(n_5512));
 NAND2xp5_ASAP7_75t_SL g109 (.A(n_5513),
    .B(n_5514),
    .Y(n_5516));
 AND2x2_ASAP7_75t_SL g11 (.A(n_8801),
    .B(n_8799),
    .Y(n_17443));
 NOR2xp33_ASAP7_75t_SL g110 (.A(n_5513),
    .B(n_5514),
    .Y(n_5515));
 OR5x1_ASAP7_75t_SL g11039__2398 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[7]),
    .B(u_NV_NVDLA_cmac_u_reg_req_pd[2]),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[9]),
    .D(u_NV_NVDLA_cmac_u_reg_req_pd[8]),
    .E(n_53),
    .Y(n_2083));
 AOI21xp5_ASAP7_75t_SL g11040__5107 (.A1(n_854),
    .A2(u_NV_NVDLA_cmac_u_core_wt1_actv_pvld[7]),
    .B(n_817),
    .Y(n_2082));
 AOI21xp5_ASAP7_75t_SL g11041__6260 (.A1(n_854),
    .A2(u_NV_NVDLA_cmac_u_core_wt2_actv_pvld[7]),
    .B(n_579),
    .Y(n_2081));
 AOI21xp5_ASAP7_75t_SL g11042__4319 (.A1(n_854),
    .A2(u_NV_NVDLA_cmac_u_core_wt0_actv_pvld[7]),
    .B(n_819),
    .Y(n_2080));
 AOI22xp5_ASAP7_75t_SL g11043__8428 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[0]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .B2(n_823),
    .Y(n_2079));
 AOI22xp5_ASAP7_75t_SL g11044__5526 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[1]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .B2(n_823),
    .Y(n_2078));
 AOI22xp5_ASAP7_75t_SL g11045__6783 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[2]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .B2(n_823),
    .Y(n_2077));
 AOI22xp5_ASAP7_75t_SL g11046__3680 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[3]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .B2(n_823),
    .Y(n_2076));
 AOI22xp5_ASAP7_75t_SL g11047__1617 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[4]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .B2(n_823),
    .Y(n_2075));
 AOI22xp5_ASAP7_75t_SL g11048__2802 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[5]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .B2(n_823),
    .Y(n_2074));
 AOI22xp5_ASAP7_75t_SL g11049__1705 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[6]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .B2(n_823),
    .Y(n_2073));
 AOI21xp5_ASAP7_75t_SL g1105 (.A1(n_22512),
    .A2(n_7051),
    .B(n_7063),
    .Y(n_7064));
 AOI22xp5_ASAP7_75t_SL g11050__5122 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_mask[7]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .B2(n_823),
    .Y(n_2072));
 AOI22xp5_ASAP7_75t_SL g11051__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[0]),
    .A2(n_586),
    .B1(sc2mac_wt_sel[0]),
    .B2(n_585),
    .Y(n_2071));
 AOI22xp5_ASAP7_75t_SL g11052__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[1]),
    .A2(n_586),
    .B1(sc2mac_wt_sel[1]),
    .B2(n_585),
    .Y(n_2070));
 AOI22xp5_ASAP7_75t_SL g11053__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[2]),
    .A2(n_586),
    .B1(sc2mac_wt_sel[2]),
    .B2(n_585),
    .Y(n_2069));
 AOI22xp5_ASAP7_75t_SL g11054__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[3]),
    .A2(n_586),
    .B1(sc2mac_wt_sel[3]),
    .B2(n_585),
    .Y(n_2068));
 AOI22xp5_ASAP7_75t_SL g11055__5115 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_sel[0]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[0]),
    .B2(n_823),
    .Y(n_2067));
 AOI22xp5_ASAP7_75t_SL g11056__7482 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_sel[1]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[1]),
    .B2(n_823),
    .Y(n_2066));
 AOI22xp5_ASAP7_75t_SL g11057__4733 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_sel[2]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[2]),
    .B2(n_823),
    .Y(n_2065));
 AOI22xp5_ASAP7_75t_SL g11058__6161 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_sel[3]),
    .A2(n_824),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[3]),
    .B2(n_823),
    .Y(n_2064));
 AOI22xp5_ASAP7_75t_SL g11059__9315 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[0]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .B2(n_821),
    .Y(n_2063));
 XNOR2xp5_ASAP7_75t_SL g1106 (.A(n_7061),
    .B(n_22512),
    .Y(n_7062));
 AOI22xp5_ASAP7_75t_SL g11060__9945 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[1]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .B2(n_821),
    .Y(n_2062));
 AOI22xp5_ASAP7_75t_SL g11061__2883 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[2]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .B2(n_821),
    .Y(n_2061));
 AOI22xp5_ASAP7_75t_SL g11062__2346 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[3]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .B2(n_821),
    .Y(n_2060));
 AOI22xp5_ASAP7_75t_SL g11063__1666 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[4]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .B2(n_821),
    .Y(n_2059));
 AOI22xp5_ASAP7_75t_SL g11064__7410 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[5]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .B2(n_821),
    .Y(n_2058));
 AOI22xp5_ASAP7_75t_SL g11065__6417 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[6]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .B2(n_821),
    .Y(n_2057));
 AOI22xp5_ASAP7_75t_SL g11066__5477 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_mask[7]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .B2(n_821),
    .Y(n_2056));
 AOI22xp5_ASAP7_75t_SL g11067__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[0]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[0]),
    .B2(n_583),
    .Y(n_2055));
 AOI22xp5_ASAP7_75t_SL g11068__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[1]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[1]),
    .B2(n_583),
    .Y(n_2054));
 AOI22xp5_ASAP7_75t_SL g11069__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[2]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[2]),
    .B2(n_583),
    .Y(n_2053));
 AOI22xp5_ASAP7_75t_SL g11070__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[3]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[3]),
    .B2(n_583),
    .Y(n_2052));
 AOI22xp5_ASAP7_75t_SL g11071__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[4]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[4]),
    .B2(n_583),
    .Y(n_2051));
 AOI22xp5_ASAP7_75t_SL g11072__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[5]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[5]),
    .B2(n_583),
    .Y(n_2050));
 AOI22xp5_ASAP7_75t_SL g11073__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[6]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[6]),
    .B2(n_583),
    .Y(n_2049));
 AOI22xp5_ASAP7_75t_SL g11074__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[7]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[7]),
    .B2(n_583),
    .Y(n_2048));
 AOI22xp5_ASAP7_75t_SL g11075__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[8]),
    .A2(n_584),
    .B1(sc2mac_dat_pd[8]),
    .B2(n_583),
    .Y(n_2047));
 AOI22xp5_ASAP7_75t_SL g11076__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[0]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[0]),
    .B2(n_821),
    .Y(n_2046));
 AOI22xp5_ASAP7_75t_SL g11077__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[1]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[1]),
    .B2(n_821),
    .Y(n_2045));
 AOI22xp5_ASAP7_75t_SL g11078__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[2]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[2]),
    .B2(n_821),
    .Y(n_2044));
 AOI22xp5_ASAP7_75t_SL g11079__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[3]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[3]),
    .B2(n_821),
    .Y(n_2043));
 AOI22xp5_ASAP7_75t_SL g11080__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[4]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[4]),
    .B2(n_821),
    .Y(n_2042));
 AOI22xp5_ASAP7_75t_SL g11081__6131 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_stripe_st),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[5]),
    .B2(n_821),
    .Y(n_2041));
 AOI22xp5_ASAP7_75t_SL g11082__1881 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_stripe_end),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[6]),
    .B2(n_821),
    .Y(n_2040));
 AOI22xp5_ASAP7_75t_SL g11083__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[7]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[7]),
    .B2(n_821),
    .Y(n_2039));
 AOI22xp5_ASAP7_75t_SL g11084__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[8]),
    .A2(n_822),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[8]),
    .B2(n_821),
    .Y(n_2038));
 AOI21xp5_ASAP7_75t_SL g11085__4733 (.A1(u_NV_NVDLA_cmac_u_reg_n_1258),
    .A2(cmac_a2csb_resp_pd[33]),
    .B(n_4416),
    .Y(n_2037));
 OAI33xp33_ASAP7_75t_SL g11090__2346 (.A1(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .A2(n_662),
    .A3(n_338),
    .B1(n_336),
    .B2(n_332),
    .B3(n_333),
    .Y(n_2032));
 AOI22xp5_ASAP7_75t_SL g11091__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[0]),
    .B2(n_582),
    .Y(n_2031));
 AOI22xp5_ASAP7_75t_SL g11092__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[1]),
    .B2(n_582),
    .Y(n_2030));
 AOI22xp5_ASAP7_75t_SL g11093__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[2]),
    .B2(n_582),
    .Y(n_2029));
 AOI22xp5_ASAP7_75t_SL g11094__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[3]),
    .B2(n_582),
    .Y(n_2028));
 AOI22xp5_ASAP7_75t_SL g11095__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[4]),
    .B2(n_582),
    .Y(n_2027));
 AOI22xp5_ASAP7_75t_SL g11096__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[5]),
    .B2(n_582),
    .Y(n_2026));
 AOI22xp5_ASAP7_75t_SL g11097__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[6]),
    .B2(n_582),
    .Y(n_2025));
 AOI22xp5_ASAP7_75t_SL g11098__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .A2(n_581),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[7]),
    .B2(n_582),
    .Y(n_2024));
 AOI22xp5_ASAP7_75t_SL g11099__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[0]),
    .B2(n_17240),
    .Y(n_2023));
 INVx1_ASAP7_75t_SL g111 (.A(n_18927),
    .Y(n_5513));
 NAND3x1_ASAP7_75t_SL g1110 (.A(n_7049),
    .B(n_22512),
    .C(n_7051),
    .Y(n_7052));
 AOI22xp5_ASAP7_75t_SL g11100__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[1]),
    .B2(n_17240),
    .Y(n_2022));
 AOI22xp5_ASAP7_75t_SL g11101__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[2]),
    .B2(n_17240),
    .Y(n_2021));
 AOI22xp5_ASAP7_75t_SL g11102__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[3]),
    .B2(n_17240),
    .Y(n_2020));
 AOI22xp5_ASAP7_75t_SL g11103__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[4]),
    .B2(n_17240),
    .Y(n_2019));
 AOI22xp5_ASAP7_75t_SL g11104__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[5]),
    .B2(n_17240),
    .Y(n_2018));
 AOI22xp5_ASAP7_75t_SL g11105__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[6]),
    .B2(n_17240),
    .Y(n_2017));
 AOI22xp5_ASAP7_75t_SL g11106__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .A2(n_817),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[7]),
    .B2(n_17240),
    .Y(n_2016));
 AOI22xp5_ASAP7_75t_SL g11107__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[0]),
    .B2(n_580),
    .Y(n_2015));
 AOI22xp5_ASAP7_75t_SL g11108__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[1]),
    .B2(n_580),
    .Y(n_2014));
 AOI22xp5_ASAP7_75t_SL g11109__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[2]),
    .B2(n_580),
    .Y(n_2013));
 AND2x2_ASAP7_75t_SL g1111 (.A(n_7049),
    .B(n_23021),
    .Y(n_7060));
 AOI22xp5_ASAP7_75t_SL g11110__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[3]),
    .B2(n_580),
    .Y(n_2012));
 AOI22xp5_ASAP7_75t_SL g11111__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[4]),
    .B2(n_580),
    .Y(n_2011));
 AOI22xp5_ASAP7_75t_SL g11112__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[5]),
    .B2(n_580),
    .Y(n_2010));
 AOI22xp5_ASAP7_75t_SL g11113__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[6]),
    .B2(n_580),
    .Y(n_2009));
 AOI22xp5_ASAP7_75t_SL g11114__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .A2(n_579),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[7]),
    .B2(n_580),
    .Y(n_2008));
 AOI22xp5_ASAP7_75t_SL g11115__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[0]),
    .B2(n_820),
    .Y(n_2007));
 AOI22xp5_ASAP7_75t_SL g11116__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[1]),
    .B2(n_820),
    .Y(n_2006));
 AOI22xp5_ASAP7_75t_SL g11117__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[2]),
    .B2(n_820),
    .Y(n_2005));
 AOI22xp5_ASAP7_75t_SL g11118__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[3]),
    .B2(n_820),
    .Y(n_2004));
 AOI22xp5_ASAP7_75t_SL g11119__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[4]),
    .B2(n_820),
    .Y(n_2003));
 NAND2xp5_ASAP7_75t_SL g1112 (.A(n_7051),
    .B(n_7053),
    .Y(n_7061));
 AOI22xp5_ASAP7_75t_SL g11120__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[5]),
    .B2(n_820),
    .Y(n_2002));
 AOI22xp5_ASAP7_75t_SL g11121__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[6]),
    .B2(n_820),
    .Y(n_2001));
 AOI22xp5_ASAP7_75t_SL g11122__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .A2(n_819),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[7]),
    .B2(n_820),
    .Y(n_2000));
 AOI22xp5_ASAP7_75t_SL g11123__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[6]),
    .B2(n_620),
    .Y(n_1999));
 AOI22xp5_ASAP7_75t_SL g11124__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[7]),
    .B2(n_620),
    .Y(n_1998));
 AOI22xp5_ASAP7_75t_SL g11125__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[8]),
    .B2(n_646),
    .Y(n_1997));
 AOI22xp5_ASAP7_75t_SL g11126__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[9]),
    .B2(n_646),
    .Y(n_1996));
 AOI22xp5_ASAP7_75t_SL g11127__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[10]),
    .B2(n_646),
    .Y(n_1995));
 AOI22xp5_ASAP7_75t_SL g11128__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[11]),
    .B2(n_646),
    .Y(n_1994));
 AOI22xp5_ASAP7_75t_SL g11129__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[12]),
    .B2(n_646),
    .Y(n_1993));
 AOI22xp5_ASAP7_75t_SL g11130__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[14]),
    .B2(n_646),
    .Y(n_1992));
 AOI22xp5_ASAP7_75t_SL g11131__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[13]),
    .B2(n_646),
    .Y(n_1991));
 AOI22xp5_ASAP7_75t_SL g11132__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]),
    .A2(n_645),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[15]),
    .B2(n_646),
    .Y(n_1990));
 AOI22xp5_ASAP7_75t_SL g11133__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[16]),
    .B2(n_598),
    .Y(n_1989));
 AOI22xp5_ASAP7_75t_SL g11134__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[17]),
    .B2(n_598),
    .Y(n_1988));
 AOI22xp5_ASAP7_75t_SL g11135__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[18]),
    .B2(n_598),
    .Y(n_1987));
 AOI22xp5_ASAP7_75t_SL g11136__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[20]),
    .B2(n_598),
    .Y(n_1986));
 AOI22xp5_ASAP7_75t_SL g11137__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[19]),
    .B2(n_598),
    .Y(n_1985));
 AOI22xp5_ASAP7_75t_SL g11138__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[21]),
    .B2(n_598),
    .Y(n_1984));
 AOI22xp5_ASAP7_75t_SL g11139__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[22]),
    .B2(n_598),
    .Y(n_1983));
 INVx2_ASAP7_75t_SL g1114 (.A(n_11781),
    .Y(n_7049));
 AOI22xp5_ASAP7_75t_SL g11140__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]),
    .A2(n_597),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[23]),
    .B2(n_598),
    .Y(n_1982));
 AOI22xp5_ASAP7_75t_SL g11141__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[0]),
    .B2(n_650),
    .Y(n_1981));
 AOI22xp5_ASAP7_75t_SL g11142__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[1]),
    .B2(n_650),
    .Y(n_1980));
 AOI22xp5_ASAP7_75t_SL g11143__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[24]),
    .B2(n_648),
    .Y(n_1979));
 AOI22xp5_ASAP7_75t_SL g11144__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[2]),
    .B2(n_650),
    .Y(n_1978));
 AOI22xp5_ASAP7_75t_SL g11145__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[3]),
    .B2(n_650),
    .Y(n_1977));
 AOI22xp5_ASAP7_75t_SL g11146__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[4]),
    .B2(n_650),
    .Y(n_1976));
 AOI22xp5_ASAP7_75t_SL g11147__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[5]),
    .B2(n_650),
    .Y(n_1975));
 AOI22xp5_ASAP7_75t_SL g11148__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[6]),
    .B2(n_650),
    .Y(n_1974));
 AOI22xp5_ASAP7_75t_SL g11149__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]),
    .A2(n_649),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[7]),
    .B2(n_650),
    .Y(n_1973));
 AOI22xp5_ASAP7_75t_SL g11150__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[25]),
    .B2(n_648),
    .Y(n_1972));
 AOI22xp5_ASAP7_75t_SL g11151__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[26]),
    .B2(n_648),
    .Y(n_1971));
 AOI22xp5_ASAP7_75t_SL g11152__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[8]),
    .B2(n_644),
    .Y(n_1970));
 AOI22xp5_ASAP7_75t_SL g11153__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[9]),
    .B2(n_644),
    .Y(n_1969));
 AOI22xp5_ASAP7_75t_SL g11154__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[27]),
    .B2(n_648),
    .Y(n_1968));
 AOI22xp5_ASAP7_75t_SL g11155__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[10]),
    .B2(n_644),
    .Y(n_1967));
 AOI22xp5_ASAP7_75t_SL g11156__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[11]),
    .B2(n_644),
    .Y(n_1966));
 AOI22xp5_ASAP7_75t_SL g11157__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[12]),
    .B2(n_644),
    .Y(n_1965));
 AOI22xp5_ASAP7_75t_SL g11158__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[28]),
    .B2(n_648),
    .Y(n_1964));
 AOI22xp5_ASAP7_75t_SL g11159__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[13]),
    .B2(n_644),
    .Y(n_1963));
 AOI22xp5_ASAP7_75t_SL g11160__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[14]),
    .B2(n_644),
    .Y(n_1962));
 AOI22xp5_ASAP7_75t_SL g11161__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]),
    .A2(n_643),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[15]),
    .B2(n_644),
    .Y(n_1961));
 AOI22xp5_ASAP7_75t_SL g11162__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[29]),
    .B2(n_648),
    .Y(n_1960));
 AOI22xp5_ASAP7_75t_SL g11163__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[16]),
    .B2(n_642),
    .Y(n_1959));
 AOI22xp5_ASAP7_75t_SL g11164__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[17]),
    .B2(n_642),
    .Y(n_1958));
 AOI22xp5_ASAP7_75t_SL g11165__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[18]),
    .B2(n_642),
    .Y(n_1957));
 AOI22xp5_ASAP7_75t_SL g11166__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[30]),
    .B2(n_648),
    .Y(n_1956));
 AOI22xp5_ASAP7_75t_SL g11167__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[19]),
    .B2(n_642),
    .Y(n_1955));
 AOI22xp5_ASAP7_75t_SL g11168__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[20]),
    .B2(n_642),
    .Y(n_1954));
 AOI22xp5_ASAP7_75t_SL g11169__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]),
    .A2(n_647),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[31]),
    .B2(n_648),
    .Y(n_1953));
 NAND2xp5_ASAP7_75t_SL g1117 (.A(n_11510),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_245),
    .Y(n_7051));
 AOI22xp5_ASAP7_75t_SL g11170__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[32]),
    .B2(n_640),
    .Y(n_1952));
 AOI22xp5_ASAP7_75t_SL g11171__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[21]),
    .B2(n_642),
    .Y(n_1951));
 AOI22xp5_ASAP7_75t_SL g11172__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[22]),
    .B2(n_642),
    .Y(n_1950));
 AOI22xp5_ASAP7_75t_SL g11173__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]),
    .A2(n_641),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[23]),
    .B2(n_642),
    .Y(n_1949));
 AOI22xp5_ASAP7_75t_SL g11174__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[24]),
    .B2(n_638),
    .Y(n_1948));
 AOI22xp5_ASAP7_75t_SL g11175__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[25]),
    .B2(n_638),
    .Y(n_1947));
 AOI22xp5_ASAP7_75t_SL g11176__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[26]),
    .B2(n_638),
    .Y(n_1946));
 AOI22xp5_ASAP7_75t_SL g11177__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[33]),
    .B2(n_640),
    .Y(n_1945));
 AOI22xp5_ASAP7_75t_SL g11178__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[27]),
    .B2(n_638),
    .Y(n_1944));
 AOI22xp5_ASAP7_75t_SL g11179__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[34]),
    .B2(n_640),
    .Y(n_1943));
 INVxp67_ASAP7_75t_SL g1118 (.A(n_7053),
    .Y(n_7063));
 AOI22xp5_ASAP7_75t_SL g11180__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[28]),
    .B2(n_638),
    .Y(n_1942));
 AOI22xp5_ASAP7_75t_SL g11181__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[29]),
    .B2(n_638),
    .Y(n_1941));
 AOI22xp5_ASAP7_75t_SL g11182__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[30]),
    .B2(n_638),
    .Y(n_1940));
 AOI22xp5_ASAP7_75t_SL g11183__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[35]),
    .B2(n_640),
    .Y(n_1939));
 AOI22xp5_ASAP7_75t_SL g11184__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]),
    .A2(n_637),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[31]),
    .B2(n_638),
    .Y(n_1938));
 AOI22xp5_ASAP7_75t_SL g11185__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[32]),
    .B2(n_634),
    .Y(n_1937));
 AOI22xp5_ASAP7_75t_SL g11186__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[36]),
    .B2(n_640),
    .Y(n_1936));
 AOI22xp5_ASAP7_75t_SL g11187__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[33]),
    .B2(n_634),
    .Y(n_1935));
 AOI22xp5_ASAP7_75t_SL g11188__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[34]),
    .B2(n_634),
    .Y(n_1934));
 AOI22xp5_ASAP7_75t_SL g11189__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[35]),
    .B2(n_634),
    .Y(n_1933));
 OR2x2_ASAP7_75t_SL g1119 (.A(n_11510),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_245),
    .Y(n_7053));
 AOI22xp5_ASAP7_75t_SL g11190__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[37]),
    .B2(n_640),
    .Y(n_1932));
 AOI22xp5_ASAP7_75t_SL g11191__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[36]),
    .B2(n_634),
    .Y(n_1931));
 AOI22xp5_ASAP7_75t_SL g11192__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[38]),
    .B2(n_640),
    .Y(n_1930));
 AOI22xp5_ASAP7_75t_SL g11193__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[37]),
    .B2(n_634),
    .Y(n_1929));
 AOI22xp5_ASAP7_75t_SL g11194__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[38]),
    .B2(n_634),
    .Y(n_1928));
 AOI22xp5_ASAP7_75t_SL g11195__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]),
    .A2(n_633),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[39]),
    .B2(n_634),
    .Y(n_1927));
 AOI22xp5_ASAP7_75t_SL g11196__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[40]),
    .B2(n_632),
    .Y(n_1926));
 AOI22xp5_ASAP7_75t_SL g11197__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[41]),
    .B2(n_632),
    .Y(n_1925));
 AOI22xp5_ASAP7_75t_SL g11198__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[42]),
    .B2(n_632),
    .Y(n_1924));
 AOI22xp5_ASAP7_75t_SL g11199__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]),
    .A2(n_639),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[39]),
    .B2(n_640),
    .Y(n_1923));
 INVx2_ASAP7_75t_SL g112 (.A(n_9464),
    .Y(n_5514));
 AOI22xp5_ASAP7_75t_SL g11200__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[40]),
    .B2(n_630),
    .Y(n_1922));
 AOI22xp5_ASAP7_75t_SL g11201__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[43]),
    .B2(n_632),
    .Y(n_1921));
 AOI22xp5_ASAP7_75t_SL g11202__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[44]),
    .B2(n_632),
    .Y(n_1920));
 AOI22xp5_ASAP7_75t_SL g11203__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[45]),
    .B2(n_632),
    .Y(n_1919));
 AOI22xp5_ASAP7_75t_SL g11204__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[46]),
    .B2(n_632),
    .Y(n_1918));
 AOI22xp5_ASAP7_75t_SL g11205__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[41]),
    .B2(n_630),
    .Y(n_1917));
 AOI22xp5_ASAP7_75t_SL g11206__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]),
    .A2(n_631),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[47]),
    .B2(n_632),
    .Y(n_1916));
 AOI22xp5_ASAP7_75t_SL g11207__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[48]),
    .B2(n_628),
    .Y(n_1915));
 AOI22xp5_ASAP7_75t_SL g11208__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[49]),
    .B2(n_628),
    .Y(n_1914));
 AOI22xp5_ASAP7_75t_SL g11209__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[42]),
    .B2(n_630),
    .Y(n_1913));
 AOI22xp5_ASAP7_75t_SL g11210__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[50]),
    .B2(n_628),
    .Y(n_1912));
 AOI22xp5_ASAP7_75t_SL g11211__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[51]),
    .B2(n_628),
    .Y(n_1911));
 AOI22xp5_ASAP7_75t_SL g11212__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[43]),
    .B2(n_630),
    .Y(n_1910));
 AOI22xp5_ASAP7_75t_SL g11213__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[44]),
    .B2(n_630),
    .Y(n_1909));
 AOI22xp5_ASAP7_75t_SL g11214__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[52]),
    .B2(n_628),
    .Y(n_1908));
 AOI22xp5_ASAP7_75t_SL g11215__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[53]),
    .B2(n_628),
    .Y(n_1907));
 AOI22xp5_ASAP7_75t_SL g11216__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[54]),
    .B2(n_628),
    .Y(n_1906));
 AOI22xp5_ASAP7_75t_SL g11217__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]),
    .A2(n_627),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[55]),
    .B2(n_628),
    .Y(n_1905));
 AOI22xp5_ASAP7_75t_SL g11218__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[56]),
    .B2(n_616),
    .Y(n_1904));
 AOI22xp5_ASAP7_75t_SL g11219__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[57]),
    .B2(n_616),
    .Y(n_1903));
 AOI22xp5_ASAP7_75t_SL g11220__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[45]),
    .B2(n_630),
    .Y(n_1902));
 AOI22xp5_ASAP7_75t_SL g11221__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[46]),
    .B2(n_630),
    .Y(n_1901));
 AOI22xp5_ASAP7_75t_SL g11222__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[58]),
    .B2(n_616),
    .Y(n_1900));
 AOI22xp5_ASAP7_75t_SL g11223__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[59]),
    .B2(n_616),
    .Y(n_1899));
 AOI22xp5_ASAP7_75t_SL g11224__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]),
    .A2(n_629),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[47]),
    .B2(n_630),
    .Y(n_1898));
 AOI22xp5_ASAP7_75t_SL g11225__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[60]),
    .B2(n_616),
    .Y(n_1897));
 AOI22xp5_ASAP7_75t_SL g11226__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[61]),
    .B2(n_616),
    .Y(n_1896));
 AOI22xp5_ASAP7_75t_SL g11227__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[62]),
    .B2(n_616),
    .Y(n_1895));
 AOI22xp5_ASAP7_75t_SL g11228__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[48]),
    .B2(n_600),
    .Y(n_1894));
 AOI22xp5_ASAP7_75t_SL g11229__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]),
    .A2(n_615),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[63]),
    .B2(n_616),
    .Y(n_1893));
 AOI22xp5_ASAP7_75t_SL g11230__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[49]),
    .B2(n_600),
    .Y(n_1892));
 AOI22xp5_ASAP7_75t_SL g11231__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[50]),
    .B2(n_600),
    .Y(n_1891));
 AOI22xp5_ASAP7_75t_SL g11232__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[52]),
    .B2(n_600),
    .Y(n_1890));
 AOI22xp5_ASAP7_75t_SL g11233__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[51]),
    .B2(n_600),
    .Y(n_1889));
 AOI22xp5_ASAP7_75t_SL g11234__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[53]),
    .B2(n_600),
    .Y(n_1888));
 AOI22xp5_ASAP7_75t_SL g11235__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[54]),
    .B2(n_600),
    .Y(n_1887));
 AOI22xp5_ASAP7_75t_SL g11236__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[56]),
    .B2(n_623),
    .Y(n_1886));
 AOI22xp5_ASAP7_75t_SL g11237__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]),
    .A2(n_599),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[55]),
    .B2(n_600),
    .Y(n_1885));
 AOI22xp5_ASAP7_75t_SL g11238__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[57]),
    .B2(n_623),
    .Y(n_1884));
 AOI22xp5_ASAP7_75t_SL g11239__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[58]),
    .B2(n_623),
    .Y(n_1883));
 AOI22xp5_ASAP7_75t_SL g11240__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[59]),
    .B2(n_623),
    .Y(n_1882));
 AOI22xp5_ASAP7_75t_SL g11241__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[60]),
    .B2(n_623),
    .Y(n_1881));
 AOI22xp5_ASAP7_75t_SL g11242__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[61]),
    .B2(n_623),
    .Y(n_1880));
 AOI22xp5_ASAP7_75t_SL g11243__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[62]),
    .B2(n_623),
    .Y(n_1879));
 AOI22xp5_ASAP7_75t_SL g11244__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]),
    .A2(n_622),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[63]),
    .B2(n_623),
    .Y(n_1878));
 AOI22xp5_ASAP7_75t_SL g11245__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[0]),
    .B2(n_614),
    .Y(n_1877));
 AOI22xp5_ASAP7_75t_SL g11246__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[1]),
    .B2(n_614),
    .Y(n_1876));
 AOI22xp5_ASAP7_75t_SL g11247__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[2]),
    .B2(n_614),
    .Y(n_1875));
 AOI22xp5_ASAP7_75t_SL g11248__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[3]),
    .B2(n_614),
    .Y(n_1874));
 AOI22xp5_ASAP7_75t_SL g11249__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[4]),
    .B2(n_614),
    .Y(n_1873));
 XNOR2xp5_ASAP7_75t_SL g1125 (.A(n_20640),
    .B(n_23128),
    .Y(n_20656));
 AOI22xp5_ASAP7_75t_SL g11250__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[5]),
    .B2(n_614),
    .Y(n_1872));
 AOI22xp5_ASAP7_75t_SL g11251__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[6]),
    .B2(n_614),
    .Y(n_1871));
 AOI22xp5_ASAP7_75t_SL g11252__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]),
    .A2(n_613),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[7]),
    .B2(n_614),
    .Y(n_1870));
 AOI22xp5_ASAP7_75t_SL g11253__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[8]),
    .B2(n_612),
    .Y(n_1869));
 AOI22xp5_ASAP7_75t_SL g11254__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[9]),
    .B2(n_612),
    .Y(n_1868));
 AOI22xp5_ASAP7_75t_SL g11255__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[10]),
    .B2(n_612),
    .Y(n_1867));
 AOI22xp5_ASAP7_75t_SL g11256__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[11]),
    .B2(n_612),
    .Y(n_1866));
 AOI22xp5_ASAP7_75t_SL g11257__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[12]),
    .B2(n_612),
    .Y(n_1865));
 AOI22xp5_ASAP7_75t_SL g11258__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[13]),
    .B2(n_612),
    .Y(n_1864));
 AOI22xp5_ASAP7_75t_SL g11259__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[14]),
    .B2(n_612),
    .Y(n_1863));
 AOI22xp5_ASAP7_75t_SL g11260__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]),
    .A2(n_611),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[15]),
    .B2(n_612),
    .Y(n_1862));
 AOI22xp5_ASAP7_75t_SL g11261__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[16]),
    .B2(n_610),
    .Y(n_1861));
 AOI22xp5_ASAP7_75t_SL g11262__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[17]),
    .B2(n_610),
    .Y(n_1860));
 AOI22xp5_ASAP7_75t_SL g11263__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[18]),
    .B2(n_610),
    .Y(n_1859));
 AOI22xp5_ASAP7_75t_SL g11264__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[19]),
    .B2(n_610),
    .Y(n_1858));
 AOI22xp5_ASAP7_75t_SL g11265__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[20]),
    .B2(n_610),
    .Y(n_1857));
 AOI22xp5_ASAP7_75t_SL g11266__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[21]),
    .B2(n_610),
    .Y(n_1856));
 AOI22xp5_ASAP7_75t_SL g11267__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[22]),
    .B2(n_610),
    .Y(n_1855));
 AOI22xp5_ASAP7_75t_SL g11268__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]),
    .A2(n_609),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[23]),
    .B2(n_610),
    .Y(n_1854));
 AOI22xp5_ASAP7_75t_SL g11269__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[24]),
    .B2(n_625),
    .Y(n_1853));
 AOI21xp5_ASAP7_75t_SL g1127 (.A1(n_18168),
    .A2(n_6024),
    .B(n_6032),
    .Y(n_6033));
 AOI22xp5_ASAP7_75t_SL g11270__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[25]),
    .B2(n_625),
    .Y(n_1852));
 AOI22xp5_ASAP7_75t_SL g11271__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[26]),
    .B2(n_625),
    .Y(n_1851));
 AOI22xp5_ASAP7_75t_SL g11272__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[27]),
    .B2(n_625),
    .Y(n_1850));
 AOI22xp5_ASAP7_75t_SL g11273__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[28]),
    .B2(n_625),
    .Y(n_1849));
 AOI22xp5_ASAP7_75t_SL g11274__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[29]),
    .B2(n_625),
    .Y(n_1848));
 AOI22xp5_ASAP7_75t_SL g11275__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[30]),
    .B2(n_625),
    .Y(n_1847));
 AOI22xp5_ASAP7_75t_SL g11276__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]),
    .A2(n_624),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[31]),
    .B2(n_625),
    .Y(n_1846));
 AOI22xp5_ASAP7_75t_SL g11277__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[32]),
    .B2(n_636),
    .Y(n_1845));
 AOI22xp5_ASAP7_75t_SL g11278__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[33]),
    .B2(n_636),
    .Y(n_1844));
 AOI22xp5_ASAP7_75t_SL g11279__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[34]),
    .B2(n_636),
    .Y(n_1843));
 INVx1_ASAP7_75t_SL g1128 (.A(n_13008),
    .Y(n_6030));
 AOI22xp5_ASAP7_75t_SL g11280__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[35]),
    .B2(n_636),
    .Y(n_1842));
 AOI22xp5_ASAP7_75t_SL g11281__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[36]),
    .B2(n_636),
    .Y(n_1841));
 AOI22xp5_ASAP7_75t_SL g11282__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[37]),
    .B2(n_636),
    .Y(n_1840));
 AOI22xp5_ASAP7_75t_SL g11283__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[38]),
    .B2(n_636),
    .Y(n_1839));
 AOI22xp5_ASAP7_75t_SL g11284__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]),
    .A2(n_635),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[39]),
    .B2(n_636),
    .Y(n_1838));
 AOI22xp5_ASAP7_75t_SL g11285__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[40]),
    .B2(n_608),
    .Y(n_1837));
 AOI22xp5_ASAP7_75t_SL g11286__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[41]),
    .B2(n_608),
    .Y(n_1836));
 AOI22xp5_ASAP7_75t_SL g11287__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[42]),
    .B2(n_608),
    .Y(n_1835));
 AOI22xp5_ASAP7_75t_SL g11288__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[43]),
    .B2(n_608),
    .Y(n_1834));
 AOI22xp5_ASAP7_75t_SL g11289__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[44]),
    .B2(n_608),
    .Y(n_1833));
 INVxp67_ASAP7_75t_SL g1129 (.A(n_20653),
    .Y(n_20654));
 AOI22xp5_ASAP7_75t_SL g11290__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[45]),
    .B2(n_608),
    .Y(n_1832));
 AOI22xp5_ASAP7_75t_SL g11291__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[46]),
    .B2(n_608),
    .Y(n_1831));
 AOI22xp5_ASAP7_75t_SL g11292__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]),
    .A2(n_607),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[47]),
    .B2(n_608),
    .Y(n_1830));
 AOI22xp5_ASAP7_75t_SL g11293__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[48]),
    .B2(n_594),
    .Y(n_1829));
 AOI22xp5_ASAP7_75t_SL g11294__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[49]),
    .B2(n_594),
    .Y(n_1828));
 AOI22xp5_ASAP7_75t_SL g11295__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[50]),
    .B2(n_594),
    .Y(n_1827));
 AOI22xp5_ASAP7_75t_SL g11296__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[51]),
    .B2(n_594),
    .Y(n_1826));
 AOI22xp5_ASAP7_75t_SL g11297__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[52]),
    .B2(n_594),
    .Y(n_1825));
 AOI22xp5_ASAP7_75t_SL g11298__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[53]),
    .B2(n_594),
    .Y(n_1824));
 AOI22xp5_ASAP7_75t_SL g11299__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[54]),
    .B2(n_594),
    .Y(n_1823));
 INVx1_ASAP7_75t_SL g113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_43),
    .Y(n_5511));
 XNOR2xp5_ASAP7_75t_SL g1130 (.A(n_6034),
    .B(n_18168),
    .Y(n_6035));
 AOI22xp5_ASAP7_75t_SL g11300__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]),
    .A2(n_593),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[55]),
    .B2(n_594),
    .Y(n_1822));
 AOI22xp5_ASAP7_75t_SL g11301__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[56]),
    .B2(n_606),
    .Y(n_1821));
 AOI22xp5_ASAP7_75t_SL g11302__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[57]),
    .B2(n_606),
    .Y(n_1820));
 AOI22xp5_ASAP7_75t_SL g11303__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[58]),
    .B2(n_606),
    .Y(n_1819));
 AOI22xp5_ASAP7_75t_SL g11304__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[59]),
    .B2(n_606),
    .Y(n_1818));
 AOI22xp5_ASAP7_75t_SL g11305__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[60]),
    .B2(n_606),
    .Y(n_1817));
 AOI22xp5_ASAP7_75t_SL g11306__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[61]),
    .B2(n_606),
    .Y(n_1816));
 AOI22xp5_ASAP7_75t_SL g11307__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[62]),
    .B2(n_606),
    .Y(n_1815));
 AOI22xp5_ASAP7_75t_SL g11308__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]),
    .A2(n_605),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[63]),
    .B2(n_606),
    .Y(n_1814));
 AOI22xp5_ASAP7_75t_SL g11309__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[0]),
    .B2(n_658),
    .Y(n_1813));
 INVxp67_ASAP7_75t_SL g1131 (.A(n_20645),
    .Y(n_20651));
 AOI22xp5_ASAP7_75t_SL g11310__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[1]),
    .B2(n_658),
    .Y(n_1812));
 AOI22xp5_ASAP7_75t_SL g11311__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[2]),
    .B2(n_658),
    .Y(n_1811));
 AOI22xp5_ASAP7_75t_SL g11312__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[3]),
    .B2(n_658),
    .Y(n_1810));
 AOI22xp5_ASAP7_75t_SL g11313__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[4]),
    .B2(n_658),
    .Y(n_1809));
 AOI22xp5_ASAP7_75t_SL g11314__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[5]),
    .B2(n_658),
    .Y(n_1808));
 AOI22xp5_ASAP7_75t_SL g11315__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[6]),
    .B2(n_658),
    .Y(n_1807));
 AOI22xp5_ASAP7_75t_SL g11316__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]),
    .A2(n_657),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[7]),
    .B2(n_658),
    .Y(n_1806));
 AOI22xp5_ASAP7_75t_SL g11317__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[8]),
    .B2(n_596),
    .Y(n_1805));
 AOI22xp5_ASAP7_75t_SL g11318__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[9]),
    .B2(n_596),
    .Y(n_1804));
 AOI22xp5_ASAP7_75t_SL g11319__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[10]),
    .B2(n_596),
    .Y(n_1803));
 NAND3x2_ASAP7_75t_SL g1132 (.B(n_18168),
    .C(n_6024),
    .Y(n_6025),
    .A(n_6022));
 AOI22xp5_ASAP7_75t_SL g11320__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[11]),
    .B2(n_596),
    .Y(n_1802));
 AOI22xp5_ASAP7_75t_SL g11321__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[12]),
    .B2(n_596),
    .Y(n_1801));
 AOI22xp5_ASAP7_75t_SL g11322__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[13]),
    .B2(n_596),
    .Y(n_1800));
 AOI22xp5_ASAP7_75t_SL g11323__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[14]),
    .B2(n_596),
    .Y(n_1799));
 AOI22xp5_ASAP7_75t_SL g11324__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]),
    .A2(n_595),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[15]),
    .B2(n_596),
    .Y(n_1798));
 AOI22xp5_ASAP7_75t_SL g11325__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[16]),
    .B2(n_604),
    .Y(n_1797));
 AOI22xp5_ASAP7_75t_SL g11326__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[17]),
    .B2(n_604),
    .Y(n_1796));
 AOI22xp5_ASAP7_75t_SL g11327__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[18]),
    .B2(n_604),
    .Y(n_1795));
 AOI22xp5_ASAP7_75t_SL g11328__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[19]),
    .B2(n_604),
    .Y(n_1794));
 AOI22xp5_ASAP7_75t_SL g11329__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[20]),
    .B2(n_604),
    .Y(n_1793));
 AND2x2_ASAP7_75t_SL g1133 (.A(n_6022),
    .B(n_12152),
    .Y(n_6031));
 AOI22xp5_ASAP7_75t_SL g11330__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[21]),
    .B2(n_604),
    .Y(n_1792));
 AOI22xp5_ASAP7_75t_SL g11331__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[22]),
    .B2(n_604),
    .Y(n_1791));
 AOI22xp5_ASAP7_75t_SL g11332__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]),
    .A2(n_603),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[23]),
    .B2(n_604),
    .Y(n_1790));
 AOI22xp5_ASAP7_75t_SL g11333__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[24]),
    .B2(n_652),
    .Y(n_1789));
 AOI22xp5_ASAP7_75t_SL g11334__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[25]),
    .B2(n_652),
    .Y(n_1788));
 AOI22xp5_ASAP7_75t_SL g11335__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[26]),
    .B2(n_652),
    .Y(n_1787));
 AOI22xp5_ASAP7_75t_SL g11336__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[27]),
    .B2(n_652),
    .Y(n_1786));
 AOI22xp5_ASAP7_75t_SL g11337__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[28]),
    .B2(n_652),
    .Y(n_1785));
 AOI22xp5_ASAP7_75t_SL g11338__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[29]),
    .B2(n_652),
    .Y(n_1784));
 AOI22xp5_ASAP7_75t_SL g11339__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[30]),
    .B2(n_652),
    .Y(n_1783));
 NAND2xp5_ASAP7_75t_SL g1134 (.A(n_6024),
    .B(n_6019),
    .Y(n_6034));
 AOI22xp5_ASAP7_75t_SL g11340__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]),
    .A2(n_651),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[31]),
    .B2(n_652),
    .Y(n_1782));
 AOI22xp5_ASAP7_75t_SL g11341__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[32]),
    .B2(n_588),
    .Y(n_1781));
 AOI22xp5_ASAP7_75t_SL g11342__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[33]),
    .B2(n_588),
    .Y(n_1780));
 AOI22xp5_ASAP7_75t_SL g11343__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[34]),
    .B2(n_588),
    .Y(n_1779));
 AOI22xp5_ASAP7_75t_SL g11344__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[35]),
    .B2(n_588),
    .Y(n_1778));
 AOI22xp5_ASAP7_75t_SL g11345__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[36]),
    .B2(n_588),
    .Y(n_1777));
 AOI22xp5_ASAP7_75t_SL g11346__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[37]),
    .B2(n_588),
    .Y(n_1776));
 AOI22xp5_ASAP7_75t_SL g11347__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[38]),
    .B2(n_588),
    .Y(n_1775));
 AOI22xp5_ASAP7_75t_SL g11348__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]),
    .A2(n_587),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[39]),
    .B2(n_588),
    .Y(n_1774));
 AOI22xp5_ASAP7_75t_SL g11349__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[40]),
    .B2(n_592),
    .Y(n_1773));
 AOI21xp5_ASAP7_75t_SL g1135 (.A1(n_20638),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_193),
    .B(n_20639),
    .Y(n_20640));
 AOI22xp5_ASAP7_75t_SL g11350__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[41]),
    .B2(n_592),
    .Y(n_1772));
 AOI22xp5_ASAP7_75t_SL g11351__8428 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[42]),
    .B2(n_592),
    .Y(n_1771));
 AOI22xp5_ASAP7_75t_SL g11352__5526 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[43]),
    .B2(n_592),
    .Y(n_1770));
 AOI22xp5_ASAP7_75t_SL g11353__6783 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[44]),
    .B2(n_592),
    .Y(n_1769));
 AOI22xp5_ASAP7_75t_SL g11354__3680 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[45]),
    .B2(n_592),
    .Y(n_1768));
 AOI22xp5_ASAP7_75t_SL g11355__1617 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[46]),
    .B2(n_592),
    .Y(n_1767));
 AOI22xp5_ASAP7_75t_SL g11356__2802 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]),
    .A2(n_591),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[47]),
    .B2(n_592),
    .Y(n_1766));
 AOI22xp5_ASAP7_75t_SL g11357__1705 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[48]),
    .B2(n_590),
    .Y(n_1765));
 AOI22xp5_ASAP7_75t_SL g11358__5122 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[49]),
    .B2(n_590),
    .Y(n_1764));
 AOI22xp5_ASAP7_75t_SL g11359__8246 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[50]),
    .B2(n_590),
    .Y(n_1763));
 INVx2_ASAP7_75t_SL g1136 (.A(n_20758),
    .Y(n_6022));
 AOI22xp5_ASAP7_75t_SL g11360__7098 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[51]),
    .B2(n_590),
    .Y(n_1762));
 AOI22xp5_ASAP7_75t_SL g11361__6131 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[52]),
    .B2(n_590),
    .Y(n_1761));
 AOI22xp5_ASAP7_75t_SL g11362__1881 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[53]),
    .B2(n_590),
    .Y(n_1760));
 AOI22xp5_ASAP7_75t_SL g11363__5115 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[54]),
    .B2(n_590),
    .Y(n_1759));
 AOI22xp5_ASAP7_75t_SL g11364__7482 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]),
    .A2(n_589),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[55]),
    .B2(n_590),
    .Y(n_1758));
 AOI22xp5_ASAP7_75t_SL g11365__4733 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[56]),
    .B2(n_660),
    .Y(n_1757));
 AOI22xp5_ASAP7_75t_SL g11366__6161 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[57]),
    .B2(n_660),
    .Y(n_1756));
 AOI22xp5_ASAP7_75t_SL g11367__9315 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[58]),
    .B2(n_660),
    .Y(n_1755));
 AOI22xp5_ASAP7_75t_SL g11368__9945 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[59]),
    .B2(n_660),
    .Y(n_1754));
 AOI22xp5_ASAP7_75t_SL g11369__2883 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[60]),
    .B2(n_660),
    .Y(n_1753));
 AOI22xp5_ASAP7_75t_SL g11370__2346 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[61]),
    .B2(n_660),
    .Y(n_1752));
 AOI22xp5_ASAP7_75t_SL g11371__1666 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[62]),
    .B2(n_660),
    .Y(n_1751));
 AOI22xp5_ASAP7_75t_SL g11372__7410 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]),
    .A2(n_659),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[63]),
    .B2(n_660),
    .Y(n_1750));
 AOI22xp5_ASAP7_75t_SL g11373__6417 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[0]),
    .B2(n_620),
    .Y(n_1749));
 AOI22xp5_ASAP7_75t_SL g11374__5477 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[1]),
    .B2(n_620),
    .Y(n_1748));
 AOI22xp5_ASAP7_75t_SL g11375__2398 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[2]),
    .B2(n_620),
    .Y(n_1747));
 AOI22xp5_ASAP7_75t_SL g11376__5107 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[3]),
    .B2(n_620),
    .Y(n_1746));
 AOI22xp5_ASAP7_75t_SL g11377__6260 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[4]),
    .B2(n_620),
    .Y(n_1745));
 AOI22xp5_ASAP7_75t_SL g11378__4319 (.A1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]),
    .A2(n_619),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[5]),
    .B2(n_620),
    .Y(n_1744));
 AOI22xp5_ASAP7_75t_SL g11379__8428 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[0]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]),
    .B2(n_827),
    .Y(n_1743));
 AOI22xp5_ASAP7_75t_SL g11380__5526 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[1]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]),
    .B2(n_827),
    .Y(n_1742));
 AOI22xp5_ASAP7_75t_SL g11381__6783 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[2]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]),
    .B2(n_827),
    .Y(n_1741));
 AOI22xp5_ASAP7_75t_SL g11382__3680 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[3]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]),
    .B2(n_827),
    .Y(n_1740));
 AOI22xp5_ASAP7_75t_SL g11383__1617 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[4]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]),
    .B2(n_827),
    .Y(n_1739));
 AOI22xp5_ASAP7_75t_SL g11384__2802 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[5]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]),
    .B2(n_827),
    .Y(n_1738));
 AOI22xp5_ASAP7_75t_SL g11385__1705 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[6]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]),
    .B2(n_827),
    .Y(n_1737));
 AOI22xp5_ASAP7_75t_SL g11386__5122 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[7]),
    .A2(n_826),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]),
    .B2(n_827),
    .Y(n_1736));
 AOI22xp5_ASAP7_75t_SL g11387__8246 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[0]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]),
    .B2(n_830),
    .Y(n_1735));
 AOI22xp5_ASAP7_75t_SL g11388__7098 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[1]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]),
    .B2(n_830),
    .Y(n_1734));
 AOI22xp5_ASAP7_75t_SL g11389__6131 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[2]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]),
    .B2(n_830),
    .Y(n_1733));
 NAND2xp5_ASAP7_75t_SL g1139 (.A(n_11627),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_245),
    .Y(n_6024));
 AOI22xp5_ASAP7_75t_SL g11390__1881 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[3]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]),
    .B2(n_830),
    .Y(n_1732));
 AOI22xp5_ASAP7_75t_SL g11391__5115 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[4]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]),
    .B2(n_830),
    .Y(n_1731));
 AOI22xp5_ASAP7_75t_SL g11392__7482 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[5]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]),
    .B2(n_830),
    .Y(n_1730));
 AOI22xp5_ASAP7_75t_SL g11393__4733 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[6]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]),
    .B2(n_830),
    .Y(n_1729));
 AOI22xp5_ASAP7_75t_SL g11394__6161 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[7]),
    .A2(n_829),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]),
    .B2(n_830),
    .Y(n_1728));
 AOI22xp5_ASAP7_75t_SL g11395__9315 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[0]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]),
    .B2(n_832),
    .Y(n_1727));
 AOI22xp5_ASAP7_75t_SL g11396__9945 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[1]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]),
    .B2(n_832),
    .Y(n_1726));
 AOI22xp5_ASAP7_75t_SL g11397__2883 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[2]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]),
    .B2(n_832),
    .Y(n_1725));
 AOI22xp5_ASAP7_75t_SL g11398__2346 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[3]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]),
    .B2(n_832),
    .Y(n_1724));
 AOI22xp5_ASAP7_75t_SL g11399__1666 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[4]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]),
    .B2(n_832),
    .Y(n_1723));
 INVxp67_ASAP7_75t_SL g114 (.A(n_9991),
    .Y(n_6016));
 INVxp67_ASAP7_75t_SL g1140 (.A(n_6019),
    .Y(n_6032));
 AOI22xp5_ASAP7_75t_SL g11400__7410 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[5]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]),
    .B2(n_832),
    .Y(n_1722));
 AOI22xp5_ASAP7_75t_SL g11401__6417 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[6]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]),
    .B2(n_832),
    .Y(n_1721));
 AOI22xp5_ASAP7_75t_SL g11402__5477 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[7]),
    .A2(n_831),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]),
    .B2(n_832),
    .Y(n_1720));
 AOI22xp5_ASAP7_75t_SL g11403__2398 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[0]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]),
    .B2(n_842),
    .Y(n_1719));
 AOI22xp5_ASAP7_75t_SL g11404__5107 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[1]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]),
    .B2(n_842),
    .Y(n_1718));
 AOI22xp5_ASAP7_75t_SL g11405__6260 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[2]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]),
    .B2(n_842),
    .Y(n_1717));
 AOI22xp5_ASAP7_75t_SL g11406__4319 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[3]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]),
    .B2(n_842),
    .Y(n_1716));
 AOI22xp5_ASAP7_75t_SL g11407__8428 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[4]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]),
    .B2(n_842),
    .Y(n_1715));
 AOI22xp5_ASAP7_75t_SL g11408__5526 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[5]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]),
    .B2(n_842),
    .Y(n_1714));
 AOI22xp5_ASAP7_75t_SL g11409__6783 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[6]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]),
    .B2(n_842),
    .Y(n_1713));
 OR2x2_ASAP7_75t_SL g1141 (.A(n_11627),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_245),
    .Y(n_6019));
 AOI22xp5_ASAP7_75t_SL g11410__3680 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[7]),
    .A2(n_841),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]),
    .B2(n_842),
    .Y(n_1712));
 AOI22xp5_ASAP7_75t_SL g11411__1617 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[0]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]),
    .B2(n_837),
    .Y(n_1711));
 AOI22xp5_ASAP7_75t_SL g11412__2802 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[1]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]),
    .B2(n_837),
    .Y(n_1710));
 AOI22xp5_ASAP7_75t_SL g11413__1705 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[2]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]),
    .B2(n_837),
    .Y(n_1709));
 AOI22xp5_ASAP7_75t_SL g11414__5122 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[3]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]),
    .B2(n_837),
    .Y(n_1708));
 AOI22xp5_ASAP7_75t_SL g11415__8246 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[4]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]),
    .B2(n_837),
    .Y(n_1707));
 AOI22xp5_ASAP7_75t_SL g11416__7098 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[5]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]),
    .B2(n_837),
    .Y(n_1706));
 AOI22xp5_ASAP7_75t_SL g11417__6131 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[6]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]),
    .B2(n_837),
    .Y(n_1705));
 AOI22xp5_ASAP7_75t_SL g11418__1881 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[7]),
    .A2(n_836),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]),
    .B2(n_837),
    .Y(n_1704));
 AOI22xp5_ASAP7_75t_SL g11419__5115 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[0]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]),
    .B2(n_654),
    .Y(n_1703));
 NOR2xp33_ASAP7_75t_SL g1142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_286),
    .B(n_11343),
    .Y(n_20649));
 AOI22xp5_ASAP7_75t_SL g11420__7482 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[1]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]),
    .B2(n_654),
    .Y(n_1702));
 AOI22xp5_ASAP7_75t_SL g11421__4733 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[2]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]),
    .B2(n_654),
    .Y(n_1701));
 AOI22xp5_ASAP7_75t_SL g11422__6161 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[3]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]),
    .B2(n_654),
    .Y(n_1700));
 AOI22xp5_ASAP7_75t_SL g11423__9315 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[4]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]),
    .B2(n_654),
    .Y(n_1699));
 AOI22xp5_ASAP7_75t_SL g11424__9945 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[5]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]),
    .B2(n_654),
    .Y(n_1698));
 AOI22xp5_ASAP7_75t_SL g11425__2883 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[6]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]),
    .B2(n_654),
    .Y(n_1697));
 AOI22xp5_ASAP7_75t_SL g11426__2346 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[7]),
    .A2(n_653),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]),
    .B2(n_654),
    .Y(n_1696));
 AOI22xp5_ASAP7_75t_SL g11427__1666 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[0]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]),
    .B2(n_840),
    .Y(n_1695));
 AOI22xp5_ASAP7_75t_SL g11428__7410 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[1]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]),
    .B2(n_840),
    .Y(n_1694));
 AOI22xp5_ASAP7_75t_SL g11429__6417 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[2]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]),
    .B2(n_840),
    .Y(n_1693));
 NOR2xp33_ASAP7_75t_SL g1143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_250),
    .Y(n_20639));
 AOI22xp5_ASAP7_75t_SL g11430__5477 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[3]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]),
    .B2(n_840),
    .Y(n_1692));
 AOI22xp5_ASAP7_75t_SL g11431__2398 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[4]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]),
    .B2(n_840),
    .Y(n_1691));
 AOI22xp5_ASAP7_75t_SL g11432__5107 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[5]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]),
    .B2(n_840),
    .Y(n_1690));
 AOI22xp5_ASAP7_75t_SL g11433__6260 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[6]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]),
    .B2(n_840),
    .Y(n_1689));
 AOI22xp5_ASAP7_75t_SL g11434__4319 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[7]),
    .A2(n_839),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]),
    .B2(n_840),
    .Y(n_1688));
 AOI22xp5_ASAP7_75t_SL g11435__8428 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[0]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]),
    .B2(n_844),
    .Y(n_1687));
 AOI22xp5_ASAP7_75t_SL g11436__5526 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[1]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]),
    .B2(n_844),
    .Y(n_1686));
 AOI22xp5_ASAP7_75t_SL g11437__6783 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[2]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]),
    .B2(n_844),
    .Y(n_1685));
 AOI22xp5_ASAP7_75t_SL g11438__3680 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[3]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]),
    .B2(n_844),
    .Y(n_1684));
 AOI22xp5_ASAP7_75t_SL g11439__1617 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[4]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]),
    .B2(n_844),
    .Y(n_1683));
 INVxp67_ASAP7_75t_SL g1144 (.A(n_20765),
    .Y(n_20642));
 AOI22xp5_ASAP7_75t_SL g11440__2802 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[5]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]),
    .B2(n_844),
    .Y(n_1682));
 AOI22xp5_ASAP7_75t_SL g11441__1705 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[0]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[0]),
    .B2(n_846),
    .Y(n_1681));
 AOI22xp5_ASAP7_75t_SL g11442__5122 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[6]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]),
    .B2(n_844),
    .Y(n_1680));
 AOI22xp5_ASAP7_75t_SL g11443__8246 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[7]),
    .A2(n_843),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]),
    .B2(n_844),
    .Y(n_1679));
 AOI22xp5_ASAP7_75t_SL g11444__7098 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[1]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[1]),
    .B2(n_846),
    .Y(n_1678));
 AOI22xp5_ASAP7_75t_SL g11445__6131 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[2]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[2]),
    .B2(n_846),
    .Y(n_1677));
 AOI22xp5_ASAP7_75t_SL g11446__1881 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[3]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[3]),
    .B2(n_846),
    .Y(n_1676));
 AOI22xp5_ASAP7_75t_SL g11447__5115 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[4]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[4]),
    .B2(n_846),
    .Y(n_1675));
 AOI22xp5_ASAP7_75t_SL g11448__7482 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[6]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[6]),
    .B2(n_846),
    .Y(n_1674));
 AOI22xp5_ASAP7_75t_SL g11449__4733 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[7]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[7]),
    .B2(n_846),
    .Y(n_1673));
 INVxp67_ASAP7_75t_SL g1145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_208),
    .Y(n_20641));
 AOI22xp5_ASAP7_75t_SL g11450__6161 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[5]),
    .A2(n_845),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[5]),
    .B2(n_846),
    .Y(n_1672));
 AOI22xp5_ASAP7_75t_SL g11451 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[0]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[8]),
    .B2(n_851),
    .Y(n_1671));
 AOI22xp5_ASAP7_75t_SL g11452 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[1]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[9]),
    .B2(n_851),
    .Y(n_1670));
 AOI22xp5_ASAP7_75t_SL g11453 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[2]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[10]),
    .B2(n_851),
    .Y(n_1669));
 AOI22xp5_ASAP7_75t_SL g11454 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[4]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[12]),
    .B2(n_851),
    .Y(n_1668));
 AOI22xp5_ASAP7_75t_SL g11455 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[5]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[13]),
    .B2(n_851),
    .Y(n_1667));
 AOI22xp5_ASAP7_75t_SL g11456 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[6]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[14]),
    .B2(n_851),
    .Y(n_1666));
 AOI22xp5_ASAP7_75t_SL g11457 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[7]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[15]),
    .B2(n_851),
    .Y(n_1665));
 AOI22xp5_ASAP7_75t_SL g11458 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[0]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[16]),
    .B2(n_853),
    .Y(n_1664));
 AOI22xp5_ASAP7_75t_SL g11459 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[3]),
    .A2(n_850),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[11]),
    .B2(n_851),
    .Y(n_1663));
 AOI22xp5_ASAP7_75t_SL g11460 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[2]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[18]),
    .B2(n_853),
    .Y(n_1662));
 AOI22xp5_ASAP7_75t_SL g11461 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[3]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[19]),
    .B2(n_853),
    .Y(n_1661));
 AOI22xp5_ASAP7_75t_SL g11462 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[1]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[17]),
    .B2(n_853),
    .Y(n_1660));
 AOI22xp5_ASAP7_75t_SL g11463 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[4]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[20]),
    .B2(n_853),
    .Y(n_1659));
 AOI22xp5_ASAP7_75t_SL g11464 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[5]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[21]),
    .B2(n_853),
    .Y(n_1658));
 AOI22xp5_ASAP7_75t_SL g11465 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[6]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[22]),
    .B2(n_853),
    .Y(n_1657));
 AOI22xp5_ASAP7_75t_SL g11466 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[7]),
    .A2(n_852),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[23]),
    .B2(n_853),
    .Y(n_1656));
 AOI22xp5_ASAP7_75t_SL g11467 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[0]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[24]),
    .B2(n_602),
    .Y(n_1655));
 AOI22xp5_ASAP7_75t_SL g11468 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[1]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[25]),
    .B2(n_602),
    .Y(n_1654));
 AOI22xp5_ASAP7_75t_SL g11469 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[2]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[26]),
    .B2(n_602),
    .Y(n_1653));
 HB1xp67_ASAP7_75t_SL g1147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_250),
    .Y(n_20638));
 AOI22xp5_ASAP7_75t_SL g11470 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[3]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[27]),
    .B2(n_602),
    .Y(n_1652));
 AOI22xp5_ASAP7_75t_SL g11471 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[4]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[28]),
    .B2(n_602),
    .Y(n_1651));
 AOI22xp5_ASAP7_75t_SL g11472 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[5]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[29]),
    .B2(n_602),
    .Y(n_1650));
 AOI22xp5_ASAP7_75t_SL g11473 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[6]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[30]),
    .B2(n_602),
    .Y(n_1649));
 AOI22xp5_ASAP7_75t_SL g11474 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[7]),
    .A2(n_601),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[31]),
    .B2(n_602),
    .Y(n_1648));
 AOI22xp5_ASAP7_75t_SL g11475 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[0]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[32]),
    .B2(n_618),
    .Y(n_1647));
 AOI22xp5_ASAP7_75t_SL g11476 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[1]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[33]),
    .B2(n_618),
    .Y(n_1646));
 AOI22xp5_ASAP7_75t_SL g11477 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[2]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[34]),
    .B2(n_618),
    .Y(n_1645));
 AOI22xp5_ASAP7_75t_SL g11478 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[3]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[35]),
    .B2(n_618),
    .Y(n_1644));
 AOI22xp5_ASAP7_75t_SL g11479 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[4]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[36]),
    .B2(n_618),
    .Y(n_1643));
 AOI22xp5_ASAP7_75t_SL g11480 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[5]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[37]),
    .B2(n_618),
    .Y(n_1642));
 AOI22xp5_ASAP7_75t_SL g11481 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[6]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[38]),
    .B2(n_618),
    .Y(n_1641));
 AOI22xp5_ASAP7_75t_SL g11482 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[7]),
    .A2(n_617),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[39]),
    .B2(n_618),
    .Y(n_1640));
 AOI22xp5_ASAP7_75t_SL g11483 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[0]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[40]),
    .B2(n_848),
    .Y(n_1639));
 AOI22xp5_ASAP7_75t_SL g11484 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[1]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[41]),
    .B2(n_848),
    .Y(n_1638));
 AOI22xp5_ASAP7_75t_SL g11485 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[2]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[42]),
    .B2(n_848),
    .Y(n_1637));
 AOI22xp5_ASAP7_75t_SL g11486 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[4]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[44]),
    .B2(n_848),
    .Y(n_1636));
 AOI22xp5_ASAP7_75t_SL g11487 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[3]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[43]),
    .B2(n_848),
    .Y(n_1635));
 AOI22xp5_ASAP7_75t_SL g11488 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[5]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[45]),
    .B2(n_848),
    .Y(n_1634));
 AOI22xp5_ASAP7_75t_SL g11489 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[6]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[46]),
    .B2(n_848),
    .Y(n_1633));
 AOI22xp5_ASAP7_75t_SL g11490 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[7]),
    .A2(n_847),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[47]),
    .B2(n_848),
    .Y(n_1632));
 AOI22xp5_ASAP7_75t_SL g11491 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[0]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[48]),
    .B2(n_656),
    .Y(n_1631));
 AOI22xp5_ASAP7_75t_SL g11492 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[2]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[50]),
    .B2(n_656),
    .Y(n_1630));
 AOI22xp5_ASAP7_75t_SL g11493 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[1]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[49]),
    .B2(n_656),
    .Y(n_1629));
 AOI22xp5_ASAP7_75t_SL g11494 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[3]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[51]),
    .B2(n_656),
    .Y(n_1628));
 AOI22xp5_ASAP7_75t_SL g11495 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[4]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[52]),
    .B2(n_656),
    .Y(n_1627));
 AOI22xp5_ASAP7_75t_SL g11496 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[5]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[53]),
    .B2(n_656),
    .Y(n_1626));
 AOI22xp5_ASAP7_75t_SL g11497 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[6]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[54]),
    .B2(n_656),
    .Y(n_1625));
 AOI22xp5_ASAP7_75t_SL g11498 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[7]),
    .A2(n_655),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[55]),
    .B2(n_656),
    .Y(n_1624));
 AOI22xp5_ASAP7_75t_SL g11499 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[0]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[56]),
    .B2(n_835),
    .Y(n_1623));
 AND2x2_ASAP7_75t_SL g115 (.A(n_2180),
    .B(n_8481),
    .Y(n_8482));
 AOI22xp5_ASAP7_75t_SL g11500 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[1]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[57]),
    .B2(n_835),
    .Y(n_1622));
 AOI22xp5_ASAP7_75t_SL g11501 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[2]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[58]),
    .B2(n_835),
    .Y(n_1621));
 AOI22xp5_ASAP7_75t_SL g11502 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[3]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[59]),
    .B2(n_835),
    .Y(n_1620));
 AOI22xp5_ASAP7_75t_SL g11503 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[4]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[60]),
    .B2(n_835),
    .Y(n_1619));
 AOI22xp5_ASAP7_75t_SL g11504 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[5]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[61]),
    .B2(n_835),
    .Y(n_1618));
 AOI22xp5_ASAP7_75t_SL g11505 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[6]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[62]),
    .B2(n_835),
    .Y(n_1617));
 AOI22xp5_ASAP7_75t_SL g11506 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[7]),
    .A2(n_834),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[63]),
    .B2(n_835),
    .Y(n_1616));
 AOI22xp5_ASAP7_75t_SL g11507 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .B1(sc2mac_wt_mask[0]),
    .B2(n_585),
    .Y(n_1615));
 AOI22xp5_ASAP7_75t_SL g11508 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .B1(sc2mac_wt_mask[1]),
    .B2(n_585),
    .Y(n_1614));
 AOI22xp5_ASAP7_75t_SL g11509 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .B1(sc2mac_wt_mask[2]),
    .B2(n_585),
    .Y(n_1613));
 AOI22xp5_ASAP7_75t_SL g11510 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .B1(sc2mac_wt_mask[3]),
    .B2(n_585),
    .Y(n_1612));
 AOI22xp5_ASAP7_75t_SL g11511 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .B1(sc2mac_wt_mask[4]),
    .B2(n_585),
    .Y(n_1611));
 AOI22xp5_ASAP7_75t_SL g11512 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .B1(sc2mac_wt_mask[5]),
    .B2(n_585),
    .Y(n_1610));
 AOI22xp5_ASAP7_75t_SL g11513 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .B1(sc2mac_wt_mask[6]),
    .B2(n_585),
    .Y(n_1609));
 AOI22xp5_ASAP7_75t_SL g11514 (.A1(n_586),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .B1(sc2mac_wt_mask[7]),
    .B2(n_585),
    .Y(n_1608));
 AOI22xp5_ASAP7_75t_SL g11515 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .B1(sc2mac_dat_mask[0]),
    .B2(n_583),
    .Y(n_1607));
 AOI22xp5_ASAP7_75t_SL g11516 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .B1(sc2mac_dat_mask[1]),
    .B2(n_583),
    .Y(n_1606));
 AOI22xp5_ASAP7_75t_SL g11517 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .B1(sc2mac_dat_mask[2]),
    .B2(n_583),
    .Y(n_1605));
 AOI22xp5_ASAP7_75t_SL g11518 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .B1(sc2mac_dat_mask[3]),
    .B2(n_583),
    .Y(n_1604));
 AOI22xp5_ASAP7_75t_SL g11519 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .B1(sc2mac_dat_mask[4]),
    .B2(n_583),
    .Y(n_1603));
 AOI22xp5_ASAP7_75t_SL g11520 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .B1(sc2mac_dat_mask[5]),
    .B2(n_583),
    .Y(n_1602));
 AOI22xp5_ASAP7_75t_SL g11521 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .B1(sc2mac_dat_mask[6]),
    .B2(n_583),
    .Y(n_1601));
 AOI22xp5_ASAP7_75t_SL g11522 (.A1(n_584),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .B1(sc2mac_dat_mask[7]),
    .B2(n_583),
    .Y(n_1600));
 AOI21xp5_ASAP7_75t_SL g11523 (.A1(n_854),
    .A2(u_NV_NVDLA_cmac_u_core_wt3_actv_pvld[7]),
    .B(n_581),
    .Y(n_1599));
 INVx1_ASAP7_75t_SL g116 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_243),
    .Y(n_20752));
 AOI22xp5_ASAP7_75t_SL g11654 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[0]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1598));
 AOI22xp5_ASAP7_75t_SL g11655 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[1]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[1]),
    .Y(n_1597));
 AOI22xp5_ASAP7_75t_SL g11656 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[4]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[4]),
    .Y(n_1596));
 AOI22xp5_ASAP7_75t_SL g11657 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[3]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[3]),
    .Y(n_1595));
 AOI22xp5_ASAP7_75t_SL g11658 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[3]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[3]),
    .Y(n_1594));
 AOI22xp5_ASAP7_75t_SL g11659 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[7]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[7]),
    .Y(n_1593));
 AOI22xp5_ASAP7_75t_SL g11660 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[2]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[2]),
    .Y(n_1592));
 AOI22xp5_ASAP7_75t_SL g11661 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[4]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[4]),
    .Y(n_1591));
 AOI22xp5_ASAP7_75t_SL g11662 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[3]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[3]),
    .Y(n_1590));
 AOI22xp5_ASAP7_75t_SL g11663 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[4]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[4]),
    .Y(n_1589));
 AOI22xp5_ASAP7_75t_SL g11664 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[7]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[7]),
    .Y(n_1588));
 AOI22xp5_ASAP7_75t_SL g11665 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[0]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[0]),
    .Y(n_1587));
 AOI22xp5_ASAP7_75t_SL g11666 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[1]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[1]),
    .Y(n_1586));
 AOI22xp5_ASAP7_75t_SL g11667 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[2]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[2]),
    .Y(n_1585));
 AOI22xp5_ASAP7_75t_SL g11668 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[3]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[3]),
    .Y(n_1584));
 AOI22xp5_ASAP7_75t_SL g11669 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[5]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[5]),
    .Y(n_1583));
 AOI22xp5_ASAP7_75t_SL g11670 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[6]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[6]),
    .Y(n_1582));
 AOI22xp5_ASAP7_75t_SL g11671 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[7]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[7]),
    .Y(n_1581));
 AOI22xp5_ASAP7_75t_SL g11672 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[4]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[4]),
    .Y(n_1580));
 AOI22xp5_ASAP7_75t_SL g11673 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[0]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[0]),
    .Y(n_1579));
 AOI22xp5_ASAP7_75t_SL g11674 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[1]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[1]),
    .Y(n_1578));
 AOI22xp5_ASAP7_75t_SL g11675 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[2]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[2]),
    .Y(n_1577));
 AOI22xp5_ASAP7_75t_SL g11676 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[3]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[3]),
    .Y(n_1576));
 AOI22xp5_ASAP7_75t_SL g11677 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[4]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[4]),
    .Y(n_1575));
 AOI22xp5_ASAP7_75t_SL g11678 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[5]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[5]),
    .Y(n_1574));
 AOI22xp5_ASAP7_75t_SL g11679 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[6]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[6]),
    .Y(n_1573));
 AOI22xp5_ASAP7_75t_SL g11680 (.A1(n_35),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[7]),
    .B1(sc2mac_dat_mask[1]),
    .B2(sc2mac_dat_data1[7]),
    .Y(n_1572));
 AOI22xp5_ASAP7_75t_SL g11681 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[0]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[0]),
    .Y(n_1571));
 AOI22xp5_ASAP7_75t_SL g11682 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[0]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[0]),
    .Y(n_1570));
 AOI22xp5_ASAP7_75t_SL g11683 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[1]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[1]),
    .Y(n_1569));
 AOI22xp5_ASAP7_75t_SL g11684 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[2]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[2]),
    .Y(n_1568));
 AOI22xp5_ASAP7_75t_SL g11685 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[3]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[3]),
    .Y(n_1567));
 AOI22xp5_ASAP7_75t_SL g11686 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[4]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[4]),
    .Y(n_1566));
 AOI22xp5_ASAP7_75t_SL g11687 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[5]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[5]),
    .Y(n_1565));
 AOI22xp5_ASAP7_75t_SL g11688 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[6]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[6]),
    .Y(n_1564));
 AOI22xp5_ASAP7_75t_SL g11689 (.A1(n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[7]),
    .B1(sc2mac_dat_mask[2]),
    .B2(sc2mac_dat_data2[7]),
    .Y(n_1563));
 AOI22xp5_ASAP7_75t_SL g11690 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[0]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[0]),
    .Y(n_1562));
 AOI22xp5_ASAP7_75t_SL g11691 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[1]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[1]),
    .Y(n_1561));
 AOI22xp5_ASAP7_75t_SL g11692 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[2]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[2]),
    .Y(n_1560));
 AOI22xp5_ASAP7_75t_SL g11693 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[3]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[3]),
    .Y(n_1559));
 AOI22xp5_ASAP7_75t_SL g11694 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[4]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[4]),
    .Y(n_1558));
 AOI22xp5_ASAP7_75t_SL g11695 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[5]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[5]),
    .Y(n_1557));
 AOI22xp5_ASAP7_75t_SL g11696 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[6]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[6]),
    .Y(n_1556));
 AOI22xp5_ASAP7_75t_SL g11697 (.A1(n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[7]),
    .B1(sc2mac_dat_mask[3]),
    .B2(sc2mac_dat_data3[7]),
    .Y(n_1555));
 AOI22xp5_ASAP7_75t_SL g11698 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[0]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[0]),
    .Y(n_1554));
 AOI22xp5_ASAP7_75t_SL g11699 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[1]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[1]),
    .Y(n_1553));
 AOI22xp5_ASAP7_75t_SL g117 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_156),
    .B1(n_5549),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_140),
    .Y(n_9089));
 AOI22xp5_ASAP7_75t_SL g11700 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[2]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[2]),
    .Y(n_1552));
 AOI22xp5_ASAP7_75t_SL g11701 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[4]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[4]),
    .Y(n_1551));
 AOI22xp5_ASAP7_75t_SL g11702 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[5]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[5]),
    .Y(n_1550));
 AOI22xp5_ASAP7_75t_SL g11703 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[5]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[5]),
    .Y(n_1549));
 AOI22xp5_ASAP7_75t_SL g11704 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[6]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[6]),
    .Y(n_1548));
 AOI22xp5_ASAP7_75t_SL g11705 (.A1(n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[7]),
    .B1(sc2mac_dat_mask[4]),
    .B2(sc2mac_dat_data4[7]),
    .Y(n_1547));
 AOI22xp5_ASAP7_75t_SL g11706 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[4]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[4]),
    .Y(n_1546));
 AOI22xp5_ASAP7_75t_SL g11707 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[0]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[0]),
    .Y(n_1545));
 AOI22xp5_ASAP7_75t_SL g11708 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[1]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[1]),
    .Y(n_1544));
 AOI22xp5_ASAP7_75t_SL g11709 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[2]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[2]),
    .Y(n_1543));
 AOI22xp5_ASAP7_75t_SL g11710 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[3]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[3]),
    .Y(n_1542));
 AOI22xp5_ASAP7_75t_SL g11711 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[5]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[5]),
    .Y(n_1541));
 AOI22xp5_ASAP7_75t_SL g11712 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[6]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[6]),
    .Y(n_1540));
 AOI22xp5_ASAP7_75t_SL g11713 (.A1(n_38),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[7]),
    .B1(sc2mac_dat_mask[5]),
    .B2(sc2mac_dat_data5[7]),
    .Y(n_1539));
 AOI22xp5_ASAP7_75t_SL g11714 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[1]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[1]),
    .Y(n_1538));
 AOI22xp5_ASAP7_75t_SL g11715 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[0]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[0]),
    .Y(n_1537));
 AOI22xp5_ASAP7_75t_SL g11716 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[1]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[1]),
    .Y(n_1536));
 AOI22xp5_ASAP7_75t_SL g11717 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[2]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[2]),
    .Y(n_1535));
 AOI22xp5_ASAP7_75t_SL g11718 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[3]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[3]),
    .Y(n_1534));
 AOI22xp5_ASAP7_75t_SL g11719 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[4]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[4]),
    .Y(n_1533));
 AOI22xp5_ASAP7_75t_SL g11720 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[5]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[5]),
    .Y(n_1532));
 AOI22xp5_ASAP7_75t_SL g11721 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[6]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[6]),
    .Y(n_1531));
 AOI22xp5_ASAP7_75t_SL g11722 (.A1(n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[7]),
    .B1(sc2mac_dat_mask[6]),
    .B2(sc2mac_dat_data6[7]),
    .Y(n_1530));
 AOI22xp5_ASAP7_75t_SL g11723 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[0]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[0]),
    .Y(n_1529));
 AOI22xp5_ASAP7_75t_SL g11724 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[1]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[1]),
    .Y(n_1528));
 AOI22xp5_ASAP7_75t_SL g11725 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[2]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[2]),
    .Y(n_1527));
 AOI22xp5_ASAP7_75t_SL g11726 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[3]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[3]),
    .Y(n_1526));
 AOI22xp5_ASAP7_75t_SL g11727 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[5]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[5]),
    .Y(n_1525));
 AOI22xp5_ASAP7_75t_SL g11728 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[6]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[6]),
    .Y(n_1524));
 AOI22xp5_ASAP7_75t_SL g11729 (.A1(n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[7]),
    .B1(sc2mac_dat_mask[7]),
    .B2(sc2mac_dat_data7[7]),
    .Y(n_1523));
 AOI22xp5_ASAP7_75t_SL g11730 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[0]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[0]),
    .Y(n_1522));
 AOI22xp5_ASAP7_75t_SL g11731 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[2]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[2]),
    .Y(n_1521));
 AOI22xp5_ASAP7_75t_SL g11732 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[3]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[3]),
    .Y(n_1520));
 AOI22xp5_ASAP7_75t_SL g11733 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[4]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[4]),
    .Y(n_1519));
 AOI22xp5_ASAP7_75t_SL g11734 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[5]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[5]),
    .Y(n_1518));
 AOI22xp5_ASAP7_75t_SL g11735 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[6]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[6]),
    .Y(n_1517));
 AOI22xp5_ASAP7_75t_SL g11736 (.A1(n_36),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[7]),
    .B1(sc2mac_wt_mask[0]),
    .B2(sc2mac_wt_data0[7]),
    .Y(n_1516));
 AOI22xp5_ASAP7_75t_SL g11737 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[4]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[4]),
    .Y(n_1515));
 AOI22xp5_ASAP7_75t_SL g11738 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[0]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[0]),
    .Y(n_1514));
 AOI22xp5_ASAP7_75t_SL g11739 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[1]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[1]),
    .Y(n_1513));
 AOI22xp5_ASAP7_75t_SL g11740 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[2]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[2]),
    .Y(n_1512));
 AOI22xp5_ASAP7_75t_SL g11741 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[4]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[4]),
    .Y(n_1511));
 AOI22xp5_ASAP7_75t_SL g11742 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[5]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[5]),
    .Y(n_1510));
 AOI22xp5_ASAP7_75t_SL g11743 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[6]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[6]),
    .Y(n_1509));
 AOI22xp5_ASAP7_75t_SL g11744 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[7]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[7]),
    .Y(n_1508));
 AOI22xp5_ASAP7_75t_SL g11745 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[2]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[2]),
    .Y(n_1507));
 AOI22xp5_ASAP7_75t_SL g11746 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[1]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[1]),
    .Y(n_1506));
 AOI22xp5_ASAP7_75t_SL g11747 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[0]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[0]),
    .Y(n_1505));
 AOI22xp5_ASAP7_75t_SL g11748 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[1]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[1]),
    .Y(n_1504));
 AOI22xp5_ASAP7_75t_SL g11749 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[2]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[2]),
    .Y(n_1503));
 AOI22xp5_ASAP7_75t_SL g11750 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[3]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[3]),
    .Y(n_1502));
 AOI22xp5_ASAP7_75t_SL g11751 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[4]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[4]),
    .Y(n_1501));
 AOI22xp5_ASAP7_75t_SL g11752 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[5]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[5]),
    .Y(n_1500));
 AOI22xp5_ASAP7_75t_SL g11753 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[6]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[6]),
    .Y(n_1499));
 AOI22xp5_ASAP7_75t_SL g11754 (.A1(n_30),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[7]),
    .B1(sc2mac_wt_mask[2]),
    .B2(sc2mac_wt_data2[7]),
    .Y(n_1498));
 AOI22xp5_ASAP7_75t_SL g11755 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[0]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[0]),
    .Y(n_1497));
 AOI22xp5_ASAP7_75t_SL g11756 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[1]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[1]),
    .Y(n_1496));
 AOI22xp5_ASAP7_75t_SL g11757 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[2]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[2]),
    .Y(n_1495));
 AOI22xp5_ASAP7_75t_SL g11758 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[3]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[3]),
    .Y(n_1494));
 AOI22xp5_ASAP7_75t_SL g11759 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[4]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[4]),
    .Y(n_1493));
 AOI22xp5_ASAP7_75t_SL g11760 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[5]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[5]),
    .Y(n_1492));
 AOI22xp5_ASAP7_75t_SL g11761 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[6]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[6]),
    .Y(n_1491));
 AOI22xp5_ASAP7_75t_SL g11762 (.A1(n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[7]),
    .B1(sc2mac_wt_mask[3]),
    .B2(sc2mac_wt_data3[7]),
    .Y(n_1490));
 AOI22xp5_ASAP7_75t_SL g11763 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[0]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[0]),
    .Y(n_1489));
 AOI22xp5_ASAP7_75t_SL g11764 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[3]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[3]),
    .Y(n_1488));
 AOI22xp5_ASAP7_75t_SL g11765 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[5]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[5]),
    .Y(n_1487));
 AOI22xp5_ASAP7_75t_SL g11766 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[6]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[6]),
    .Y(n_1486));
 AOI22xp5_ASAP7_75t_SL g11767 (.A1(n_34),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[7]),
    .B1(sc2mac_wt_mask[4]),
    .B2(sc2mac_wt_data4[7]),
    .Y(n_1485));
 AOI22xp5_ASAP7_75t_SL g11768 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[0]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[0]),
    .Y(n_1484));
 AOI22xp5_ASAP7_75t_SL g11769 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[2]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[2]),
    .Y(n_1483));
 AOI22xp5_ASAP7_75t_SL g11770 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[3]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[3]),
    .Y(n_1482));
 AOI22xp5_ASAP7_75t_SL g11771 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[6]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[6]),
    .Y(n_1481));
 AOI22xp5_ASAP7_75t_SL g11772 (.A1(n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[7]),
    .B1(sc2mac_wt_mask[5]),
    .B2(sc2mac_wt_data5[7]),
    .Y(n_1480));
 AOI22xp5_ASAP7_75t_SL g11773 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[1]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[1]),
    .Y(n_1479));
 AOI22xp5_ASAP7_75t_SL g11774 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[2]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[2]),
    .Y(n_1478));
 AOI22xp5_ASAP7_75t_SL g11775 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[5]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[5]),
    .Y(n_1477));
 AOI22xp5_ASAP7_75t_SL g11776 (.A1(n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[6]),
    .B1(sc2mac_wt_mask[6]),
    .B2(sc2mac_wt_data6[6]),
    .Y(n_1476));
 AOI22xp5_ASAP7_75t_SL g11777 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[0]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[0]),
    .Y(n_1475));
 AOI22xp5_ASAP7_75t_SL g11778 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[1]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[1]),
    .Y(n_1474));
 AOI22xp5_ASAP7_75t_SL g11779 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[5]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[5]),
    .Y(n_1473));
 AOI22xp5_ASAP7_75t_SL g11780 (.A1(n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[6]),
    .B1(sc2mac_wt_mask[7]),
    .B2(sc2mac_wt_data7[6]),
    .Y(n_1472));
 AOI22xp5_ASAP7_75t_SL g11781 (.A1(n_31),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[4]),
    .B1(sc2mac_dat_mask[0]),
    .B2(sc2mac_dat_data0[4]),
    .Y(n_1471));
 AOI22xp5_ASAP7_75t_SL g11782 (.A1(n_33),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[3]),
    .B1(sc2mac_wt_mask[1]),
    .B2(sc2mac_wt_data1[3]),
    .Y(n_1470));
 AOI22xp5_ASAP7_75t_SL g11783 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[1]),
    .Y(n_1469));
 AOI22xp5_ASAP7_75t_SL g11784 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[2]),
    .Y(n_1468));
 AOI22xp5_ASAP7_75t_SL g11785 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[3]),
    .Y(n_1467));
 AOI22xp5_ASAP7_75t_SL g11786 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[4]),
    .Y(n_1466));
 AOI22xp5_ASAP7_75t_SL g11787 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[5]),
    .Y(n_1465));
 AOI22xp5_ASAP7_75t_SL g11788 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[6]),
    .Y(n_1464));
 AOI22xp5_ASAP7_75t_SL g11789 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[7]),
    .Y(n_1463));
 AOI22xp5_ASAP7_75t_SL g11790 (.A1(mac2accu_pd[0]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[0]),
    .Y(n_1462));
 AOI22xp5_ASAP7_75t_SL g11791 (.A1(mac2accu_pd[1]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[1]),
    .Y(n_1461));
 AOI22xp5_ASAP7_75t_SL g11792 (.A1(mac2accu_pd[2]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[2]),
    .Y(n_1460));
 AOI22xp5_ASAP7_75t_SL g11793 (.A1(mac2accu_pd[3]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[3]),
    .Y(n_1459));
 AOI22xp5_ASAP7_75t_SL g11794 (.A1(mac2accu_pd[4]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[4]),
    .Y(n_1458));
 AOI22xp5_ASAP7_75t_SL g11795 (.A1(mac2accu_pd[5]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[5]),
    .Y(n_1457));
 AOI22xp5_ASAP7_75t_SL g11796 (.A1(mac2accu_pd[6]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[6]),
    .Y(n_1456));
 AOI22xp5_ASAP7_75t_SL g11797 (.A1(mac2accu_pd[7]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[7]),
    .Y(n_1455));
 AOI22xp5_ASAP7_75t_SL g11798 (.A1(mac2accu_pd[8]),
    .A2(n_29),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[8]),
    .Y(n_1454));
 AOI22xp5_ASAP7_75t_SL g11799 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[6]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1453));
 OAI221xp5_ASAP7_75t_SL g118 (.A1(n_16530),
    .A2(n_16532),
    .B1(n_16534),
    .B2(n_16071),
    .C(n_16535),
    .Y(n_16536));
 AOI22xp5_ASAP7_75t_SL g11800 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[5]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1452));
 AOI22xp5_ASAP7_75t_SL g11801 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[7]),
    .Y(n_1451));
 AOI22xp5_ASAP7_75t_SL g11802 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[8]),
    .Y(n_1450));
 AOI22xp5_ASAP7_75t_SL g11803 (.A1(n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[0]),
    .Y(n_1449));
 AOI22xp5_ASAP7_75t_SL g11804 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[7]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1448));
 AOI22xp5_ASAP7_75t_SL g11805 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[6]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1447));
 AOI22xp5_ASAP7_75t_SL g11806 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[6]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1446));
 AOI22xp5_ASAP7_75t_SL g11807 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[1]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1445));
 AOI22xp5_ASAP7_75t_SL g11808 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[4]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1444));
 AOI22xp5_ASAP7_75t_SL g11809 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[2]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1443));
 AOI22xp5_ASAP7_75t_SL g11810 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[6]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1442));
 AOI22xp5_ASAP7_75t_SL g11811 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[3]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1441));
 AOI22xp5_ASAP7_75t_SL g11812 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[0]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1440));
 AOI22xp5_ASAP7_75t_SL g11813 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[0]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1439));
 AOI22xp5_ASAP7_75t_SL g11814 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[1]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1438));
 AOI22xp5_ASAP7_75t_SL g11815 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[2]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1437));
 AOI22xp5_ASAP7_75t_SL g11816 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[4]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1436));
 AOI22xp5_ASAP7_75t_SL g11817 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[5]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1435));
 AOI22xp5_ASAP7_75t_SL g11818 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[6]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1434));
 AOI22xp5_ASAP7_75t_SL g11819 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[7]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1433));
 AOI22xp5_ASAP7_75t_SL g11820 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[0]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1432));
 AOI22xp5_ASAP7_75t_SL g11821 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[5]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1431));
 AOI22xp5_ASAP7_75t_SL g11822 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[1]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1430));
 AOI22xp5_ASAP7_75t_SL g11823 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[2]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1429));
 AOI22xp5_ASAP7_75t_SL g11824 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[3]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1428));
 AOI22xp5_ASAP7_75t_SL g11825 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[4]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1427));
 AOI22xp5_ASAP7_75t_SL g11826 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[7]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1426));
 AOI22xp5_ASAP7_75t_SL g11827 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[5]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1425));
 AOI22xp5_ASAP7_75t_SL g11828 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[6]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1424));
 AOI22xp5_ASAP7_75t_SL g11829 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data1[7]),
    .A2(n_324),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_1423));
 AOI22xp5_ASAP7_75t_SL g11830 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[6]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1422));
 AOI22xp5_ASAP7_75t_SL g11831 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[0]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1421));
 AOI22xp5_ASAP7_75t_SL g11832 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[1]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1420));
 AOI22xp5_ASAP7_75t_SL g11833 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[2]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1419));
 AOI22xp5_ASAP7_75t_SL g11834 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[3]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1418));
 AOI22xp5_ASAP7_75t_SL g11835 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[4]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1417));
 AOI22xp5_ASAP7_75t_SL g11836 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[5]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1416));
 AOI22xp5_ASAP7_75t_SL g11837 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[4]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1415));
 AOI22xp5_ASAP7_75t_SL g11838 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data2[7]),
    .A2(n_328),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_1414));
 AOI22xp5_ASAP7_75t_SL g11839 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[1]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1413));
 AOI22xp5_ASAP7_75t_SL g11841 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[1]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1411));
 AOI22xp5_ASAP7_75t_SL g11842 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[0]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1410));
 AOI22xp5_ASAP7_75t_SL g11843 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[2]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1409));
 AOI22xp5_ASAP7_75t_SL g11844 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[3]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1408));
 AOI22xp5_ASAP7_75t_SL g11845 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[4]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1407));
 AOI22xp5_ASAP7_75t_SL g11846 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[5]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1406));
 AOI22xp5_ASAP7_75t_SL g11847 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[6]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1405));
 AOI22xp5_ASAP7_75t_SL g11848 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data3[7]),
    .A2(n_322),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_1404));
 AOI22xp5_ASAP7_75t_SL g11849 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[0]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1403));
 AOI22xp5_ASAP7_75t_SL g11850 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[0]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1402));
 AOI22xp5_ASAP7_75t_SL g11851 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[1]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1401));
 AOI22xp5_ASAP7_75t_SL g11852 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[2]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1400));
 AOI22xp5_ASAP7_75t_SL g11853 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[3]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1399));
 AOI22xp5_ASAP7_75t_SL g11854 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[4]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1398));
 AOI22xp5_ASAP7_75t_SL g11855 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[5]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1397));
 AOI22xp5_ASAP7_75t_SL g11856 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[6]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1396));
 AOI22xp5_ASAP7_75t_SL g11857 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data4[7]),
    .A2(n_330),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_1395));
 AOI22xp5_ASAP7_75t_SL g11858 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[0]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1394));
 AOI22xp5_ASAP7_75t_SL g11859 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[1]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1393));
 AOI22xp5_ASAP7_75t_SL g11860 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[2]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1392));
 AOI22xp5_ASAP7_75t_SL g11861 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[0]),
    .Y(n_1391));
 AOI22xp5_ASAP7_75t_SL g11862 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[3]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1390));
 AOI22xp5_ASAP7_75t_SL g11863 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[4]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1389));
 AOI22xp5_ASAP7_75t_SL g11864 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[1]),
    .Y(n_1388));
 AOI22xp5_ASAP7_75t_SL g11865 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[6]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1387));
 AOI22xp5_ASAP7_75t_SL g11866 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data5[7]),
    .A2(n_327),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_1386));
 AOI22xp5_ASAP7_75t_SL g11867 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[2]),
    .Y(n_1385));
 AOI22xp5_ASAP7_75t_SL g11868 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[7]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1384));
 AOI22xp5_ASAP7_75t_SL g11869 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[0]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1383));
 AOI22xp5_ASAP7_75t_SL g11870 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[6]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1382));
 AOI22xp5_ASAP7_75t_SL g11871 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[2]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1381));
 AOI22xp5_ASAP7_75t_SL g11872 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[3]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1380));
 AOI22xp5_ASAP7_75t_SL g11873 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[4]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1379));
 AOI22xp5_ASAP7_75t_SL g11874 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[5]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1378));
 AOI22xp5_ASAP7_75t_SL g11875 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[6]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1377));
 AOI22xp5_ASAP7_75t_SL g11876 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[3]),
    .Y(n_1376));
 AOI22xp5_ASAP7_75t_SL g11877 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[7]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1375));
 AOI22xp5_ASAP7_75t_SL g11878 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[2]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1374));
 AOI22xp5_ASAP7_75t_SL g11879 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[0]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1373));
 AOI22xp5_ASAP7_75t_SL g11880 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[4]),
    .Y(n_1372));
 AOI22xp5_ASAP7_75t_SL g11881 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[1]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1371));
 AOI22xp5_ASAP7_75t_SL g11882 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[1]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1370));
 AOI22xp5_ASAP7_75t_SL g11883 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[2]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1369));
 AOI22xp5_ASAP7_75t_SL g11884 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[3]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1368));
 AOI22xp5_ASAP7_75t_SL g11885 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[4]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1367));
 AOI22xp5_ASAP7_75t_SL g11886 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data7[5]),
    .A2(n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_1366));
 AOI22xp5_ASAP7_75t_SL g11887 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[5]),
    .Y(n_1365));
 AOI22xp5_ASAP7_75t_SL g11888 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[6]),
    .Y(n_1364));
 AOI22xp5_ASAP7_75t_SL g11889 (.A1(n_27),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[8]),
    .Y(n_1363));
 AOI22xp5_ASAP7_75t_SL g11890 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data0[3]),
    .A2(n_320),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_1362));
 AOI22xp5_ASAP7_75t_SL g11891 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[0]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1361));
 AOI22xp5_ASAP7_75t_SL g11892 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[1]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1360));
 AOI22xp5_ASAP7_75t_SL g11893 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[2]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1359));
 AOI22xp5_ASAP7_75t_SL g11894 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[3]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1358));
 AOI22xp5_ASAP7_75t_SL g11895 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[4]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1357));
 AOI22xp5_ASAP7_75t_SL g11896 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[5]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1356));
 AOI22xp5_ASAP7_75t_SL g11897 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[6]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1355));
 AOI22xp5_ASAP7_75t_SL g11898 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[0]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1354));
 AOI22xp5_ASAP7_75t_SL g11899 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[2]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1353));
 XNOR2xp5_ASAP7_75t_SL g119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_152),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_189),
    .Y(n_12616));
 AOI22xp5_ASAP7_75t_SL g11900 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[3]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1352));
 AOI22xp5_ASAP7_75t_SL g11901 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[4]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1351));
 AOI22xp5_ASAP7_75t_SL g11902 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[5]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1350));
 AOI22xp5_ASAP7_75t_SL g11903 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[6]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1349));
 AOI22xp5_ASAP7_75t_SL g11904 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[6]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1348));
 AOI22xp5_ASAP7_75t_SL g11905 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[0]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1347));
 AOI22xp5_ASAP7_75t_SL g11906 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[1]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1346));
 AOI22xp5_ASAP7_75t_SL g11907 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[2]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1345));
 AOI22xp5_ASAP7_75t_SL g11908 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[3]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1344));
 AOI22xp5_ASAP7_75t_SL g11909 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[5]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1343));
 AOI22xp5_ASAP7_75t_SL g11910 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[4]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1342));
 AOI22xp5_ASAP7_75t_SL g11911 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[5]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1341));
 AOI22xp5_ASAP7_75t_SL g11912 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[6]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[6]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1340));
 AOI22xp5_ASAP7_75t_SL g11913 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[4]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1339));
 AOI22xp5_ASAP7_75t_SL g11914 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[0]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1338));
 AOI22xp5_ASAP7_75t_SL g11915 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[2]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1337));
 AOI22xp5_ASAP7_75t_SL g11916 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[3]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1336));
 AOI22xp5_ASAP7_75t_SL g11917 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[1]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1335));
 AOI22xp5_ASAP7_75t_SL g11918 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data3[7]),
    .A2(n_319),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_1334));
 AOI22xp5_ASAP7_75t_SL g11919 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[4]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1333));
 AOI22xp5_ASAP7_75t_SL g11920 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data4[5]),
    .A2(n_323),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_1332));
 AOI22xp5_ASAP7_75t_SL g11921 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[2]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1331));
 AOI22xp5_ASAP7_75t_SL g11922 (.A1(u_NV_NVDLA_cmac_u_core_in_dat_data6[1]),
    .A2(n_318),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_1330));
 AOI22xp5_ASAP7_75t_SL g11923 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data5[3]),
    .A2(n_325),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_1329));
 AOI22xp5_ASAP7_75t_SL g11924 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[1]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1328));
 AOI22xp5_ASAP7_75t_SL g11925 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[2]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1327));
 AOI22xp5_ASAP7_75t_SL g11926 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[3]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1326));
 AOI22xp5_ASAP7_75t_SL g11927 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data2[7]),
    .A2(n_317),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_1325));
 AOI22xp5_ASAP7_75t_SL g11928 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[4]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[4]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1324));
 AOI22xp5_ASAP7_75t_SL g11929 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[5]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1323));
 AOI22xp5_ASAP7_75t_SL g11930 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data6[7]),
    .A2(n_321),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_1322));
 AOI22xp5_ASAP7_75t_SL g11931 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[0]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1321));
 AOI22xp5_ASAP7_75t_SL g11932 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[3]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1320));
 AOI22xp5_ASAP7_75t_SL g11933 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[5]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[5]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1319));
 AOI22xp5_ASAP7_75t_SL g11934 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data7[7]),
    .A2(n_326),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_1318));
 AOI22xp5_ASAP7_75t_SL g11935 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[7]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1317));
 AOI22xp5_ASAP7_75t_SL g11936 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data1[1]),
    .A2(n_316),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_1316));
 AOI22xp5_ASAP7_75t_SL g11937 (.A1(u_NV_NVDLA_cmac_u_core_in_wt_data0[7]),
    .A2(n_329),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[7]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_1315));
 AOI22xp5_ASAP7_75t_SL g11938 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[0]),
    .Y(n_1314));
 AOI22xp5_ASAP7_75t_SL g11939 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[1]),
    .Y(n_1313));
 AOI22xp5_ASAP7_75t_SL g11940 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[2]),
    .Y(n_1312));
 AOI22xp5_ASAP7_75t_SL g11941 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[3]),
    .Y(n_1311));
 AOI22xp5_ASAP7_75t_SL g11942 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[4]),
    .Y(n_1310));
 AOI22xp5_ASAP7_75t_SL g11943 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[5]),
    .Y(n_1309));
 AOI22xp5_ASAP7_75t_SL g11944 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[6]),
    .Y(n_1308));
 AOI22xp5_ASAP7_75t_SL g11945 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .A2(n_26),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[7]),
    .Y(n_1307));
 AOI22xp33_ASAP7_75t_SL g11946 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[0]),
    .Y(n_1306));
 AOI22xp33_ASAP7_75t_SL g11947 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[1]),
    .Y(n_1305));
 AOI22xp33_ASAP7_75t_SL g11948 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[2]),
    .Y(n_1304));
 AOI22xp33_ASAP7_75t_SL g11949 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[3]),
    .Y(n_1303));
 AOI22xp33_ASAP7_75t_SL g11950 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[4]),
    .Y(n_1302));
 AOI22xp33_ASAP7_75t_SL g11951 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[5]),
    .Y(n_1301));
 AOI22xp33_ASAP7_75t_SL g11952 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[6]),
    .Y(n_1300));
 AOI22xp33_ASAP7_75t_SL g11953 (.A1(n_25),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_wt_mask[7]),
    .Y(n_1299));
 AOI22xp33_ASAP7_75t_SL g11954 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[0]),
    .Y(n_1298));
 AOI22xp5_ASAP7_75t_SL g11955 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[6]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[6]),
    .Y(n_1297));
 AOI22xp5_ASAP7_75t_SL g11956 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[34]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[34]),
    .Y(n_1296));
 AOI22xp5_ASAP7_75t_SL g11957 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[9]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[9]),
    .Y(n_1295));
 AOI22xp5_ASAP7_75t_SL g11958 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[54]),
    .Y(n_1294));
 AOI22xp5_ASAP7_75t_SL g11959 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[22]),
    .Y(n_1293));
 AOI22xp5_ASAP7_75t_SL g11960 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[2]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[2]),
    .Y(n_1292));
 AOI22xp5_ASAP7_75t_SL g11961 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[5]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[5]),
    .Y(n_1291));
 AOI22xp5_ASAP7_75t_SL g11962 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[35]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[35]),
    .Y(n_1290));
 AOI22xp5_ASAP7_75t_SL g11963 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[55]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[55]),
    .Y(n_1289));
 AOI22xp5_ASAP7_75t_SL g11964 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[4]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[4]),
    .Y(n_1288));
 AOI22xp5_ASAP7_75t_SL g11965 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[3]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[3]),
    .Y(n_1287));
 AOI22xp5_ASAP7_75t_SL g11966 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[1]),
    .Y(n_1286));
 AOI22xp5_ASAP7_75t_SL g11967 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[7]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[7]),
    .Y(n_1285));
 AOI22xp5_ASAP7_75t_SL g11968 (.A1(n_24),
    .A2(u_NV_NVDLA_cmac_u_reg_req_pd[8]),
    .B1(csb2cmac_a_req_pvld),
    .B2(csb2cmac_a_req_pd[8]),
    .Y(n_1284));
 AOI22xp5_ASAP7_75t_SL g11969 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[6]),
    .Y(n_1283));
 AOI22xp5_ASAP7_75t_SL g11970 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[1]),
    .Y(n_1282));
 AOI22xp5_ASAP7_75t_SL g11971 (.A1(mac2accu_data3[7]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[7]),
    .Y(n_1281));
 AOI22xp5_ASAP7_75t_SL g11972 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[18]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[18]),
    .Y(n_1280));
 AOI22xp5_ASAP7_75t_SL g11973 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[16]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[16]),
    .Y(n_1279));
 AOI22xp5_ASAP7_75t_SL g11974 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[15]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[15]),
    .Y(n_1278));
 AOI22xp5_ASAP7_75t_SL g11975 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[10]),
    .Y(n_1277));
 AOI22xp5_ASAP7_75t_SL g11976 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[9]),
    .Y(n_1276));
 AOI22xp5_ASAP7_75t_SL g11977 (.A1(mac2accu_data3[18]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[18]),
    .Y(n_1275));
 AOI22xp5_ASAP7_75t_SL g11978 (.A1(mac2accu_data3[16]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[16]),
    .Y(n_1274));
 AOI22xp5_ASAP7_75t_SL g11979 (.A1(mac2accu_data3[15]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[15]),
    .Y(n_1273));
 AOI22xp5_ASAP7_75t_SL g11981 (.A1(mac2accu_data3[12]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[12]),
    .Y(n_1271));
 AOI22xp5_ASAP7_75t_SL g11982 (.A1(mac2accu_data3[13]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[13]),
    .Y(n_1270));
 AOI22xp5_ASAP7_75t_SL g11984 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[12]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[12]),
    .Y(n_1268));
 AOI22xp5_ASAP7_75t_SL g11985 (.A1(mac2accu_data3[10]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[10]),
    .Y(n_1267));
 AOI22xp5_ASAP7_75t_SL g11986 (.A1(mac2accu_data3[9]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[9]),
    .Y(n_1266));
 AOI22xp5_ASAP7_75t_SL g11987 (.A1(mac2accu_data3[6]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[6]),
    .Y(n_1265));
 AOI22xp5_ASAP7_75t_SL g11988 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_173),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[3]),
    .B2(n_17876),
    .Y(n_1264));
 AOI22xp5_ASAP7_75t_SL g11989 (.A1(mac2accu_data3[4]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[4]),
    .Y(n_1263));
 AOI22xp5_ASAP7_75t_SL g11990 (.A1(mac2accu_data3[3]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[3]),
    .Y(n_1262));
 AOI22xp5_ASAP7_75t_SL g11991 (.A1(mac2accu_data3[0]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[0]),
    .Y(n_1261));
 AOI22xp5_ASAP7_75t_SL g11992 (.A1(mac2accu_data3[1]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[1]),
    .Y(n_1260));
 AOI22xp5_ASAP7_75t_SL g11993 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[17]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[17]),
    .Y(n_1259));
 AOI22xp5_ASAP7_75t_SL g11994 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[14]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[14]),
    .Y(n_1258));
 AOI22xp5_ASAP7_75t_SL g11995 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[15]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[15]),
    .Y(n_1257));
 AOI22xp5_ASAP7_75t_SL g11996 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[13]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[13]),
    .Y(n_1256));
 AOI22xp5_ASAP7_75t_SL g11997 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[11]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[11]),
    .Y(n_1255));
 AOI22xp5_ASAP7_75t_SL g11998 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[8]),
    .Y(n_1254));
 AOI22xp5_ASAP7_75t_SL g11999 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[9]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[9]),
    .Y(n_1253));
 AND2x2_ASAP7_75t_SRAM g12 (.A(n_3112),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(n_14029));
 OAI21x1_ASAP7_75t_SL g120 (.A1(n_5491),
    .A2(n_5492),
    .B(n_5493),
    .Y(n_5494));
 AOI22xp5_ASAP7_75t_SL g12000 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[5]),
    .Y(n_1252));
 AOI22xp5_ASAP7_75t_SL g12001 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[7]),
    .Y(n_1251));
 AOI22xp5_ASAP7_75t_SL g12003 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_171),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[1]),
    .B2(n_17870),
    .Y(n_1249));
 AOI22xp5_ASAP7_75t_SL g12004 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[7]),
    .Y(n_1248));
 AOI22xp5_ASAP7_75t_SL g12005 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_172),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[2]),
    .B2(n_17870),
    .Y(n_1247));
 AOI22xp5_ASAP7_75t_SL g12006 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_173),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[3]),
    .B2(n_17870),
    .Y(n_1246));
 AOI22xp5_ASAP7_75t_SL g12007 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_174),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[4]),
    .B2(n_17870),
    .Y(n_1245));
 AOI22xp5_ASAP7_75t_SL g12008 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[6]),
    .Y(n_1244));
 AOI22xp5_ASAP7_75t_SL g12009 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_175),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[5]),
    .B2(n_17870),
    .Y(n_1243));
 AOI22xp5_ASAP7_75t_SL g12010 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_176),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[6]),
    .Y(n_1242));
 AOI22xp5_ASAP7_75t_SL g12011 (.A1(n_17869),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_n_177),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[7]),
    .Y(n_1241));
 AOI22xp5_ASAP7_75t_SL g12012 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_n_178),
    .A2(n_17869),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[8]),
    .Y(n_1240));
 AOI22xp5_ASAP7_75t_SL g12014 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_n_180),
    .A2(n_17869),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[10]),
    .Y(n_1238));
 AOI22xp5_ASAP7_75t_SL g12015 (.A1(n_16597),
    .A2(n_17869),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[11]),
    .Y(n_1237));
 AOI22xp5_ASAP7_75t_SL g12016 (.A1(n_17869),
    .A2(n_18804),
    .B1(n_17870),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[12]),
    .Y(n_1236));
 AOI22xp5_ASAP7_75t_SL g12023 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[0]),
    .Y(n_1230));
 AOI22xp5_ASAP7_75t_SL g12024 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[1]),
    .Y(n_1229));
 AOI22xp5_ASAP7_75t_SL g12025 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[2]),
    .Y(n_1228));
 AOI22xp5_ASAP7_75t_SL g12027 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[4]),
    .Y(n_1226));
 AOI22xp5_ASAP7_75t_SL g12028 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[3]),
    .Y(n_1225));
 AOI22xp5_ASAP7_75t_SL g12029 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[5]),
    .Y(n_1224));
 AOI22xp5_ASAP7_75t_SL g12030 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[16]),
    .Y(n_1223));
 AOI22xp5_ASAP7_75t_SL g12031 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[6]),
    .Y(n_1222));
 AOI22xp5_ASAP7_75t_SL g12032 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[7]),
    .Y(n_1221));
 AOI22xp5_ASAP7_75t_SL g12033 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[8]),
    .Y(n_1220));
 AOI22xp5_ASAP7_75t_SL g12034 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[2]),
    .Y(n_1219));
 AOI22xp5_ASAP7_75t_SL g12035 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[9]),
    .Y(n_1218));
 AOI22xp5_ASAP7_75t_SL g12036 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[10]),
    .Y(n_1217));
 AOI22xp5_ASAP7_75t_SL g12037 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[11]),
    .Y(n_1216));
 AOI22xp5_ASAP7_75t_SL g12038 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[12]),
    .Y(n_1215));
 AOI22xp5_ASAP7_75t_SL g12039 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[13]),
    .Y(n_1214));
 AOI22xp5_ASAP7_75t_SL g12040 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[14]),
    .Y(n_1213));
 AOI22xp5_ASAP7_75t_SL g12041 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[15]),
    .Y(n_1212));
 AOI22xp5_ASAP7_75t_SL g12042 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[16]),
    .Y(n_1211));
 AOI22xp5_ASAP7_75t_SL g12043 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[17]),
    .Y(n_1210));
 AOI22xp5_ASAP7_75t_SL g12044 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[18]),
    .Y(n_1209));
 AOI22xp5_ASAP7_75t_SL g12045 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[0]),
    .Y(n_1208));
 AOI22xp5_ASAP7_75t_SL g12046 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[1]),
    .Y(n_1207));
 AOI22xp5_ASAP7_75t_SL g12047 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[2]),
    .Y(n_1206));
 AOI22xp5_ASAP7_75t_SL g12048 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[3]),
    .Y(n_1205));
 AOI22xp5_ASAP7_75t_SL g12049 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[4]),
    .Y(n_1204));
 AOI22xp5_ASAP7_75t_SL g12050 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[5]),
    .Y(n_1203));
 AOI22xp5_ASAP7_75t_SL g12051 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[6]),
    .Y(n_1202));
 AOI22xp5_ASAP7_75t_SL g12052 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[7]),
    .Y(n_1201));
 AOI22xp5_ASAP7_75t_SL g12053 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[8]),
    .Y(n_1200));
 AOI22xp5_ASAP7_75t_SL g12054 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[9]),
    .Y(n_1199));
 AOI22xp5_ASAP7_75t_SL g12055 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[0]),
    .Y(n_1198));
 AOI22xp5_ASAP7_75t_SL g12056 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[10]),
    .Y(n_1197));
 AOI22xp5_ASAP7_75t_SL g12057 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[11]),
    .Y(n_1196));
 AOI22xp5_ASAP7_75t_SL g12058 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[12]),
    .Y(n_1195));
 AOI22xp5_ASAP7_75t_SL g12059 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[13]),
    .Y(n_1194));
 AOI22xp5_ASAP7_75t_SL g12060 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[14]),
    .Y(n_1193));
 AOI22xp5_ASAP7_75t_SL g12061 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[15]),
    .Y(n_1192));
 AOI22xp5_ASAP7_75t_SL g12062 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[16]),
    .Y(n_1191));
 AOI22xp5_ASAP7_75t_SL g12063 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[17]),
    .Y(n_1190));
 AOI22xp5_ASAP7_75t_SL g12064 (.A1(n_13),
    .A2(u_NV_NVDLA_cmac_u_core_out_data0[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[18]),
    .Y(n_1189));
 AOI22xp5_ASAP7_75t_SL g12065 (.A1(n_17936),
    .A2(n_19083),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[0]),
    .B2(n_5332),
    .Y(n_1188));
 AOI22xp5_ASAP7_75t_SL g12066 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_171),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[1]),
    .B2(n_5332),
    .Y(n_1187));
 AOI22xp5_ASAP7_75t_SL g12067 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_172),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[2]),
    .B2(n_5332),
    .Y(n_1186));
 AOI22xp5_ASAP7_75t_SL g12068 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_173),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[3]),
    .B2(n_5332),
    .Y(n_1185));
 AOI22xp5_ASAP7_75t_SL g12069 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_174),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[4]),
    .B2(n_5332),
    .Y(n_1184));
 AOI22xp5_ASAP7_75t_SL g12070 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_175),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[5]),
    .B2(n_5332),
    .Y(n_1183));
 AOI22xp5_ASAP7_75t_SL g12071 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_176),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[6]),
    .Y(n_1182));
 AOI22xp5_ASAP7_75t_SL g12072 (.A1(n_17936),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_177),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[7]),
    .Y(n_1181));
 AOI22xp5_ASAP7_75t_SL g12073 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_n_178),
    .A2(n_17936),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[8]),
    .Y(n_1180));
 AOI22xp5_ASAP7_75t_SL g12075 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_n_180),
    .A2(n_17936),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[10]),
    .Y(n_1178));
 AOI22xp5_ASAP7_75t_SL g12077 (.A1(n_20741),
    .A2(n_17936),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[12]),
    .Y(n_1176));
 AOI22xp5_ASAP7_75t_SL g12084 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[0]),
    .Y(n_1169));
 AOI22xp5_ASAP7_75t_SL g12085 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[1]),
    .Y(n_1168));
 AOI22xp5_ASAP7_75t_SL g12086 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[2]),
    .Y(n_1167));
 AOI22xp5_ASAP7_75t_SL g12087 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[3]),
    .Y(n_1166));
 AOI22xp5_ASAP7_75t_SL g12088 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[4]),
    .Y(n_1165));
 AOI22xp5_ASAP7_75t_SL g12089 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[5]),
    .Y(n_1164));
 AOI22xp5_ASAP7_75t_SL g12090 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[6]),
    .Y(n_1163));
 AOI22xp5_ASAP7_75t_SL g12091 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[7]),
    .Y(n_1162));
 AOI22xp5_ASAP7_75t_SL g12092 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[8]),
    .Y(n_1161));
 AOI22xp5_ASAP7_75t_SL g12093 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[9]),
    .Y(n_1160));
 AOI22xp5_ASAP7_75t_SL g12094 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[10]),
    .Y(n_1159));
 AOI22xp5_ASAP7_75t_SL g12095 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[11]),
    .Y(n_1158));
 AOI22xp5_ASAP7_75t_SL g12096 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[12]),
    .Y(n_1157));
 AOI22xp5_ASAP7_75t_SL g12097 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[13]),
    .Y(n_1156));
 AOI22xp5_ASAP7_75t_SL g12098 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[7]),
    .Y(n_1155));
 AOI22xp5_ASAP7_75t_SL g12099 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[14]),
    .Y(n_1154));
 OR2x2_ASAP7_75t_SL g121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_581),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_677),
    .Y(n_5493));
 AOI22xp5_ASAP7_75t_SL g12100 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[15]),
    .Y(n_1153));
 AOI22xp5_ASAP7_75t_SL g12101 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[16]),
    .Y(n_1152));
 AOI22xp5_ASAP7_75t_SL g12102 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[17]),
    .Y(n_1151));
 AOI22xp5_ASAP7_75t_SL g12103 (.A1(n_15),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[18]),
    .Y(n_1150));
 AOI22xp5_ASAP7_75t_SL g12104 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[2]),
    .Y(n_1149));
 AOI22xp5_ASAP7_75t_SL g12105 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[0]),
    .Y(n_1148));
 AOI22xp5_ASAP7_75t_SL g12106 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[1]),
    .Y(n_1147));
 AOI22xp5_ASAP7_75t_SL g12107 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[2]),
    .Y(n_1146));
 AOI22xp5_ASAP7_75t_SL g12109 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[3]),
    .Y(n_1144));
 AOI22xp5_ASAP7_75t_SL g12110 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[9]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[9]),
    .Y(n_1143));
 AOI22xp5_ASAP7_75t_SL g12111 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[4]),
    .Y(n_1142));
 AOI22xp5_ASAP7_75t_SL g12112 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[5]),
    .Y(n_1141));
 AOI22xp5_ASAP7_75t_SL g12113 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[6]),
    .Y(n_1140));
 AOI22xp5_ASAP7_75t_SL g12114 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[7]),
    .Y(n_1139));
 AOI22xp5_ASAP7_75t_SL g12115 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[8]),
    .Y(n_1138));
 AOI22xp5_ASAP7_75t_SL g12116 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[9]),
    .Y(n_1137));
 AOI22xp5_ASAP7_75t_SL g12117 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[10]),
    .Y(n_1136));
 AOI22xp5_ASAP7_75t_SL g12118 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[11]),
    .Y(n_1135));
 AOI22xp5_ASAP7_75t_SL g12119 (.A1(mac2accu_data2[11]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[11]),
    .Y(n_1134));
 AOI22xp5_ASAP7_75t_SL g12120 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[12]),
    .Y(n_1133));
 AOI22xp5_ASAP7_75t_SL g12121 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[13]),
    .Y(n_1132));
 AOI22xp5_ASAP7_75t_SL g12122 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[14]),
    .Y(n_1131));
 AOI22xp5_ASAP7_75t_SL g12123 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[15]),
    .Y(n_1130));
 AOI22xp5_ASAP7_75t_SL g12124 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[16]),
    .Y(n_1129));
 AOI22xp5_ASAP7_75t_SL g12125 (.A1(mac2accu_data2[9]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[9]),
    .Y(n_1128));
 AOI22xp5_ASAP7_75t_SL g12126 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[17]),
    .Y(n_1127));
 AOI22xp5_ASAP7_75t_SL g12127 (.A1(n_10),
    .A2(u_NV_NVDLA_cmac_u_core_out_data1[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[18]),
    .Y(n_1126));
 AOI22xp5_ASAP7_75t_SL g12129 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_171),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[1]),
    .B2(n_17882),
    .Y(n_1124));
 A2O1A1Ixp33_ASAP7_75t_SL g1213 (.A1(n_19377),
    .A2(n_15816),
    .B(n_12676),
    .C(n_19378),
    .Y(n_12680));
 AOI22xp5_ASAP7_75t_SL g12130 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_172),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[2]),
    .B2(n_17882),
    .Y(n_1123));
 AOI22xp5_ASAP7_75t_SL g12131 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_173),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[3]),
    .B2(n_17882),
    .Y(n_1122));
 AOI22xp5_ASAP7_75t_SL g12132 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_174),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[4]),
    .B2(n_17882),
    .Y(n_1121));
 AOI22xp5_ASAP7_75t_SL g12133 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_175),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[5]),
    .B2(n_17882),
    .Y(n_1120));
 AOI22xp5_ASAP7_75t_SL g12134 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_176),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[6]),
    .Y(n_1119));
 AOI22xp5_ASAP7_75t_SL g12135 (.A1(n_23932),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_n_177),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[7]),
    .Y(n_1118));
 AOI22xp5_ASAP7_75t_SL g12136 (.A1(n_17077),
    .A2(n_23932),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[8]),
    .Y(n_1117));
 AOI22xp5_ASAP7_75t_SL g12137 (.A1(n_23932),
    .A2(n_26256),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[9]),
    .Y(n_1116));
 AOI22xp5_ASAP7_75t_SL g12138 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_n_180),
    .A2(n_23932),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[10]),
    .Y(n_1115));
 OAI21xp5_ASAP7_75t_SL g1214 (.A1(n_12667),
    .A2(n_12669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_280),
    .Y(n_12676));
 AOI22xp5_ASAP7_75t_SL g12142 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_n_184),
    .A2(n_23932),
    .B1(n_17882),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[14]),
    .Y(n_1111));
 AOI22xp5_ASAP7_75t_SL g12146 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[0]),
    .Y(n_1107));
 AOI22xp5_ASAP7_75t_SL g12147 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[1]),
    .Y(n_1106));
 AOI22xp5_ASAP7_75t_SL g12148 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[3]),
    .Y(n_1105));
 AOI22xp5_ASAP7_75t_SL g12149 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[4]),
    .Y(n_1104));
 AOI22xp5_ASAP7_75t_SL g12150 (.A1(mac2accu_data2[5]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[5]),
    .Y(n_1103));
 AOI22xp5_ASAP7_75t_SL g12151 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[5]),
    .Y(n_1102));
 AOI22xp5_ASAP7_75t_SL g12152 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[6]),
    .Y(n_1101));
 AOI22xp5_ASAP7_75t_SL g12153 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[7]),
    .Y(n_1100));
 AOI22xp5_ASAP7_75t_SL g12154 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[8]),
    .Y(n_1099));
 AOI22xp5_ASAP7_75t_SL g12155 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[9]),
    .Y(n_1098));
 AOI22xp5_ASAP7_75t_SL g12156 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[10]),
    .Y(n_1097));
 AOI22xp5_ASAP7_75t_SL g12157 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[11]),
    .Y(n_1096));
 AOI22xp5_ASAP7_75t_SL g12158 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[12]),
    .Y(n_1095));
 AOI22xp5_ASAP7_75t_SL g12159 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[13]),
    .Y(n_1094));
 AOI22xp5_ASAP7_75t_SL g12160 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[14]),
    .Y(n_1093));
 AOI22xp5_ASAP7_75t_SL g12161 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[15]),
    .Y(n_1092));
 AOI22xp5_ASAP7_75t_SL g12162 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[17]),
    .Y(n_1091));
 AOI22xp5_ASAP7_75t_SL g12163 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[11]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[11]),
    .Y(n_1090));
 AOI22xp5_ASAP7_75t_SL g12164 (.A1(n_4),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[18]),
    .Y(n_1089));
 AOI22xp5_ASAP7_75t_SL g12165 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[0]),
    .Y(n_1088));
 AOI22xp5_ASAP7_75t_SL g12166 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[1]),
    .Y(n_1087));
 AOI22xp5_ASAP7_75t_SL g12167 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[2]),
    .Y(n_1086));
 AOI22xp5_ASAP7_75t_SL g12168 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[3]),
    .Y(n_1085));
 AOI22xp5_ASAP7_75t_SL g12169 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[4]),
    .Y(n_1084));
 NAND2xp5_ASAP7_75t_SL g1217 (.A(n_12672),
    .B(n_12674),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_280));
 AOI22xp5_ASAP7_75t_SL g12170 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[5]),
    .Y(n_1083));
 AOI22xp5_ASAP7_75t_SL g12171 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[6]),
    .Y(n_1082));
 AOI22xp5_ASAP7_75t_SL g12172 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[7]),
    .Y(n_1081));
 AOI22xp5_ASAP7_75t_SL g12173 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[8]),
    .Y(n_1080));
 AOI22xp5_ASAP7_75t_SL g12174 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[9]),
    .Y(n_1079));
 AOI22xp5_ASAP7_75t_SL g12175 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[10]),
    .Y(n_1078));
 AOI22xp5_ASAP7_75t_SL g12176 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[11]),
    .Y(n_1077));
 AOI22xp5_ASAP7_75t_SL g12177 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[12]),
    .Y(n_1076));
 AOI22xp5_ASAP7_75t_SL g12178 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[13]),
    .Y(n_1075));
 AOI22xp5_ASAP7_75t_SL g12179 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[14]),
    .Y(n_1074));
 NOR2xp33_ASAP7_75t_SL g1218 (.A(n_12667),
    .B(n_12669),
    .Y(n_12681));
 AOI22xp5_ASAP7_75t_SL g12180 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[15]),
    .Y(n_1073));
 AOI22xp5_ASAP7_75t_SL g12181 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[16]),
    .Y(n_1072));
 AOI22xp5_ASAP7_75t_SL g12182 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[17]),
    .Y(n_1071));
 AOI22xp5_ASAP7_75t_SL g12183 (.A1(n_5),
    .A2(u_NV_NVDLA_cmac_u_core_out_data2[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[18]),
    .Y(n_1070));
 AOI22xp5_ASAP7_75t_SL g12185 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_171),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[1]),
    .B2(n_17876),
    .Y(n_1068));
 AOI22xp5_ASAP7_75t_SL g12186 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_172),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[2]),
    .B2(n_17876),
    .Y(n_1067));
 AOI22xp5_ASAP7_75t_SL g12187 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_174),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[4]),
    .B2(n_17876),
    .Y(n_1066));
 AOI22xp5_ASAP7_75t_SL g12188 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_175),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[5]),
    .B2(n_17876),
    .Y(n_1065));
 AOI22xp5_ASAP7_75t_SL g12189 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_176),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[6]),
    .Y(n_1064));
 AOI22xp5_ASAP7_75t_SL g12190 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_177),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[7]),
    .Y(n_1063));
 AOI22xp5_ASAP7_75t_SL g12191 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[17]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[17]),
    .Y(n_1062));
 AOI22xp5_ASAP7_75t_SL g12192 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_n_178),
    .A2(n_17874),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[8]),
    .Y(n_1061));
 AOI22xp5_ASAP7_75t_SL g12194 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_181),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[11]),
    .Y(n_1059));
 AOI22xp5_ASAP7_75t_SL g12195 (.A1(n_17874),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_182),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[12]),
    .Y(n_1058));
 AOI22xp5_ASAP7_75t_SL g12196 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[12]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[12]),
    .Y(n_1057));
 AOI22xp5_ASAP7_75t_SL g12197 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_n_184),
    .A2(n_17874),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[14]),
    .Y(n_1056));
 AOI22xp5_ASAP7_75t_SL g12198 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[16]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[16]),
    .Y(n_1055));
 AND2x2_ASAP7_75t_SL g122 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_677),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_581),
    .Y(n_5491));
 AOI22xp5_ASAP7_75t_SL g12203 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[0]),
    .Y(n_1050));
 AOI22xp5_ASAP7_75t_SL g12204 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[1]),
    .Y(n_1049));
 AOI22xp5_ASAP7_75t_SL g12205 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[2]),
    .Y(n_1048));
 AOI22xp5_ASAP7_75t_SL g12206 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[3]),
    .Y(n_1047));
 AOI22xp5_ASAP7_75t_SL g12207 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[4]),
    .Y(n_1046));
 AOI22xp5_ASAP7_75t_SL g12208 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[5]),
    .Y(n_1045));
 AOI22xp5_ASAP7_75t_SL g12209 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[6]),
    .Y(n_1044));
 MAJIxp5_ASAP7_75t_SL g1221 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_239),
    .B(n_13575),
    .C(n_25503),
    .Y(n_12672));
 AOI22xp5_ASAP7_75t_SL g12210 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[7]),
    .Y(n_1043));
 AOI22xp5_ASAP7_75t_SL g12211 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[8]),
    .Y(n_1042));
 AOI22xp5_ASAP7_75t_SL g12212 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[14]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[14]),
    .Y(n_1041));
 AOI22xp5_ASAP7_75t_SL g12213 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[11]),
    .Y(n_1040));
 AOI22xp5_ASAP7_75t_SL g12214 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[12]),
    .Y(n_1039));
 AOI22xp5_ASAP7_75t_SL g12215 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[13]),
    .Y(n_1038));
 AOI22xp5_ASAP7_75t_SL g12216 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[14]),
    .Y(n_1037));
 AOI22xp5_ASAP7_75t_SL g12217 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[15]),
    .Y(n_1036));
 AOI22xp5_ASAP7_75t_SL g12218 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[16]),
    .Y(n_1035));
 AOI22xp5_ASAP7_75t_SL g12219 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[17]),
    .Y(n_1034));
 MAJIxp5_ASAP7_75t_SL g1222 (.A(n_25504),
    .B(n_9452),
    .C(n_9453),
    .Y(n_12667));
 AOI22xp5_ASAP7_75t_SL g12220 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[12]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[12]),
    .Y(n_1033));
 AOI22xp5_ASAP7_75t_SL g12221 (.A1(n_18),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[18]),
    .Y(n_1032));
 AOI22xp5_ASAP7_75t_SL g12222 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[0]),
    .Y(n_1031));
 AOI22xp5_ASAP7_75t_SL g12223 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[1]),
    .Y(n_1030));
 AOI22xp5_ASAP7_75t_SL g12224 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[2]),
    .Y(n_1029));
 AOI22xp5_ASAP7_75t_SL g12225 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[3]),
    .Y(n_1028));
 AOI22xp5_ASAP7_75t_SL g12226 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[4]),
    .Y(n_1027));
 AOI22xp5_ASAP7_75t_SL g12227 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[5]),
    .Y(n_1026));
 AOI22xp5_ASAP7_75t_SL g12228 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[9]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[9]),
    .Y(n_1025));
 AOI22xp5_ASAP7_75t_SL g12229 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[6]),
    .Y(n_1024));
 AOI22xp5_ASAP7_75t_SL g12230 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[7]),
    .Y(n_1023));
 AOI22xp5_ASAP7_75t_SL g12231 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[8]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[8]),
    .Y(n_1022));
 AOI22xp5_ASAP7_75t_SL g12232 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[9]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[9]),
    .Y(n_1021));
 AOI22xp5_ASAP7_75t_SL g12233 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[11]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[11]),
    .Y(n_1020));
 AOI22xp5_ASAP7_75t_SL g12234 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[12]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[12]),
    .Y(n_1019));
 AOI22xp5_ASAP7_75t_SL g12235 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[13]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[13]),
    .Y(n_1018));
 AOI22xp5_ASAP7_75t_SL g12236 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[14]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[14]),
    .Y(n_1017));
 AOI22xp5_ASAP7_75t_SL g12237 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[15]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[15]),
    .Y(n_1016));
 AOI22xp5_ASAP7_75t_SL g12238 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[16]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[16]),
    .Y(n_1015));
 AOI22xp5_ASAP7_75t_SL g12239 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[17]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[17]),
    .Y(n_1014));
 XOR2x2_ASAP7_75t_SL g1224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_250),
    .B(n_25503),
    .Y(n_12669));
 AOI22xp5_ASAP7_75t_SL g12240 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[18]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[18]),
    .Y(n_1013));
 AOI22xp5_ASAP7_75t_SL g12241 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[3]),
    .Y(n_1012));
 AOI22xp5_ASAP7_75t_SL g12242 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[2]),
    .Y(n_1011));
 AOI22xp5_ASAP7_75t_SL g12243 (.A1(mac2accu_data0[0]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[0]),
    .Y(n_1010));
 AOI22xp5_ASAP7_75t_SL g12244 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[4]),
    .Y(n_1009));
 AOI22xp5_ASAP7_75t_SL g12245 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[4]),
    .Y(n_1008));
 AOI22xp5_ASAP7_75t_SL g12246 (.A1(mac2accu_data1[18]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[18]),
    .Y(n_1007));
 AOI22xp5_ASAP7_75t_SL g12247 (.A1(mac2accu_data1[17]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[17]),
    .Y(n_1006));
 AOI22xp5_ASAP7_75t_SL g12248 (.A1(mac2accu_data1[15]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[15]),
    .Y(n_1005));
 AOI22xp5_ASAP7_75t_SL g12249 (.A1(mac2accu_data1[12]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[12]),
    .Y(n_1004));
 AOI22xp5_ASAP7_75t_SL g12250 (.A1(mac2accu_data1[11]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[11]),
    .Y(n_1003));
 AOI22xp5_ASAP7_75t_SL g12251 (.A1(mac2accu_data1[6]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[6]),
    .Y(n_1002));
 AOI22xp5_ASAP7_75t_SL g12252 (.A1(mac2accu_data1[9]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[9]),
    .Y(n_1001));
 AOI22xp5_ASAP7_75t_SL g12253 (.A1(mac2accu_data1[8]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[8]),
    .Y(n_1000));
 AOI22xp5_ASAP7_75t_SL g12254 (.A1(mac2accu_data1[0]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[0]),
    .Y(n_999));
 AOI22xp5_ASAP7_75t_SL g12255 (.A1(mac2accu_data1[2]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[2]),
    .Y(n_998));
 AOI22xp5_ASAP7_75t_SL g12256 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[17]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[17]),
    .Y(n_997));
 AOI22xp5_ASAP7_75t_SL g12257 (.A1(mac2accu_data1[3]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[3]),
    .Y(n_996));
 AOI22xp5_ASAP7_75t_SL g12258 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[8]),
    .Y(n_995));
 AOI22xp5_ASAP7_75t_SL g12259 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[18]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[18]),
    .Y(n_994));
 XNOR2x1_ASAP7_75t_SL g1226 (.B(n_18786),
    .Y(n_12674),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_15));
 AOI22xp5_ASAP7_75t_SL g12260 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[13]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[13]),
    .Y(n_993));
 AOI22xp5_ASAP7_75t_SL g12261 (.A1(n_12),
    .A2(u_NV_NVDLA_cmac_u_core_out_data3[10]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[10]),
    .Y(n_992));
 AOI22xp5_ASAP7_75t_SL g12262 (.A1(mac2accu_data1[14]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[14]),
    .Y(n_991));
 AOI22xp5_ASAP7_75t_SL g12263 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[0]),
    .Y(n_990));
 AOI22xp5_ASAP7_75t_SL g12264 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[1]),
    .Y(n_989));
 AOI22xp5_ASAP7_75t_SL g12265 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[5]),
    .Y(n_988));
 AOI22xp5_ASAP7_75t_SL g12266 (.A1(mac2accu_data1[16]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[16]),
    .Y(n_987));
 AOI22xp5_ASAP7_75t_SL g12267 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[5]),
    .Y(n_986));
 AOI22xp5_ASAP7_75t_SL g12268 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[9]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[9]),
    .Y(n_985));
 AOI22xp5_ASAP7_75t_SL g12269 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[10]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[10]),
    .Y(n_984));
 AOI22xp5_ASAP7_75t_SL g12270 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[11]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[11]),
    .Y(n_983));
 AOI22xp5_ASAP7_75t_SL g12271 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[2]),
    .Y(n_982));
 AOI22xp5_ASAP7_75t_SL g12272 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[13]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[13]),
    .Y(n_981));
 AOI22xp5_ASAP7_75t_SL g12273 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[14]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[14]),
    .Y(n_980));
 AOI22xp5_ASAP7_75t_SL g12274 (.A1(n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[17]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data0[17]),
    .Y(n_979));
 AOI22xp5_ASAP7_75t_SL g12275 (.A1(mac2accu_data0[7]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[7]),
    .Y(n_978));
 AOI22xp5_ASAP7_75t_SL g12276 (.A1(mac2accu_data0[8]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[8]),
    .Y(n_977));
 AOI22xp5_ASAP7_75t_SL g12277 (.A1(mac2accu_data0[9]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[9]),
    .Y(n_976));
 AOI22xp5_ASAP7_75t_SL g12278 (.A1(mac2accu_data0[10]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[10]),
    .Y(n_975));
 AOI22xp5_ASAP7_75t_SL g12279 (.A1(mac2accu_data0[11]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[11]),
    .Y(n_974));
 AOI22xp5_ASAP7_75t_SL g12280 (.A1(mac2accu_data0[12]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[12]),
    .Y(n_973));
 AOI22xp5_ASAP7_75t_SL g12281 (.A1(mac2accu_data0[13]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[13]),
    .Y(n_972));
 AOI22xp5_ASAP7_75t_SL g12282 (.A1(mac2accu_data0[14]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[14]),
    .Y(n_971));
 AOI22xp5_ASAP7_75t_SL g12283 (.A1(mac2accu_data0[15]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[15]),
    .Y(n_970));
 AOI22xp5_ASAP7_75t_SL g12284 (.A1(mac2accu_data0[16]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[16]),
    .Y(n_969));
 AOI22xp5_ASAP7_75t_SL g12285 (.A1(mac2accu_data0[17]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[17]),
    .Y(n_968));
 AOI22xp5_ASAP7_75t_SL g12286 (.A1(mac2accu_data0[18]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[18]),
    .Y(n_967));
 AOI22xp5_ASAP7_75t_SL g12287 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[0]),
    .Y(n_966));
 AOI22xp5_ASAP7_75t_SL g12288 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[1]),
    .Y(n_965));
 AOI22xp5_ASAP7_75t_SL g12289 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[2]),
    .Y(n_964));
 AOI22xp5_ASAP7_75t_SL g12290 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[3]),
    .Y(n_963));
 AOI22xp5_ASAP7_75t_SL g12291 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[4]),
    .Y(n_962));
 AOI22xp5_ASAP7_75t_SL g12292 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[6]),
    .Y(n_961));
 AOI22xp5_ASAP7_75t_SL g12293 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[8]),
    .Y(n_960));
 AOI22xp5_ASAP7_75t_SL g12294 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[10]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[10]),
    .Y(n_959));
 AOI22xp5_ASAP7_75t_SL g12295 (.A1(mac2accu_data1[5]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[5]),
    .Y(n_958));
 AOI22xp5_ASAP7_75t_SL g12296 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[14]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[14]),
    .Y(n_957));
 AOI22xp5_ASAP7_75t_SL g12297 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[15]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[15]),
    .Y(n_956));
 AOI22xp5_ASAP7_75t_SL g12298 (.A1(n_22),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[16]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data1[16]),
    .Y(n_955));
 AOI22xp5_ASAP7_75t_SL g12299 (.A1(mac2accu_data1[1]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[1]),
    .Y(n_954));
 OAI21xp33_ASAP7_75t_SL g123 (.A1(n_13571),
    .A2(n_5427),
    .B(n_5431),
    .Y(n_5432));
 AOI22xp5_ASAP7_75t_SL g12300 (.A1(mac2accu_data1[4]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[4]),
    .Y(n_953));
 AOI22xp5_ASAP7_75t_SL g12301 (.A1(mac2accu_data1[7]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[7]),
    .Y(n_952));
 AOI22xp5_ASAP7_75t_SL g12302 (.A1(mac2accu_data1[10]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[10]),
    .Y(n_951));
 AOI22xp5_ASAP7_75t_SL g12303 (.A1(mac2accu_data1[13]),
    .A2(n_14),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[13]),
    .Y(n_950));
 AOI22xp5_ASAP7_75t_SL g12304 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[0]),
    .Y(n_949));
 AOI22xp5_ASAP7_75t_SL g12305 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[1]),
    .Y(n_948));
 AOI22xp5_ASAP7_75t_SL g12306 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[3]),
    .Y(n_947));
 AOI22xp5_ASAP7_75t_SL g12307 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[5]),
    .Y(n_946));
 AOI22xp5_ASAP7_75t_SL g12308 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[7]),
    .Y(n_945));
 AOI22xp5_ASAP7_75t_SL g12309 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[10]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[10]),
    .Y(n_944));
 AOI22xp5_ASAP7_75t_SL g12310 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[11]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[11]),
    .Y(n_943));
 AOI22xp5_ASAP7_75t_SL g12311 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[13]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[13]),
    .Y(n_942));
 AOI22xp5_ASAP7_75t_SL g12312 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[15]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[15]),
    .Y(n_941));
 AOI22xp5_ASAP7_75t_SL g12313 (.A1(n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[18]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data2[18]),
    .Y(n_940));
 AOI22xp5_ASAP7_75t_SL g12314 (.A1(mac2accu_data2[0]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[0]),
    .Y(n_939));
 AOI22xp5_ASAP7_75t_SL g12315 (.A1(mac2accu_data2[1]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[1]),
    .Y(n_938));
 AOI22xp5_ASAP7_75t_SL g12316 (.A1(mac2accu_data2[2]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[2]),
    .Y(n_937));
 AOI22xp5_ASAP7_75t_SL g12317 (.A1(mac2accu_data2[3]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[3]),
    .Y(n_936));
 AOI22xp5_ASAP7_75t_SL g12318 (.A1(mac2accu_data2[4]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[4]),
    .Y(n_935));
 AOI22xp5_ASAP7_75t_SL g12319 (.A1(mac2accu_data2[6]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[6]),
    .Y(n_934));
 AOI22xp5_ASAP7_75t_SL g12320 (.A1(mac2accu_data2[7]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[7]),
    .Y(n_933));
 AOI22xp5_ASAP7_75t_SL g12321 (.A1(mac2accu_data2[8]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[8]),
    .Y(n_932));
 AOI22xp5_ASAP7_75t_SL g12322 (.A1(mac2accu_data2[10]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[10]),
    .Y(n_931));
 AOI22xp5_ASAP7_75t_SL g12323 (.A1(mac2accu_data2[12]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[12]),
    .Y(n_930));
 AOI22xp5_ASAP7_75t_SL g12324 (.A1(mac2accu_data2[13]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[13]),
    .Y(n_929));
 AOI22xp5_ASAP7_75t_SL g12325 (.A1(mac2accu_data2[14]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[14]),
    .Y(n_928));
 AOI22xp5_ASAP7_75t_SL g12326 (.A1(mac2accu_data2[15]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[15]),
    .Y(n_927));
 AOI22xp5_ASAP7_75t_SL g12327 (.A1(mac2accu_data2[16]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[16]),
    .Y(n_926));
 AOI22xp5_ASAP7_75t_SL g12328 (.A1(mac2accu_data2[17]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[17]),
    .Y(n_925));
 AOI22xp5_ASAP7_75t_SL g12329 (.A1(mac2accu_data2[18]),
    .A2(n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[18]),
    .Y(n_924));
 AOI22xp5_ASAP7_75t_SL g12330 (.A1(mac2accu_data0[6]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[6]),
    .Y(n_923));
 AOI22xp5_ASAP7_75t_SL g12331 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[4]),
    .Y(n_922));
 AOI22xp5_ASAP7_75t_SL g12332 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[6]),
    .Y(n_921));
 AOI22xp5_ASAP7_75t_SL g12333 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[8]),
    .Y(n_920));
 AOI22xp5_ASAP7_75t_SL g12334 (.A1(mac2accu_data0[5]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[5]),
    .Y(n_919));
 AOI22xp5_ASAP7_75t_SL g12335 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[10]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[10]),
    .Y(n_918));
 AOI22xp5_ASAP7_75t_SL g12336 (.A1(mac2accu_data0[1]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[1]),
    .Y(n_917));
 AOI22xp5_ASAP7_75t_SL g12337 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[12]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[12]),
    .Y(n_916));
 AOI22xp5_ASAP7_75t_SL g12338 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[16]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[16]),
    .Y(n_915));
 AOI22xp5_ASAP7_75t_SL g12339 (.A1(n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[18]),
    .B1(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .B2(u_NV_NVDLA_cmac_u_core_out_data3[18]),
    .Y(n_914));
 AOI22xp5_ASAP7_75t_SL g12340 (.A1(mac2accu_data0[4]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[4]),
    .Y(n_913));
 AOI22xp5_ASAP7_75t_SL g12341 (.A1(mac2accu_data3[2]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[2]),
    .Y(n_912));
 AOI22xp5_ASAP7_75t_SL g12342 (.A1(mac2accu_data3[5]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[5]),
    .Y(n_911));
 AOI22xp5_ASAP7_75t_SL g12343 (.A1(mac2accu_data3[8]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[8]),
    .Y(n_910));
 AOI22xp5_ASAP7_75t_SL g12344 (.A1(mac2accu_data0[3]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[3]),
    .Y(n_909));
 AOI22xp5_ASAP7_75t_SL g12345 (.A1(mac2accu_data3[11]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[11]),
    .Y(n_908));
 AOI22xp5_ASAP7_75t_SL g12346 (.A1(mac2accu_data3[14]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[14]),
    .Y(n_907));
 AOI22xp5_ASAP7_75t_SL g12347 (.A1(mac2accu_data3[17]),
    .A2(n_17),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[17]),
    .Y(n_906));
 AOI22xp5_ASAP7_75t_SL g12348 (.A1(mac2accu_data0[2]),
    .A2(n_6),
    .B1(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[2]),
    .Y(n_905));
 AOI22xp5_ASAP7_75t_SL g12349 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[0]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[0]),
    .Y(n_904));
 AOI22xp5_ASAP7_75t_SL g12350 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[1]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[1]),
    .Y(n_903));
 AOI22xp5_ASAP7_75t_SL g12351 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[4]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[4]),
    .Y(n_902));
 AOI22xp5_ASAP7_75t_SL g12352 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[0]),
    .Y(n_901));
 AOI22xp5_ASAP7_75t_SL g12353 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[1]),
    .Y(n_900));
 AOI22xp5_ASAP7_75t_SL g12354 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[2]),
    .Y(n_899));
 AOI22xp5_ASAP7_75t_SL g12355 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[3]),
    .Y(n_898));
 AOI22xp5_ASAP7_75t_SL g12356 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[5]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_stripe_st),
    .Y(n_897));
 AOI22xp5_ASAP7_75t_SL g12357 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[4]),
    .Y(n_896));
 AOI22xp5_ASAP7_75t_SL g12358 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[5]),
    .Y(n_895));
 AOI22xp5_ASAP7_75t_SL g12359 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[6]),
    .Y(n_894));
 AOI22xp5_ASAP7_75t_SL g12360 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_mask[7]),
    .Y(n_893));
 AOI22xp5_ASAP7_75t_SL g12361 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[2]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[2]),
    .Y(n_892));
 AOI22xp5_ASAP7_75t_SL g12362 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[7]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[7]),
    .Y(n_891));
 AOI22xp5_ASAP7_75t_SL g12363 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[8]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[8]),
    .Y(n_890));
 AOI22xp5_ASAP7_75t_SL g12364 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[3]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[3]),
    .Y(n_889));
 AOI22xp5_ASAP7_75t_SL g12365 (.A1(n_3),
    .A2(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[6]),
    .B1(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B2(u_NV_NVDLA_cmac_u_core_in_dat_stripe_end),
    .Y(n_888));
 AOI22xp33_ASAP7_75t_SL g12366 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_887));
 AOI22xp33_ASAP7_75t_SL g12367 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_886));
 AOI22xp33_ASAP7_75t_SL g12368 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_885));
 AOI22xp33_ASAP7_75t_SL g12369 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_884));
 AOI22xp33_ASAP7_75t_SL g12370 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_883));
 AOI22xp33_ASAP7_75t_SL g12371 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_882));
 AOI22xp33_ASAP7_75t_SL g12372 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_881));
 AOI22xp33_ASAP7_75t_SL g12373 (.A1(n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_880));
 AOI22xp33_ASAP7_75t_SL g12374 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_879));
 AOI22xp33_ASAP7_75t_SL g12375 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_878));
 AOI22xp33_ASAP7_75t_SL g12376 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_877));
 AOI22xp33_ASAP7_75t_SL g12377 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_876));
 AOI22xp33_ASAP7_75t_SL g12378 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_875));
 AOI22xp33_ASAP7_75t_SL g12379 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_874));
 AOI21xp5_ASAP7_75t_SL g1238 (.A1(n_24203),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_445),
    .B(n_25449),
    .Y(n_5941));
 AOI22xp33_ASAP7_75t_SL g12380 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_873));
 AOI22xp33_ASAP7_75t_SL g12381 (.A1(n_314),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_872));
 AOI22xp33_ASAP7_75t_SL g12382 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_871));
 AOI22xp33_ASAP7_75t_SL g12383 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_870));
 AOI22xp33_ASAP7_75t_SL g12384 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_869));
 AOI22xp33_ASAP7_75t_SL g12385 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_868));
 AOI22xp33_ASAP7_75t_SL g12386 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_867));
 AOI22xp33_ASAP7_75t_SL g12387 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_866));
 AOI22xp33_ASAP7_75t_SL g12388 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_865));
 AOI22xp33_ASAP7_75t_SL g12389 (.A1(n_313),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_864));
 NAND2xp5_ASAP7_75t_SL g1239 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_445),
    .B(n_24203),
    .Y(n_5944));
 AOI22xp33_ASAP7_75t_SL g12390 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_863));
 AOI22xp33_ASAP7_75t_SL g12391 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_862));
 AOI22xp33_ASAP7_75t_SL g12392 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_861));
 AOI22xp33_ASAP7_75t_SL g12393 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_860));
 AOI22xp33_ASAP7_75t_SL g12394 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_859));
 AOI22xp33_ASAP7_75t_SL g12395 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_858));
 AOI22xp33_ASAP7_75t_SL g12396 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_857));
 AOI22xp33_ASAP7_75t_SL g12397 (.A1(n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .B1(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B2(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_856));
 AOI22xp5_ASAP7_75t_SL g12398 (.A1(n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[3]),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[3]),
    .Y(n_855));
 INVx1_ASAP7_75t_SL g12399 (.A(n_853),
    .Y(n_852));
 AOI21xp5_ASAP7_75t_SL g124 (.A1(n_13571),
    .A2(n_5429),
    .B(n_5430),
    .Y(n_5431));
 AOI31xp33_ASAP7_75t_SL g1240 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .A2(n_20633),
    .A3(n_5379),
    .B(n_5935),
    .Y(n_5936));
 INVx1_ASAP7_75t_SL g12400 (.A(n_851),
    .Y(n_850));
 INVx1_ASAP7_75t_SL g12401 (.A(n_848),
    .Y(n_847));
 INVx1_ASAP7_75t_SL g12402 (.A(n_846),
    .Y(n_845));
 INVx1_ASAP7_75t_SL g12403 (.A(n_844),
    .Y(n_843));
 INVx1_ASAP7_75t_SL g12404 (.A(n_842),
    .Y(n_841));
 INVx1_ASAP7_75t_SL g12405 (.A(n_840),
    .Y(n_839));
 INVx1_ASAP7_75t_SL g12406 (.A(n_837),
    .Y(n_836));
 INVx1_ASAP7_75t_SL g12407 (.A(n_835),
    .Y(n_834));
 INVx1_ASAP7_75t_SL g12408 (.A(n_832),
    .Y(n_831));
 INVx1_ASAP7_75t_SL g12409 (.A(n_830),
    .Y(n_829));
 AOI21xp33_ASAP7_75t_SL g1241 (.A1(n_20633),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .B(n_5380),
    .Y(n_5943));
 INVx1_ASAP7_75t_SL g12410 (.A(n_827),
    .Y(n_826));
 INVx1_ASAP7_75t_SL g12411 (.A(n_824),
    .Y(n_823));
 INVx1_ASAP7_75t_SL g12412 (.A(n_822),
    .Y(n_821));
 INVx1_ASAP7_75t_SL g12413 (.A(n_820),
    .Y(n_819));
 INVx1_ASAP7_75t_SL g12414 (.A(n_17240),
    .Y(n_817));
 NAND2xp5_ASAP7_75t_SL g12415 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_816));
 NAND2xp5_ASAP7_75t_SL g12416 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_815));
 NAND2xp5_ASAP7_75t_SL g12417 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_814));
 NAND2xp5_ASAP7_75t_SL g12418 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_813));
 NAND2xp5_ASAP7_75t_SL g12419 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_812));
 NAND2xp5_ASAP7_75t_SL g12420 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_811));
 NAND2xp5_ASAP7_75t_SL g12421 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_810));
 NAND2xp5_ASAP7_75t_SL g12422 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_809));
 NAND2xp5_ASAP7_75t_SL g12423 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_808));
 NAND2xp5_ASAP7_75t_SL g12424 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_807));
 NAND2xp5_ASAP7_75t_SL g12425 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_806));
 NAND2xp5_ASAP7_75t_SL g12426 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_805));
 NAND2xp5_ASAP7_75t_SL g12427 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_804));
 NAND2xp5_ASAP7_75t_SL g12428 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_803));
 NAND2xp5_ASAP7_75t_SL g12429 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_802));
 NAND2xp5_ASAP7_75t_SL g12430 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_801));
 NAND2xp5_ASAP7_75t_SL g12431 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_800));
 NAND2xp5_ASAP7_75t_SL g12432 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_799));
 NAND2xp5_ASAP7_75t_SL g12433 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_798));
 NAND2xp5_ASAP7_75t_SL g12434 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_797));
 NAND2xp5_ASAP7_75t_SL g12435 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_796));
 NAND2xp5_ASAP7_75t_SL g12436 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_795));
 NAND2xp5_ASAP7_75t_SL g12437 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_794));
 NAND2xp5_ASAP7_75t_SL g12438 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_793));
 NAND2xp5_ASAP7_75t_SL g12439 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_792));
 NAND2xp5_ASAP7_75t_SL g12440 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_791));
 NAND2xp5_ASAP7_75t_SL g12441 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_790));
 NAND2xp5_ASAP7_75t_SL g12442 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_789));
 NAND2xp5_ASAP7_75t_SL g12443 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_788));
 NAND2xp5_ASAP7_75t_SL g12444 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_787));
 NAND2xp5_ASAP7_75t_SL g12445 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_786));
 NAND2xp5_ASAP7_75t_SL g12446 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_785));
 NAND2xp5_ASAP7_75t_SL g12447 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_784));
 NAND2xp5_ASAP7_75t_SL g12448 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_783));
 NAND2xp5_ASAP7_75t_SL g12449 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_782));
 NAND2xp5_ASAP7_75t_SL g12450 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_781));
 NAND2xp5_ASAP7_75t_SL g12451 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_780));
 NAND2xp5_ASAP7_75t_SL g12452 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_779));
 NAND2xp5_ASAP7_75t_SL g12453 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_778));
 NAND2xp5_ASAP7_75t_SL g12454 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_777));
 NAND2xp5_ASAP7_75t_SL g12455 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_776));
 NAND2xp5_ASAP7_75t_SL g12456 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_775));
 NAND2xp5_ASAP7_75t_SL g12457 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_774));
 NAND2xp5_ASAP7_75t_SL g12458 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_773));
 NAND2xp5_ASAP7_75t_SL g12459 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_772));
 NAND2xp5_ASAP7_75t_SL g12460 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_771));
 NAND2xp5_ASAP7_75t_SL g12461 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_770));
 NAND2xp5_ASAP7_75t_SL g12462 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_769));
 NAND2xp5_ASAP7_75t_SL g12463 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_768));
 NAND2xp5_ASAP7_75t_SL g12464 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_767));
 NAND2xp5_ASAP7_75t_SL g12465 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_766));
 NAND2xp5_ASAP7_75t_SL g12466 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_765));
 NAND2xp5_ASAP7_75t_SL g12467 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_764));
 NAND2xp5_ASAP7_75t_SL g12468 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_763));
 NAND2xp5_ASAP7_75t_SL g12469 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_762));
 INVxp67_ASAP7_75t_SL g1247 (.A(n_5383),
    .Y(n_5935));
 NAND2xp5_ASAP7_75t_SL g12470 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_761));
 NAND2xp5_ASAP7_75t_SL g12471 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_760));
 NAND2xp5_ASAP7_75t_SL g12472 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_759));
 NAND2xp5_ASAP7_75t_SL g12473 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_758));
 NAND2xp5_ASAP7_75t_SL g12474 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_757));
 NAND2xp5_ASAP7_75t_SL g12475 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_756));
 NAND2xp5_ASAP7_75t_SL g12476 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_755));
 NAND2xp5_ASAP7_75t_SL g12477 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_754));
 NAND2xp5_ASAP7_75t_SL g12478 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_753));
 NAND2xp5_ASAP7_75t_SL g12479 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_752));
 NAND2xp5_ASAP7_75t_SL g12480 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_751));
 NAND2xp5_ASAP7_75t_SL g12481 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_750));
 NAND2xp5_ASAP7_75t_SL g12482 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_749));
 NAND2xp5_ASAP7_75t_SL g12483 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_748));
 NAND2xp5_ASAP7_75t_SL g12484 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_747));
 NAND2xp5_ASAP7_75t_SL g12485 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_746));
 NAND2xp5_ASAP7_75t_SL g12486 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_745));
 NAND2xp5_ASAP7_75t_SL g12487 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_744));
 NAND2xp5_ASAP7_75t_SL g12488 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_743));
 NAND2xp5_ASAP7_75t_SL g12489 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_742));
 NAND2xp5_ASAP7_75t_SL g12490 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_741));
 NAND2xp5_ASAP7_75t_SL g12491 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_740));
 NAND2xp5_ASAP7_75t_SL g12492 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_739));
 NAND2xp5_ASAP7_75t_SL g12493 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_738));
 NAND2xp5_ASAP7_75t_SL g12494 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .Y(n_737));
 NAND2xp5_ASAP7_75t_SL g12495 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_736));
 NAND2xp5_ASAP7_75t_SL g12496 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_735));
 NAND2xp5_ASAP7_75t_SL g12497 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_734));
 NAND2xp33_ASAP7_75t_SL g12498 (.A(u_NV_NVDLA_cmac_dp2reg_done),
    .B(n_334),
    .Y(n_733));
 NAND2xp5_ASAP7_75t_SL g12499 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_732));
 NAND2xp33_ASAP7_75t_SL g125 (.A(n_5426),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_449),
    .Y(n_5427));
 NAND2xp5_ASAP7_75t_SL g12500 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_731));
 NAND2xp5_ASAP7_75t_SL g12501 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .Y(n_730));
 NAND2xp5_ASAP7_75t_SL g12502 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_729));
 NAND2xp5_ASAP7_75t_SL g12503 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_728));
 NAND2xp5_ASAP7_75t_SL g12504 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_727));
 NAND2xp5_ASAP7_75t_SL g12505 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_726));
 NAND2xp5_ASAP7_75t_SL g12506 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_725));
 NAND2xp5_ASAP7_75t_SL g12507 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_724));
 NAND2xp5_ASAP7_75t_SL g12508 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_723));
 NAND2xp5_ASAP7_75t_SL g12509 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_722));
 NAND2xp5_ASAP7_75t_SL g12510 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_721));
 NAND2xp5_ASAP7_75t_SL g12511 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_720));
 NAND2xp5_ASAP7_75t_SL g12512 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_719));
 NAND2xp5_ASAP7_75t_SL g12513 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_718));
 NAND2xp5_ASAP7_75t_SL g12514 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_717));
 NAND2xp5_ASAP7_75t_SL g12515 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_716));
 NAND2xp5_ASAP7_75t_SL g12516 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_715));
 NAND2xp5_ASAP7_75t_SL g12517 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_714));
 NAND2xp5_ASAP7_75t_SL g12518 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_713));
 NAND2xp5_ASAP7_75t_SL g12519 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .Y(n_712));
 NAND2xp5_ASAP7_75t_SL g12520 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_711));
 NAND2xp5_ASAP7_75t_SL g12521 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_710));
 NAND2xp5_ASAP7_75t_SL g12522 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_709));
 NAND2xp5_ASAP7_75t_SL g12523 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .Y(n_708));
 NAND2xp5_ASAP7_75t_SL g12524 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_707));
 NAND2xp5_ASAP7_75t_SL g12525 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_706));
 NAND2xp5_ASAP7_75t_SL g12526 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_705));
 NAND2xp5_ASAP7_75t_SL g12527 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_704));
 NAND2xp5_ASAP7_75t_SL g12528 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_703));
 NAND2xp5_ASAP7_75t_SL g12529 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_702));
 NAND2xp5_ASAP7_75t_SL g12530 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_701));
 NAND2xp5_ASAP7_75t_SL g12531 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_700));
 NAND2xp5_ASAP7_75t_SL g12532 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_699));
 NAND2xp5_ASAP7_75t_SL g12533 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_698));
 NAND2xp5_ASAP7_75t_SL g12534 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_697));
 NAND2xp5_ASAP7_75t_SL g12535 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_696));
 NAND2xp5_ASAP7_75t_SL g12536 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_695));
 NAND2xp5_ASAP7_75t_SL g12537 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_694));
 NAND2xp5_ASAP7_75t_SL g12538 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_693));
 NAND2xp5_ASAP7_75t_SL g12539 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_692));
 NAND2xp5_ASAP7_75t_SL g12540 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_691));
 NAND2xp5_ASAP7_75t_SL g12541 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_690));
 NAND2xp5_ASAP7_75t_SL g12542 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_689));
 NAND2xp5_ASAP7_75t_SL g12543 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_688));
 NAND2xp5_ASAP7_75t_SL g12545 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_686));
 NAND2xp5_ASAP7_75t_SL g12546 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_685));
 NAND2xp5_ASAP7_75t_SL g12547 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_684));
 NAND2xp5_ASAP7_75t_SL g12548 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_683));
 NAND2xp5_ASAP7_75t_SL g12549 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_682));
 NAND2xp5_ASAP7_75t_SL g12550 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_681));
 NAND2xp5_ASAP7_75t_SL g12551 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_680));
 NAND2xp5_ASAP7_75t_SL g12552 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_679));
 NAND2xp5_ASAP7_75t_SL g12553 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_678));
 NAND2xp5_ASAP7_75t_SL g12554 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_677));
 NAND2xp5_ASAP7_75t_SL g12555 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_676));
 NAND2xp5_ASAP7_75t_SL g12556 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_675));
 NAND2xp5_ASAP7_75t_SL g12557 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_674));
 NAND2xp5_ASAP7_75t_SL g12558 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_673));
 NOR2xp33_ASAP7_75t_SL g12559 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_actv_stripe_end),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_st_3519),
    .Y(n_854));
 NAND2xp5_ASAP7_75t_SL g12560 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[2]),
    .Y(n_853));
 NAND2xp5_ASAP7_75t_SL g12561 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[1]),
    .Y(n_851));
 NAND2xp5_ASAP7_75t_SL g12562 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[5]),
    .Y(n_849));
 NAND2xp5_ASAP7_75t_SL g12563 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[5]),
    .Y(n_848));
 NAND2xp5_ASAP7_75t_SL g12564 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[0]),
    .Y(n_846));
 NAND2xp5_ASAP7_75t_SL g12565 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[7]),
    .Y(n_844));
 NAND2xp5_ASAP7_75t_SL g12566 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[3]),
    .Y(n_842));
 NAND2xp5_ASAP7_75t_SL g12567 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[6]),
    .Y(n_840));
 NAND2xp5_ASAP7_75t_SL g12568 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[4]),
    .Y(n_838));
 NAND2xp5_ASAP7_75t_SL g12569 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[4]),
    .Y(n_837));
 A2O1A1O1Ixp25_ASAP7_75t_SL g1257 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_268),
    .A2(n_11586),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_270),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_197),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_191),
    .Y(n_11590));
 NAND2xp5_ASAP7_75t_SL g12570 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[7]),
    .Y(n_835));
 NAND2xp5_ASAP7_75t_SL g12571 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[1]),
    .Y(n_833));
 NAND2xp5_ASAP7_75t_SL g12572 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[2]),
    .Y(n_832));
 NAND2xp5_ASAP7_75t_SL g12573 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[1]),
    .Y(n_830));
 NAND2xp5_ASAP7_75t_SL g12574 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[7]),
    .Y(n_828));
 NAND2xp5_ASAP7_75t_SL g12575 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[0]),
    .Y(n_827));
 NOR2xp33_ASAP7_75t_SL g12577 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .Y(n_824));
 NOR2xp33_ASAP7_75t_L g12578 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .Y(n_822));
 OR2x2_ASAP7_75t_SL g12579 (.A(n_46),
    .B(n_448),
    .Y(n_820));
 OAI22xp33_ASAP7_75t_SL g1258 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_264),
    .A2(n_11586),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_265),
    .B2(n_11583),
    .Y(n_11587));
 INVx1_ASAP7_75t_SL g12582 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_st_3519),
    .Y(n_46));
 INVx1_ASAP7_75t_SL g12585 (.A(n_660),
    .Y(n_659));
 INVx1_ASAP7_75t_SL g12586 (.A(n_658),
    .Y(n_657));
 INVx1_ASAP7_75t_SL g12587 (.A(n_656),
    .Y(n_655));
 INVx1_ASAP7_75t_SL g12588 (.A(n_654),
    .Y(n_653));
 INVx1_ASAP7_75t_SL g12589 (.A(n_652),
    .Y(n_651));
 OAI21x1_ASAP7_75t_SL g1259 (.A1(n_11568),
    .A2(n_11583),
    .B(n_11584),
    .Y(n_11585));
 INVx1_ASAP7_75t_SL g12590 (.A(n_650),
    .Y(n_649));
 INVx1_ASAP7_75t_SL g12591 (.A(n_648),
    .Y(n_647));
 INVx1_ASAP7_75t_SL g12592 (.A(n_646),
    .Y(n_645));
 INVx1_ASAP7_75t_SL g12593 (.A(n_644),
    .Y(n_643));
 INVx1_ASAP7_75t_SL g12594 (.A(n_642),
    .Y(n_641));
 INVx1_ASAP7_75t_SL g12595 (.A(n_640),
    .Y(n_639));
 INVx1_ASAP7_75t_SL g12596 (.A(n_638),
    .Y(n_637));
 INVx1_ASAP7_75t_SL g12597 (.A(n_636),
    .Y(n_635));
 INVx1_ASAP7_75t_SL g12598 (.A(n_634),
    .Y(n_633));
 INVx1_ASAP7_75t_SL g12599 (.A(n_632),
    .Y(n_631));
 NOR2xp33_ASAP7_75t_SL g126 (.A(n_5428),
    .B(n_17936),
    .Y(n_5430));
 INVx1_ASAP7_75t_SL g12600 (.A(n_630),
    .Y(n_629));
 INVx1_ASAP7_75t_SL g12601 (.A(n_628),
    .Y(n_627));
 INVx1_ASAP7_75t_SL g12602 (.A(n_625),
    .Y(n_624));
 INVx1_ASAP7_75t_SL g12603 (.A(n_623),
    .Y(n_622));
 INVx1_ASAP7_75t_SL g12604 (.A(n_620),
    .Y(n_619));
 INVx1_ASAP7_75t_SL g12605 (.A(n_618),
    .Y(n_617));
 INVx1_ASAP7_75t_SL g12606 (.A(n_616),
    .Y(n_615));
 INVx1_ASAP7_75t_SL g12607 (.A(n_614),
    .Y(n_613));
 INVx1_ASAP7_75t_SL g12608 (.A(n_612),
    .Y(n_611));
 INVx1_ASAP7_75t_SL g12609 (.A(n_610),
    .Y(n_609));
 OA21x2_ASAP7_75t_SL g1261 (.A1(n_11570),
    .A2(n_11574),
    .B(n_11582),
    .Y(n_11583));
 INVx1_ASAP7_75t_SL g12610 (.A(n_608),
    .Y(n_607));
 INVx1_ASAP7_75t_SL g12611 (.A(n_606),
    .Y(n_605));
 INVx1_ASAP7_75t_SL g12612 (.A(n_604),
    .Y(n_603));
 INVx1_ASAP7_75t_SL g12613 (.A(n_602),
    .Y(n_601));
 INVx1_ASAP7_75t_SL g12614 (.A(n_600),
    .Y(n_599));
 INVx1_ASAP7_75t_SL g12615 (.A(n_598),
    .Y(n_597));
 INVx1_ASAP7_75t_SL g12616 (.A(n_596),
    .Y(n_595));
 INVx1_ASAP7_75t_SL g12617 (.A(n_594),
    .Y(n_593));
 INVx1_ASAP7_75t_SL g12618 (.A(n_592),
    .Y(n_591));
 INVx1_ASAP7_75t_SL g12619 (.A(n_590),
    .Y(n_589));
 INVx1_ASAP7_75t_SL g12620 (.A(n_588),
    .Y(n_587));
 INVx1_ASAP7_75t_SL g12621 (.A(n_586),
    .Y(n_585));
 INVx1_ASAP7_75t_SL g12622 (.A(n_584),
    .Y(n_583));
 INVx1_ASAP7_75t_SL g12623 (.A(n_582),
    .Y(n_581));
 INVx1_ASAP7_75t_SL g12624 (.A(n_580),
    .Y(n_579));
 NAND2xp5_ASAP7_75t_SL g12625 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_578));
 NAND2xp5_ASAP7_75t_SL g12626 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_577));
 NOR2xp33_ASAP7_75t_SL g12627 (.A(u_NV_NVDLA_cmac_u_reg_dp2reg_consumer),
    .B(n_336),
    .Y(n_576));
 NAND2xp5_ASAP7_75t_SL g12628 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_575));
 NAND2xp5_ASAP7_75t_SL g12629 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_574));
 OAI21xp5_ASAP7_75t_SL g1263 (.A1(n_8159),
    .A2(n_11570),
    .B(n_18717),
    .Y(n_11592));
 NOR2xp33_ASAP7_75t_SL g12630 (.A(u_NV_NVDLA_cmac_u_reg_dp2reg_consumer),
    .B(n_338),
    .Y(n_573));
 NAND2xp5_ASAP7_75t_SL g12631 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_572));
 NAND2xp5_ASAP7_75t_SL g12632 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_571));
 NAND2xp5_ASAP7_75t_SL g12633 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_570));
 NAND2xp5_ASAP7_75t_SL g12634 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_569));
 NAND2xp5_ASAP7_75t_SL g12635 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_568));
 NAND2xp5_ASAP7_75t_SL g12636 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_567));
 NAND2xp5_ASAP7_75t_SL g12637 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_566));
 NAND2xp5_ASAP7_75t_SL g12638 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_565));
 NAND2xp5_ASAP7_75t_SL g12639 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_564));
 AOI21xp5_ASAP7_75t_SL g1264 (.A1(n_11576),
    .A2(n_11579),
    .B(n_11581),
    .Y(n_11582));
 NAND2xp5_ASAP7_75t_SL g12640 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_563));
 NAND2xp5_ASAP7_75t_SL g12641 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_562));
 NAND2xp5_ASAP7_75t_SL g12642 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_561));
 NAND2xp5_ASAP7_75t_SL g12643 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_560));
 NAND2xp5_ASAP7_75t_SL g12644 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_559));
 NAND2xp5_ASAP7_75t_SL g12645 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_558));
 NAND2xp5_ASAP7_75t_SL g12646 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_557));
 NAND2xp5_ASAP7_75t_SL g12647 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_556));
 NAND2xp5_ASAP7_75t_SL g12648 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_555));
 NAND2xp5_ASAP7_75t_SL g12649 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_554));
 AOI22xp5_ASAP7_75t_SL g1265 (.A1(n_24034),
    .A2(n_8161),
    .B1(n_11596),
    .B2(n_11579),
    .Y(n_11597));
 NAND2xp5_ASAP7_75t_SL g12650 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_553));
 NAND2xp5_ASAP7_75t_SL g12651 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_552));
 NAND2xp5_ASAP7_75t_SL g12652 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_551));
 NAND2xp5_ASAP7_75t_SL g12653 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_550));
 NAND2xp5_ASAP7_75t_SL g12654 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_549));
 NAND2xp5_ASAP7_75t_SL g12655 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_548));
 NAND2xp5_ASAP7_75t_SL g12656 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_547));
 NAND2xp5_ASAP7_75t_SL g12657 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_546));
 NAND2xp5_ASAP7_75t_SL g12658 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_545));
 NAND2xp5_ASAP7_75t_SL g12659 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_544));
 NAND2xp5_ASAP7_75t_SL g1266 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259),
    .B(n_11598),
    .Y(n_11599));
 NAND2xp5_ASAP7_75t_SL g12660 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_543));
 NAND2xp5_ASAP7_75t_SL g12661 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_542));
 NAND2xp5_ASAP7_75t_SL g12662 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .Y(n_541));
 NAND2xp5_ASAP7_75t_SL g12663 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_540));
 NAND2xp5_ASAP7_75t_SL g12664 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_539));
 NAND2xp5_ASAP7_75t_SL g12665 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_538));
 NAND2xp5_ASAP7_75t_SL g12666 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .Y(n_537));
 NAND2xp5_ASAP7_75t_SL g12667 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_536));
 NAND2xp5_ASAP7_75t_SL g12668 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_535));
 NAND2xp5_ASAP7_75t_SL g12669 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_534));
 NAND2xp5_ASAP7_75t_SL g1267 (.A(n_11573),
    .B(n_8161),
    .Y(n_11574));
 NAND2xp5_ASAP7_75t_SL g12670 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_533));
 NAND2xp5_ASAP7_75t_SL g12671 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_532));
 NAND2xp5_ASAP7_75t_SL g12672 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_531));
 NAND2xp5_ASAP7_75t_SL g12673 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_530));
 NAND2xp5_ASAP7_75t_SL g12674 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_529));
 NAND2xp5_ASAP7_75t_SL g12675 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_528));
 NAND2xp5_ASAP7_75t_SL g12676 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_527));
 NAND2xp5_ASAP7_75t_SL g12677 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_526));
 NAND2xp5_ASAP7_75t_SL g12678 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_525));
 NAND2xp5_ASAP7_75t_SL g12679 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_524));
 AO21x1_ASAP7_75t_SL g1268 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_276),
    .B(n_11580),
    .Y(n_11581));
 NAND2xp5_ASAP7_75t_SL g12680 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_523));
 NAND2xp5_ASAP7_75t_SL g12681 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_522));
 NAND2xp5_ASAP7_75t_SL g12682 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_521));
 NAND2xp5_ASAP7_75t_SL g12683 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_520));
 NAND2xp5_ASAP7_75t_SL g12684 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_519));
 NAND2xp5_ASAP7_75t_SL g12685 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_518));
 NAND2xp5_ASAP7_75t_SL g12686 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_517));
 NAND2xp5_ASAP7_75t_SL g12687 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_516));
 NAND2xp5_ASAP7_75t_SL g12688 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .Y(n_515));
 NOR2xp33_ASAP7_75t_SL g1269 (.A(n_11575),
    .B(n_4079),
    .Y(n_11576));
 NAND2xp5_ASAP7_75t_SL g12690 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .Y(n_513));
 NAND2xp5_ASAP7_75t_SL g12691 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .Y(n_512));
 NAND2xp5_ASAP7_75t_SL g12692 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_511));
 NAND2xp5_ASAP7_75t_SL g12693 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_510));
 NAND2xp5_ASAP7_75t_SL g12694 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_509));
 NAND2xp5_ASAP7_75t_SL g12695 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_508));
 NAND2xp5_ASAP7_75t_SL g12696 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .Y(n_507));
 NAND2xp5_ASAP7_75t_SL g12697 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .Y(n_506));
 NAND2xp5_ASAP7_75t_SL g12698 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_505));
 NAND2xp5_ASAP7_75t_SL g12699 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_504));
 NOR2xp33_ASAP7_75t_SL g127 (.A(n_5428),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_449),
    .Y(n_5429));
 NAND2xp5_ASAP7_75t_SL g12700 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_503));
 NAND2xp5_ASAP7_75t_SL g12701 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .Y(n_502));
 NAND2xp5_ASAP7_75t_SL g12702 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .Y(n_501));
 NAND2xp5_ASAP7_75t_SL g12703 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .Y(n_500));
 NAND2xp5_ASAP7_75t_SL g12704 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .Y(n_499));
 NAND2xp5_ASAP7_75t_SL g12705 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_498));
 NAND2xp5_ASAP7_75t_SL g12706 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .Y(n_497));
 NAND2xp5_ASAP7_75t_SL g12707 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_496));
 NAND2xp5_ASAP7_75t_SL g12708 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_495));
 NAND2xp5_ASAP7_75t_SL g12709 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .Y(n_494));
 HB1xp67_ASAP7_75t_SL g1271 (.A(n_24034),
    .Y(n_11593));
 NAND2xp5_ASAP7_75t_SL g12710 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .Y(n_493));
 NAND2xp5_ASAP7_75t_SL g12711 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_492));
 NAND2xp5_ASAP7_75t_SL g12712 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_491));
 NAND2xp5_ASAP7_75t_SL g12713 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .Y(n_490));
 NAND2xp5_ASAP7_75t_SL g12714 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_489));
 NAND2xp5_ASAP7_75t_SL g12715 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_488));
 NAND2xp5_ASAP7_75t_SL g12716 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_487));
 NAND2xp5_ASAP7_75t_SL g12717 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_486));
 NAND2xp5_ASAP7_75t_SL g12718 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_485));
 NAND2xp5_ASAP7_75t_SL g12719 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_484));
 NAND2xp5_ASAP7_75t_SL g12720 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .Y(n_483));
 NAND2xp5_ASAP7_75t_SL g12721 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_482));
 NAND2xp5_ASAP7_75t_SL g12722 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_481));
 NAND2xp5_ASAP7_75t_SL g12723 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_480));
 NAND2xp5_ASAP7_75t_SL g12724 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_479));
 NAND2xp5_ASAP7_75t_SL g12725 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .Y(n_478));
 NAND2xp5_ASAP7_75t_SL g12726 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_477));
 NAND2xp5_ASAP7_75t_SL g12727 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .Y(n_476));
 NAND2xp5_ASAP7_75t_SL g12728 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .Y(n_475));
 NAND2xp5_ASAP7_75t_SL g12729 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_474));
 INVx1_ASAP7_75t_SL g1273 (.A(n_24034),
    .Y(n_11570));
 NAND2xp5_ASAP7_75t_SL g12730 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_473));
 NAND2xp5_ASAP7_75t_SL g12731 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_472));
 NAND2xp5_ASAP7_75t_SL g12732 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .Y(n_471));
 NAND2xp5_ASAP7_75t_SL g12733 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .Y(n_470));
 NAND2xp5_ASAP7_75t_SL g12734 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .Y(n_469));
 NAND2xp5_ASAP7_75t_SL g12735 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_468));
 NAND2xp5_ASAP7_75t_SL g12736 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .Y(n_467));
 NAND2xp5_ASAP7_75t_SL g12737 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .Y(n_466));
 NAND2xp5_ASAP7_75t_SL g12738 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .Y(n_465));
 NAND2xp5_ASAP7_75t_SL g12739 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .Y(n_464));
 NAND2xp5_ASAP7_75t_SL g12740 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .Y(n_463));
 NOR2xp33_ASAP7_75t_SL g12742 (.A(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .B(u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en),
    .Y(n_670));
 NOR2xp33_ASAP7_75t_SL g12743 (.A(n_332),
    .B(u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en),
    .Y(n_669));
 NOR2xp33_ASAP7_75t_SL g12747 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .B(n_334),
    .Y(n_662));
 NAND2xp5_ASAP7_75t_SL g12748 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[0]),
    .Y(n_661));
 NAND2xp5_ASAP7_75t_SL g12749 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_660));
 NAND2xp5_ASAP7_75t_SL g1275 (.A(n_18717),
    .B(n_11578),
    .Y(n_11579));
 NAND2xp5_ASAP7_75t_SL g12750 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_658));
 NAND2xp5_ASAP7_75t_SL g12751 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[6]),
    .Y(n_656));
 NAND2xp5_ASAP7_75t_SL g12752 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_wt_mask[5]),
    .Y(n_654));
 NAND2xp5_ASAP7_75t_SL g12753 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_652));
 NAND2xp5_ASAP7_75t_SL g12754 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_650));
 NAND2xp5_ASAP7_75t_SL g12755 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_648));
 NAND2xp5_ASAP7_75t_SL g12756 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_646));
 NAND2xp5_ASAP7_75t_SL g12757 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_644));
 NAND2xp5_ASAP7_75t_SL g12758 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_642));
 NAND2xp5_ASAP7_75t_SL g12759 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_640));
 INVxp67_ASAP7_75t_SL g1276 (.A(n_11580),
    .Y(n_11598));
 NAND2xp5_ASAP7_75t_SL g12760 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_638));
 NAND2xp5_ASAP7_75t_SL g12761 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_636));
 NAND2xp5_ASAP7_75t_SL g12762 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_634));
 NAND2xp5_ASAP7_75t_SL g12763 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_632));
 NAND2xp5_ASAP7_75t_SL g12764 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_630));
 NAND2xp5_ASAP7_75t_SL g12765 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_628));
 NAND2xp5_ASAP7_75t_SL g12766 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[3]),
    .Y(n_626));
 NAND2xp5_ASAP7_75t_SL g12767 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .Y(n_625));
 NAND2xp5_ASAP7_75t_SL g12768 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_623));
 NAND2xp5_ASAP7_75t_SL g12769 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[2]),
    .Y(n_621));
 NOR2xp33_ASAP7_75t_SL g1277 (.A(n_26231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_249),
    .Y(n_11580));
 NAND2xp5_ASAP7_75t_SL g12770 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_620));
 NAND2xp5_ASAP7_75t_SL g12771 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[4]),
    .Y(n_618));
 NAND2xp5_ASAP7_75t_SL g12772 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_616));
 NAND2xp5_ASAP7_75t_SL g12773 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .Y(n_614));
 NAND2xp5_ASAP7_75t_SL g12774 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_612));
 NAND2xp5_ASAP7_75t_SL g12775 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_610));
 NAND2xp5_ASAP7_75t_SL g12776 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_608));
 NAND2xp5_ASAP7_75t_SL g12777 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .Y(n_606));
 NAND2xp5_ASAP7_75t_SL g12778 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_604));
 NAND2xp5_ASAP7_75t_SL g12779 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_in_dat_mask[3]),
    .Y(n_602));
 NOR2xp33_ASAP7_75t_SL g1278 (.A(n_11571),
    .B(n_4079),
    .Y(n_11573));
 NAND2xp5_ASAP7_75t_SL g12780 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_600));
 NAND2xp5_ASAP7_75t_SL g12781 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .Y(n_598));
 NAND2xp5_ASAP7_75t_SL g12782 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .Y(n_596));
 NAND2xp5_ASAP7_75t_SL g12783 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_594));
 NAND2xp5_ASAP7_75t_SL g12784 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .Y(n_592));
 NAND2xp5_ASAP7_75t_SL g12785 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .Y(n_590));
 NAND2xp5_ASAP7_75t_SL g12786 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .Y(n_588));
 NOR2xp33_ASAP7_75t_SL g12787 (.A(sc2mac_wt_pvld),
    .B(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1),
    .Y(n_586));
 NOR2xp33_ASAP7_75t_L g12788 (.A(sc2mac_dat_pvld),
    .B(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1),
    .Y(n_584));
 OR2x2_ASAP7_75t_SL g12789 (.A(n_46),
    .B(n_440),
    .Y(n_582));
 NAND2xp5_ASAP7_75t_SL g1279 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259),
    .B(n_11596),
    .Y(n_11575));
 OR2x2_ASAP7_75t_SL g12790 (.A(n_46),
    .B(n_441),
    .Y(n_580));
 INVxp67_ASAP7_75t_SL g12793 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[2]),
    .Y(n_460));
 INVxp67_ASAP7_75t_SL g12797 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[51]),
    .Y(n_457));
 INVx1_ASAP7_75t_SL g128 (.A(n_5426),
    .Y(n_5428));
 INVxp67_ASAP7_75t_SL g1280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_270),
    .Y(n_11584));
 INVxp67_ASAP7_75t_SL g12801 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[42]),
    .Y(n_453));
 INVxp67_ASAP7_75t_SL g12802 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[5]),
    .Y(n_452));
 INVxp67_ASAP7_75t_SL g12808 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[55]),
    .Y(n_449));
 INVx1_ASAP7_75t_SL g12810 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_pvld_3195),
    .Y(n_448));
 INVxp67_ASAP7_75t_SL g12814 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[22]),
    .Y(n_446));
 INVx1_ASAP7_75t_SL g12816 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_pvld_3196),
    .Y(n_445));
 INVxp67_ASAP7_75t_SL g12817 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[29]),
    .Y(n_444));
 INVxp67_ASAP7_75t_SL g12818 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[10]),
    .Y(n_443));
 INVxp67_ASAP7_75t_SL g1282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259),
    .Y(n_11571));
 INVx1_ASAP7_75t_SL g12820 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_pvld_3197),
    .Y(n_441));
 INVx1_ASAP7_75t_SL g12821 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_pvld_3198),
    .Y(n_440));
 INVxp67_ASAP7_75t_SL g12827 (.A(n_19396),
    .Y(n_434));
 INVxp67_ASAP7_75t_SL g12828 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[15]),
    .Y(n_433));
 INVxp67_ASAP7_75t_SL g12829 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[11]),
    .Y(n_432));
 INVxp67_ASAP7_75t_SL g12830 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[41]),
    .Y(n_431));
 INVxp67_ASAP7_75t_SL g12832 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[24]),
    .Y(n_429));
 INVxp67_ASAP7_75t_SL g12833 (.A(n_9273),
    .Y(n_428));
 INVxp67_ASAP7_75t_SL g12836 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[45]),
    .Y(n_425));
 INVxp67_ASAP7_75t_SL g12838 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[47]),
    .Y(n_423));
 INVxp67_ASAP7_75t_SL g12839 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[34]),
    .Y(n_422));
 INVxp67_ASAP7_75t_SL g12843 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[16]),
    .Y(n_418));
 INVxp67_ASAP7_75t_SL g12844 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[63]),
    .Y(n_417));
 INVxp67_ASAP7_75t_SL g12845 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[4]),
    .Y(n_416));
 INVxp67_ASAP7_75t_SL g12847 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[25]),
    .Y(n_414));
 INVxp67_ASAP7_75t_SL g12848 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[54]),
    .Y(n_413));
 INVx1_ASAP7_75t_SL g1285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_23),
    .Y(n_4079));
 INVxp67_ASAP7_75t_SL g12850 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[13]),
    .Y(n_411));
 INVxp67_ASAP7_75t_SL g12854 (.A(n_9154),
    .Y(n_407));
 INVxp67_ASAP7_75t_SL g12855 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[30]),
    .Y(n_406));
 INVxp67_ASAP7_75t_SL g12856 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[31]),
    .Y(n_405));
 INVxp67_ASAP7_75t_SL g12858 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[62]),
    .Y(n_403));
 INVxp67_ASAP7_75t_SL g12859 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[23]),
    .Y(n_402));
 INVx1_ASAP7_75t_SL g1286 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_267),
    .Y(n_11578));
 INVxp67_ASAP7_75t_SL g12861 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[28]),
    .Y(n_400));
 INVxp67_ASAP7_75t_SL g12863 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[59]),
    .Y(n_398));
 INVxp67_ASAP7_75t_SL g12864 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[9]),
    .Y(n_397));
 INVxp67_ASAP7_75t_SL g12866 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[35]),
    .Y(n_395));
 INVxp67_ASAP7_75t_SL g12870 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[0]),
    .Y(n_391));
 INVxp67_ASAP7_75t_SL g12873 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[58]),
    .Y(n_388));
 INVxp67_ASAP7_75t_SL g12876 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[43]),
    .Y(n_385));
 INVxp67_ASAP7_75t_SL g12879 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[12]),
    .Y(n_382));
 INVxp67_ASAP7_75t_SL g12880 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[27]),
    .Y(n_381));
 INVxp67_ASAP7_75t_SL g12885 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[57]),
    .Y(n_376));
 INVxp67_ASAP7_75t_SL g12887 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[14]),
    .Y(n_374));
 INVxp67_ASAP7_75t_SL g12888 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[39]),
    .Y(n_373));
 INVxp67_ASAP7_75t_SL g12889 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[32]),
    .Y(n_372));
 INVxp67_ASAP7_75t_SL g12891 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[26]),
    .Y(n_370));
 INVxp67_ASAP7_75t_SL g12893 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[20]),
    .Y(n_368));
 INVxp67_ASAP7_75t_SL g12895 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[44]),
    .Y(n_366));
 INVxp67_ASAP7_75t_SL g12896 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[61]),
    .Y(n_365));
 INVxp67_ASAP7_75t_SL g12897 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[6]),
    .Y(n_364));
 NAND2xp5_ASAP7_75t_SL g129 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[15]),
    .B(n_17882),
    .Y(n_5504));
 INVxp67_ASAP7_75t_SL g12901 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[18]),
    .Y(n_360));
 INVxp67_ASAP7_75t_SL g12902 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[40]),
    .Y(n_359));
 INVxp67_ASAP7_75t_SL g12903 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[8]),
    .Y(n_358));
 INVxp67_ASAP7_75t_SL g12906 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[56]),
    .Y(n_355));
 INVxp67_ASAP7_75t_SL g12907 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[46]),
    .Y(n_354));
 INVxp67_ASAP7_75t_SL g12908 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[38]),
    .Y(n_353));
 INVxp67_ASAP7_75t_SL g12910 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[60]),
    .Y(n_351));
 INVxp67_ASAP7_75t_SL g12913 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[37]),
    .Y(n_348));
 INVxp67_ASAP7_75t_SL g12914 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[53]),
    .Y(n_347));
 INVxp67_ASAP7_75t_SL g12915 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[36]),
    .Y(n_346));
 INVxp67_ASAP7_75t_SL g12917 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[49]),
    .Y(n_344));
 INVxp67_ASAP7_75t_SL g12918 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[52]),
    .Y(n_343));
 INVxp67_ASAP7_75t_SL g12920 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[48]),
    .Y(n_341));
 INVxp67_ASAP7_75t_SL g12922 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[7]),
    .Y(n_339));
 INVx1_ASAP7_75t_SL g12925 (.A(u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en),
    .Y(n_338));
 INVx1_ASAP7_75t_SL g12926 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .Y(n_337));
 INVxp67_ASAP7_75t_SL g12927 (.A(u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en),
    .Y(n_336));
 INVx1_ASAP7_75t_SL g12933 (.A(u_NV_NVDLA_cmac_u_reg_dp2reg_consumer),
    .Y(n_334));
 INVx1_ASAP7_75t_SL g12934 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .Y(n_333));
 INVx1_ASAP7_75t_SL g12935 (.A(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .Y(n_332));
 INVx1_ASAP7_75t_SL g12936 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .Y(n_331));
 INVx1_ASAP7_75t_SL g12937 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .Y(n_330));
 INVx1_ASAP7_75t_SL g12938 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .Y(n_329));
 INVx1_ASAP7_75t_SL g12939 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .Y(n_328));
 INVx1_ASAP7_75t_SL g12940 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .Y(n_327));
 INVx1_ASAP7_75t_SL g12941 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .Y(n_326));
 INVx1_ASAP7_75t_SL g12942 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .Y(n_325));
 INVx1_ASAP7_75t_SL g12943 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .Y(n_324));
 INVx1_ASAP7_75t_SL g12944 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .Y(n_323));
 INVx1_ASAP7_75t_SL g12945 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .Y(n_322));
 INVx1_ASAP7_75t_SL g12946 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .Y(n_321));
 INVx1_ASAP7_75t_SL g12947 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .Y(n_320));
 INVx1_ASAP7_75t_SL g12948 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .Y(n_319));
 INVx1_ASAP7_75t_SL g12949 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .Y(n_318));
 INVx1_ASAP7_75t_SL g12950 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .Y(n_317));
 INVx1_ASAP7_75t_SL g12951 (.A(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .Y(n_316));
 INVx1_ASAP7_75t_SL g12952 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .Y(n_315));
 INVx1_ASAP7_75t_SL g12953 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .Y(n_314));
 INVx1_ASAP7_75t_SL g12954 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .Y(n_313));
 INVx1_ASAP7_75t_SL g12955 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .Y(n_312));
 INVxp67_ASAP7_75t_SL g12956 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .Y(n_311));
 INVxp67_ASAP7_75t_SL g12957 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .Y(n_310));
 INVxp67_ASAP7_75t_SL g12958 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .Y(n_309));
 INVxp67_ASAP7_75t_SL g12959 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .Y(n_308));
 INVxp67_ASAP7_75t_SL g12960 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .Y(n_307));
 INVxp67_ASAP7_75t_SL g12961 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .Y(n_306));
 INVxp67_ASAP7_75t_SL g12962 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .Y(n_305));
 INVxp67_ASAP7_75t_SL g12963 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .Y(n_304));
 INVxp67_ASAP7_75t_SL g12964 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_47));
 INVxp67_ASAP7_75t_SL g12966 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .Y(n_301));
 INVxp67_ASAP7_75t_SL g12967 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .Y(n_300));
 INVxp67_ASAP7_75t_SL g12968 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .Y(n_299));
 INVxp67_ASAP7_75t_SL g12969 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .Y(n_298));
 INVxp67_ASAP7_75t_SL g12970 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .Y(n_297));
 INVxp67_ASAP7_75t_SL g12971 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .Y(n_296));
 INVxp67_ASAP7_75t_SL g12972 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .Y(n_295));
 INVxp67_ASAP7_75t_SL g12973 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .Y(n_294));
 INVxp67_ASAP7_75t_SL g12974 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .Y(n_293));
 INVxp67_ASAP7_75t_SL g12975 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .Y(n_292));
 INVxp67_ASAP7_75t_SL g12976 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .Y(n_291));
 INVxp67_ASAP7_75t_SL g12977 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .Y(n_290));
 INVxp67_ASAP7_75t_SL g12978 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .Y(n_289));
 INVxp67_ASAP7_75t_SL g12979 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .Y(n_288));
 INVxp67_ASAP7_75t_SL g12980 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .Y(n_287));
 INVxp67_ASAP7_75t_SL g12981 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .Y(n_286));
 INVxp67_ASAP7_75t_SL g12982 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .Y(n_285));
 INVxp67_ASAP7_75t_SL g12983 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .Y(n_284));
 INVxp67_ASAP7_75t_SL g12984 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .Y(n_283));
 INVxp67_ASAP7_75t_SL g12986 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .Y(n_281));
 INVxp67_ASAP7_75t_SL g12987 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .Y(n_280));
 INVxp67_ASAP7_75t_SL g12988 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .Y(n_279));
 INVxp67_ASAP7_75t_SL g12989 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_47));
 INVxp67_ASAP7_75t_SL g12990 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .Y(n_277));
 INVxp67_ASAP7_75t_SL g12991 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .Y(n_276));
 INVxp67_ASAP7_75t_SL g12992 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .Y(n_275));
 INVxp67_ASAP7_75t_SL g12994 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .Y(n_273));
 INVxp67_ASAP7_75t_SL g12995 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .Y(n_272));
 INVxp67_ASAP7_75t_SL g12997 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_46));
 INVxp67_ASAP7_75t_SL g12998 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .Y(n_269));
 INVxp33_ASAP7_75t_SRAM g12999 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .Y(n_268));
 INVxp67_ASAP7_75t_R g13 (.A(n_22012),
    .Y(n_22013));
 INVxp67_ASAP7_75t_SL g13000 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .Y(n_267));
 INVxp67_ASAP7_75t_SL g13001 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .Y(n_266));
 INVxp67_ASAP7_75t_SL g13002 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .Y(n_265));
 INVxp67_ASAP7_75t_SL g13003 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_47));
 INVxp67_ASAP7_75t_SL g13004 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .Y(n_263));
 INVxp67_ASAP7_75t_SL g13005 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .Y(n_262));
 INVxp67_ASAP7_75t_SL g13006 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .Y(n_261));
 INVxp67_ASAP7_75t_SL g13007 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .Y(n_260));
 INVxp67_ASAP7_75t_SL g13008 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .Y(n_259));
 INVxp67_ASAP7_75t_SL g13009 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .Y(n_258));
 INVxp67_ASAP7_75t_SL g13010 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .Y(n_257));
 INVxp67_ASAP7_75t_SL g13011 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .Y(n_256));
 INVxp67_ASAP7_75t_SL g13012 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .Y(n_255));
 INVxp67_ASAP7_75t_SL g13013 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .Y(n_254));
 INVxp67_ASAP7_75t_SL g13014 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[25]),
    .Y(n_253));
 INVxp67_ASAP7_75t_SL g13015 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .Y(n_252));
 INVxp67_ASAP7_75t_SL g13016 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .Y(n_251));
 INVxp67_ASAP7_75t_SL g13017 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .Y(n_250));
 INVxp33_ASAP7_75t_SRAM g13021 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .Y(n_246));
 INVxp67_ASAP7_75t_SL g13022 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .Y(n_245));
 INVxp67_ASAP7_75t_SL g13023 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .Y(n_244));
 INVxp67_ASAP7_75t_SL g13024 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .Y(n_243));
 INVxp67_ASAP7_75t_SL g13025 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .Y(n_242));
 INVxp67_ASAP7_75t_SL g13027 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .Y(n_240));
 INVxp67_ASAP7_75t_SL g13029 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .Y(n_238));
 INVxp67_ASAP7_75t_SL g13030 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .Y(n_237));
 INVxp67_ASAP7_75t_SL g13031 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .Y(n_236));
 INVxp67_ASAP7_75t_SL g13034 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_47));
 INVxp67_ASAP7_75t_SL g13035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .Y(n_232));
 INVxp67_ASAP7_75t_SL g13036 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .Y(n_231));
 INVxp67_ASAP7_75t_SL g13037 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .Y(n_230));
 INVxp67_ASAP7_75t_SL g13038 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .Y(n_229));
 INVxp67_ASAP7_75t_SL g13039 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .Y(n_228));
 INVxp67_ASAP7_75t_SL g13041 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .Y(n_226));
 INVxp67_ASAP7_75t_SL g13042 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .Y(n_225));
 INVxp67_ASAP7_75t_SL g13043 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .Y(n_224));
 INVxp67_ASAP7_75t_SL g13044 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .Y(n_223));
 INVxp67_ASAP7_75t_SL g13045 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .Y(n_222));
 INVxp67_ASAP7_75t_SL g13046 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .Y(n_221));
 INVxp67_ASAP7_75t_SL g13047 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .Y(n_220));
 INVxp67_ASAP7_75t_SL g13048 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .Y(n_219));
 INVxp67_ASAP7_75t_SL g13049 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .Y(n_218));
 INVxp67_ASAP7_75t_SL g13050 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .Y(n_217));
 INVxp67_ASAP7_75t_SL g13051 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .Y(n_216));
 INVxp67_ASAP7_75t_SL g13052 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .Y(n_215));
 INVxp67_ASAP7_75t_SL g13053 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[25]),
    .Y(n_214));
 INVxp67_ASAP7_75t_SL g13054 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .Y(n_213));
 INVxp67_ASAP7_75t_SL g13056 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .Y(n_211));
 INVxp67_ASAP7_75t_SL g13057 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .Y(n_210));
 INVxp67_ASAP7_75t_SL g13058 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .Y(n_209));
 INVxp67_ASAP7_75t_SL g13059 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .Y(n_208));
 INVxp67_ASAP7_75t_SL g13060 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .Y(n_207));
 INVxp67_ASAP7_75t_SL g13061 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .Y(n_206));
 INVxp67_ASAP7_75t_SL g13062 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .Y(n_205));
 INVxp67_ASAP7_75t_SL g13064 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .Y(n_203));
 INVxp67_ASAP7_75t_SL g13065 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(n_202));
 INVxp67_ASAP7_75t_SL g13066 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .Y(n_201));
 INVxp67_ASAP7_75t_SL g13067 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .Y(n_200));
 INVxp67_ASAP7_75t_SL g13068 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .Y(n_199));
 INVxp67_ASAP7_75t_SL g13069 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .Y(n_198));
 INVxp67_ASAP7_75t_SL g13070 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_47));
 INVxp67_ASAP7_75t_SL g13071 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .Y(n_196));
 INVxp67_ASAP7_75t_SL g13072 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .Y(n_195));
 INVxp67_ASAP7_75t_SL g13073 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .Y(n_194));
 INVxp67_ASAP7_75t_SL g13074 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .Y(n_193));
 INVxp67_ASAP7_75t_SL g13075 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .Y(n_192));
 INVxp67_ASAP7_75t_SL g13076 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .Y(n_191));
 INVxp67_ASAP7_75t_SL g13077 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .Y(n_190));
 INVxp67_ASAP7_75t_SL g13078 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .Y(n_189));
 INVxp67_ASAP7_75t_SL g13079 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .Y(n_188));
 INVxp67_ASAP7_75t_SL g13080 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .Y(n_187));
 INVxp67_ASAP7_75t_SL g13081 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .Y(n_186));
 INVxp67_ASAP7_75t_SRAM g13082 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .Y(n_185));
 INVxp67_ASAP7_75t_SL g13083 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .Y(n_184));
 INVxp67_ASAP7_75t_SL g13084 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .Y(n_183));
 INVxp67_ASAP7_75t_SL g13085 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .Y(n_182));
 INVxp67_ASAP7_75t_SL g13086 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .Y(n_181));
 INVxp67_ASAP7_75t_SL g13088 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .Y(n_179));
 INVxp67_ASAP7_75t_SL g13089 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .Y(n_178));
 INVxp67_ASAP7_75t_SL g13090 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .Y(n_177));
 INVxp67_ASAP7_75t_SL g13091 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .Y(n_176));
 INVxp67_ASAP7_75t_SL g13092 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .Y(n_175));
 INVxp67_ASAP7_75t_SL g13093 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .Y(n_174));
 INVxp67_ASAP7_75t_SL g13094 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .Y(n_173));
 INVxp67_ASAP7_75t_SL g13095 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .Y(n_172));
 INVxp67_ASAP7_75t_SL g13097 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .Y(n_170));
 INVxp67_ASAP7_75t_SL g13098 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .Y(n_169));
 INVxp67_ASAP7_75t_SL g13099 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .Y(n_168));
 XOR2x2_ASAP7_75t_SL g131 (.A(n_13616),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_238),
    .Y(n_13619));
 INVxp67_ASAP7_75t_SL g13100 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_46));
 INVxp67_ASAP7_75t_SL g13101 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .Y(n_166));
 INVxp67_ASAP7_75t_SRAM g13102 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[36]),
    .Y(n_165));
 INVxp67_ASAP7_75t_SL g13103 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .Y(n_164));
 INVxp67_ASAP7_75t_SL g13104 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .Y(n_163));
 INVxp67_ASAP7_75t_SL g13105 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .Y(n_162));
 INVxp67_ASAP7_75t_SL g13106 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .Y(n_161));
 INVxp67_ASAP7_75t_SL g13107 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .Y(n_160));
 INVxp67_ASAP7_75t_SL g13108 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .Y(n_159));
 INVxp67_ASAP7_75t_SL g13109 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .Y(n_158));
 INVxp67_ASAP7_75t_SL g13110 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .Y(n_157));
 INVxp67_ASAP7_75t_SL g13111 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .Y(n_156));
 INVxp67_ASAP7_75t_SL g13112 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .Y(n_155));
 INVxp67_ASAP7_75t_SL g13113 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .Y(n_154));
 INVxp67_ASAP7_75t_SL g13114 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .Y(n_153));
 INVxp67_ASAP7_75t_SL g13115 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .Y(n_152));
 INVxp67_ASAP7_75t_SL g13116 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .Y(n_151));
 INVxp67_ASAP7_75t_SL g13117 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .Y(n_150));
 INVxp67_ASAP7_75t_SL g13118 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .Y(n_149));
 INVxp67_ASAP7_75t_SL g13119 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .Y(n_148));
 INVxp67_ASAP7_75t_SL g13120 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .Y(n_147));
 INVx1_ASAP7_75t_SL g13121 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .Y(n_146));
 INVxp67_ASAP7_75t_SL g13122 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .Y(n_145));
 INVxp67_ASAP7_75t_SL g13123 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .Y(n_144));
 INVxp67_ASAP7_75t_SL g13124 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .Y(n_143));
 INVxp67_ASAP7_75t_SL g13125 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .Y(n_142));
 INVxp67_ASAP7_75t_SL g13127 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .Y(n_140));
 INVxp67_ASAP7_75t_SL g13128 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .Y(n_139));
 INVxp67_ASAP7_75t_SL g13129 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .Y(n_138));
 INVxp67_ASAP7_75t_SL g13132 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .Y(n_135));
 INVxp67_ASAP7_75t_SL g13133 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .Y(n_134));
 INVxp67_ASAP7_75t_SL g13135 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .Y(n_132));
 INVxp67_ASAP7_75t_SL g13136 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .Y(n_131));
 INVxp67_ASAP7_75t_SL g13137 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .Y(n_130));
 INVxp67_ASAP7_75t_SL g13138 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .Y(n_129));
 INVxp67_ASAP7_75t_SL g13139 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_47));
 INVxp67_ASAP7_75t_SL g13141 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .Y(n_126));
 INVxp67_ASAP7_75t_SL g13142 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .Y(n_125));
 INVxp67_ASAP7_75t_SL g13143 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .Y(n_124));
 INVxp67_ASAP7_75t_SL g13144 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .Y(n_123));
 INVxp67_ASAP7_75t_SL g13145 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .Y(n_122));
 INVxp67_ASAP7_75t_SL g13147 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .Y(n_120));
 INVxp67_ASAP7_75t_SL g13148 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .Y(n_119));
 INVxp67_ASAP7_75t_SL g13149 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .Y(n_118));
 INVxp67_ASAP7_75t_SL g13150 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .Y(n_117));
 INVxp67_ASAP7_75t_SL g13151 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .Y(n_116));
 INVxp67_ASAP7_75t_SL g13153 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .Y(n_114));
 INVxp67_ASAP7_75t_SL g13154 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .Y(n_113));
 INVxp67_ASAP7_75t_SL g13155 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .Y(n_112));
 INVxp67_ASAP7_75t_SL g13156 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .Y(n_111));
 INVxp67_ASAP7_75t_SL g13160 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .Y(n_107));
 INVxp67_ASAP7_75t_SL g13161 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .Y(n_106));
 INVxp67_ASAP7_75t_SL g13162 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .Y(n_105));
 INVxp67_ASAP7_75t_SL g13163 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .Y(n_104));
 INVxp67_ASAP7_75t_SL g13164 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .Y(n_103));
 INVxp67_ASAP7_75t_SL g13165 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .Y(n_102));
 INVxp67_ASAP7_75t_SRAM g13166 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .Y(n_101));
 INVxp67_ASAP7_75t_SL g13167 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_46));
 INVx1_ASAP7_75t_SL g13168 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .Y(n_99));
 INVxp67_ASAP7_75t_SL g13169 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .Y(n_98));
 INVxp67_ASAP7_75t_SL g13170 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_47));
 INVxp67_ASAP7_75t_SL g13171 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .Y(n_96));
 INVxp67_ASAP7_75t_SL g13172 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .Y(n_95));
 INVxp67_ASAP7_75t_SL g13173 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .Y(n_94));
 INVxp67_ASAP7_75t_SL g13174 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .Y(n_93));
 INVxp67_ASAP7_75t_SL g13175 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .Y(n_92));
 INVxp67_ASAP7_75t_SL g13176 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .Y(n_91));
 INVxp67_ASAP7_75t_SL g13177 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .Y(n_90));
 INVxp67_ASAP7_75t_SL g13178 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .Y(n_89));
 INVxp67_ASAP7_75t_SL g13179 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .Y(n_88));
 INVxp67_ASAP7_75t_SL g13180 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .Y(n_87));
 INVxp67_ASAP7_75t_SL g13182 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .Y(n_85));
 INVxp67_ASAP7_75t_SL g13183 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .Y(n_84));
 INVxp67_ASAP7_75t_SL g13184 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .Y(n_83));
 INVxp67_ASAP7_75t_SL g13185 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .Y(n_82));
 INVxp67_ASAP7_75t_SL g13186 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_46));
 INVxp67_ASAP7_75t_SL g13187 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .Y(n_80));
 INVxp67_ASAP7_75t_SL g13188 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .Y(n_79));
 INVxp67_ASAP7_75t_SL g13189 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .Y(n_78));
 INVxp67_ASAP7_75t_SL g13190 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .Y(n_77));
 INVxp67_ASAP7_75t_SL g13191 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .Y(n_76));
 INVxp67_ASAP7_75t_SL g13193 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .Y(n_74));
 INVxp67_ASAP7_75t_SL g13194 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .Y(n_73));
 INVxp67_ASAP7_75t_SL g13195 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .Y(n_72));
 INVxp67_ASAP7_75t_SL g13196 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .Y(n_71));
 INVxp67_ASAP7_75t_SL g13197 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .Y(n_70));
 INVxp67_ASAP7_75t_SL g13199 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .Y(n_68));
 INVx1_ASAP7_75t_SL g132 (.A(n_20887),
    .Y(n_23106));
 INVxp67_ASAP7_75t_SL g13200 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .Y(n_67));
 INVxp67_ASAP7_75t_SL g13203 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .Y(n_64));
 INVxp67_ASAP7_75t_SL g13204 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .Y(n_63));
 INVxp67_ASAP7_75t_SL g13205 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .Y(n_62));
 INVxp67_ASAP7_75t_SL g13206 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .Y(n_61));
 INVxp67_ASAP7_75t_SL g13207 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .Y(n_60));
 INVxp67_ASAP7_75t_SL g13208 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[49]),
    .Y(n_59));
 INVxp67_ASAP7_75t_SL g13209 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .Y(n_58));
 INVxp67_ASAP7_75t_SL g13210 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .Y(n_57));
 INVxp67_ASAP7_75t_SL g13211 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .Y(n_56));
 INVxp67_ASAP7_75t_SL g13212 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[17]),
    .Y(n_55));
 INVxp67_ASAP7_75t_SL g13213 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[33]),
    .Y(n_54));
 INVxp67_ASAP7_75t_SL g13214 (.A(u_NV_NVDLA_cmac_u_reg_req_pvld),
    .Y(n_53));
 INVxp67_ASAP7_75t_SL g13217 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[1]),
    .Y(n_50));
 INVxp67_ASAP7_75t_SL g13218 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[21]),
    .Y(n_49));
 INVxp67_ASAP7_75t_SL g13219 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[19]),
    .Y(n_48));
 INVxp67_ASAP7_75t_SL g13220 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[3]),
    .Y(n_47));
 INVx1_ASAP7_75t_SL g13224 (.A(sc2mac_dat_mask[3]),
    .Y(n_45));
 INVx1_ASAP7_75t_SL g13225 (.A(sc2mac_wt_mask[5]),
    .Y(n_44));
 INVx1_ASAP7_75t_SL g13226 (.A(sc2mac_wt_mask[6]),
    .Y(n_43));
 INVx1_ASAP7_75t_SL g13227 (.A(sc2mac_wt_mask[7]),
    .Y(n_42));
 INVx1_ASAP7_75t_SL g13228 (.A(sc2mac_dat_mask[7]),
    .Y(n_41));
 INVx1_ASAP7_75t_SL g13229 (.A(sc2mac_wt_mask[3]),
    .Y(n_40));
 INVx1_ASAP7_75t_SL g13230 (.A(sc2mac_dat_mask[4]),
    .Y(n_39));
 INVx1_ASAP7_75t_SL g13231 (.A(sc2mac_dat_mask[5]),
    .Y(n_38));
 INVx1_ASAP7_75t_SL g13232 (.A(sc2mac_dat_mask[2]),
    .Y(n_37));
 INVx1_ASAP7_75t_SL g13233 (.A(sc2mac_wt_mask[0]),
    .Y(n_36));
 INVx1_ASAP7_75t_SL g13234 (.A(sc2mac_dat_mask[1]),
    .Y(n_35));
 INVx1_ASAP7_75t_SL g13235 (.A(sc2mac_wt_mask[4]),
    .Y(n_34));
 INVx1_ASAP7_75t_SL g13236 (.A(sc2mac_wt_mask[1]),
    .Y(n_33));
 INVx1_ASAP7_75t_SL g13237 (.A(sc2mac_dat_mask[6]),
    .Y(n_32));
 INVx1_ASAP7_75t_SL g13238 (.A(sc2mac_dat_mask[0]),
    .Y(n_31));
 INVx1_ASAP7_75t_SL g13239 (.A(sc2mac_wt_mask[2]),
    .Y(n_30));
 INVx1_ASAP7_75t_SL g13240 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .Y(n_29));
 INVx1_ASAP7_75t_SL g13241 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2),
    .Y(n_28));
 INVx1_ASAP7_75t_SL g13242 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1),
    .Y(n_27));
 INVx1_ASAP7_75t_SL g13243 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .Y(n_26));
 INVx1_ASAP7_75t_SL g13244 (.A(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .Y(n_25));
 INVx1_ASAP7_75t_SL g13245 (.A(csb2cmac_a_req_pvld),
    .Y(n_24));
 INVx1_ASAP7_75t_SL g13246 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .Y(n_23));
 INVx1_ASAP7_75t_SL g13247 (.A(u_NV_NVDLA_cmac_u_core_out_mask[1]),
    .Y(n_22));
 INVx1_ASAP7_75t_SL g13248 (.A(u_NV_NVDLA_cmac_u_core_out_mask[3]),
    .Y(n_21));
 INVx1_ASAP7_75t_SL g13250 (.A(u_NV_NVDLA_cmac_u_core_out_mask[2]),
    .Y(n_19));
 INVx1_ASAP7_75t_SL g13251 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1),
    .Y(n_18));
 INVx1_ASAP7_75t_SL g13252 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .Y(n_17));
 INVx1_ASAP7_75t_SL g13254 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1),
    .Y(n_15));
 INVx1_ASAP7_75t_SL g13255 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .Y(n_14));
 INVx1_ASAP7_75t_SL g13256 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2),
    .Y(n_13));
 INVx1_ASAP7_75t_SL g13257 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2),
    .Y(n_12));
 INVx1_ASAP7_75t_SL g13258 (.A(u_NV_NVDLA_cmac_u_core_out_mask[0]),
    .Y(n_11));
 INVx1_ASAP7_75t_SL g13259 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2),
    .Y(n_10));
 INVx1_ASAP7_75t_SL g13262 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1),
    .Y(n_7));
 INVx1_ASAP7_75t_SL g13263 (.A(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .Y(n_6));
 INVx1_ASAP7_75t_SL g13264 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2),
    .Y(n_5));
 INVx1_ASAP7_75t_SL g13265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1),
    .Y(n_4));
 INVx1_ASAP7_75t_SL g13266 (.A(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .Y(n_3));
 HB1xp67_ASAP7_75t_SL g133 (.A(n_19324),
    .Y(n_19325));
 MAJIxp5_ASAP7_75t_SL g134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_132),
    .C(n_10298),
    .Y(n_10299));
 AO21x1_ASAP7_75t_SL g135 (.A1(n_16324),
    .A2(n_16325),
    .B(n_16326),
    .Y(n_16327));
 AND2x2_ASAP7_75t_SL g136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_0),
    .Y(n_11525));
 XNOR2xp5_ASAP7_75t_SL g137 (.A(n_19316),
    .B(n_26093),
    .Y(n_19326));
 INVxp67_ASAP7_75t_SL g139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_251),
    .Y(n_5751));
 NOR2xp67_ASAP7_75t_SL g14 (.A(n_5738),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_64),
    .Y(n_5739));
 OAI221xp5_ASAP7_75t_SL g140 (.A1(n_5447),
    .A2(n_5449),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_465),
    .B2(n_5451),
    .C(n_5453),
    .Y(n_5454));
 OAI211xp5_ASAP7_75t_SL g1401 (.A1(n_14355),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_282),
    .C(n_9199),
    .Y(n_9200));
 NOR2xp33_ASAP7_75t_SL g1403 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253),
    .B(n_14355),
    .Y(n_9209));
 NAND2xp5_ASAP7_75t_SL g1404 (.A(n_18752),
    .B(n_9198),
    .Y(n_9199));
 NOR2xp33_ASAP7_75t_SL g1407 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_285),
    .Y(n_9201));
 NAND2xp5_ASAP7_75t_SL g1408 (.A(n_14355),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253),
    .Y(n_9206));
 INVx1_ASAP7_75t_SL g1409 (.A(n_8145),
    .Y(n_9198));
 NAND2xp33_ASAP7_75t_SL g141 (.A(n_23580),
    .B(n_5448),
    .Y(n_5449));
 NAND2xp5_ASAP7_75t_SL g142 (.A(n_5448),
    .B(n_5351),
    .Y(n_5453));
 AOI21xp5_ASAP7_75t_SL g14257 (.A1(n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_pvld_3198),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .Y(n_4412));
 AOI21xp5_ASAP7_75t_SL g14258 (.A1(n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_pvld_3195),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .Y(n_4413));
 AOI21xp5_ASAP7_75t_SL g14259 (.A1(n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_pvld_3196),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .Y(n_4414));
 AOI21xp5_ASAP7_75t_SL g14260 (.A1(n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_pvld_3197),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .Y(n_4415));
 NOR2xp33_ASAP7_75t_SL g14261 (.A(n_335),
    .B(u_NV_NVDLA_cmac_u_reg_n_1258),
    .Y(n_4416));
 AOI21xp5_ASAP7_75t_SL g14262 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[0]),
    .A2(n_17870),
    .B(n_19067),
    .Y(n_4417));
 AOI21xp5_ASAP7_75t_SL g14263 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[0]),
    .A2(n_17882),
    .B(n_19095),
    .Y(n_4418));
 AOI21xp5_ASAP7_75t_SL g14264 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[0]),
    .A2(n_17876),
    .B(n_19111),
    .Y(n_4419));
 NOR2xp33_ASAP7_75t_SL g14274 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_164),
    .Y(n_4429));
 NOR2xp33_ASAP7_75t_SL g14275 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_162),
    .Y(n_4430));
 NOR2xp33_ASAP7_75t_SL g14279 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_164),
    .Y(n_4434));
 NOR2xp33_ASAP7_75t_SL g14280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_162),
    .Y(n_4435));
 NOR2xp33_ASAP7_75t_SL g14283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_164),
    .Y(n_4438));
 NOR2xp33_ASAP7_75t_SL g14284 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_162),
    .Y(n_4439));
 NOR2xp33_ASAP7_75t_SL g14288 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_164),
    .Y(n_4443));
 NAND2xp5_ASAP7_75t_SL g143 (.A(n_5448),
    .B(n_5450),
    .Y(n_5451));
 NAND2xp5_ASAP7_75t_SL g144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[16]),
    .B(n_17876),
    .Y(n_5448));
 INVx1_ASAP7_75t_SL g145 (.A(n_17874),
    .Y(n_5351));
 INVx1_ASAP7_75t_SL g146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_465),
    .Y(n_5447));
 INVx1_ASAP7_75t_SL g147 (.A(n_8872),
    .Y(n_8873));
 AND2x2_ASAP7_75t_SL g14715 (.A(n_20877),
    .B(n_20886),
    .Y(n_4965));
 XNOR2x1_ASAP7_75t_SL g14717 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_101),
    .Y(n_4967),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_24));
 XNOR2x1_ASAP7_75t_SL g14719 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_69),
    .Y(n_4969),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_56));
 XOR2xp5_ASAP7_75t_SL g148 (.A(n_21165),
    .B(n_21167),
    .Y(n_21168));
 XNOR2xp5_ASAP7_75t_SL g14864 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_52),
    .Y(n_5126));
 XOR2xp5_ASAP7_75t_SL g14867 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_226),
    .B(n_23387),
    .Y(n_5129));
 MAJIxp5_ASAP7_75t_SL g149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_238),
    .B(n_10103),
    .C(n_7994),
    .Y(n_10104));
 NAND2xp33_ASAP7_75t_SL g14993 (.A(n_5329),
    .B(n_5330),
    .Y(n_5331));
 NAND2xp5_ASAP7_75t_SL g14994 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[18]),
    .B(n_5332),
    .Y(n_5329));
 INVxp33_ASAP7_75t_SL g14995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_5330));
 AND2x2_ASAP7_75t_SL g14999 (.A(n_5329),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_5334));
 NAND2xp5_ASAP7_75t_SL g15 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .B(n_5737),
    .Y(n_5738));
 XNOR2xp5_ASAP7_75t_SL g150 (.A(n_6586),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_26),
    .Y(n_19366));
 OAI21xp33_ASAP7_75t_SL g15001 (.A1(n_24206),
    .A2(n_5342),
    .B(n_5346),
    .Y(n_5347));
 NAND2xp33_ASAP7_75t_SL g15002 (.A(n_5340),
    .B(n_18721),
    .Y(n_5342));
 NAND2xp5_ASAP7_75t_SL g15003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[18]),
    .B(n_17882),
    .Y(n_5340));
 AOI21xp5_ASAP7_75t_SL g15005 (.A1(n_24206),
    .A2(n_5344),
    .B(n_5345),
    .Y(n_5346));
 NOR2xp33_ASAP7_75t_SL g15006 (.A(n_5343),
    .B(n_18721),
    .Y(n_5344));
 INVx1_ASAP7_75t_SL g15007 (.A(n_5340),
    .Y(n_5343));
 NOR2xp33_ASAP7_75t_L g15008 (.A(n_5343),
    .B(n_23932),
    .Y(n_5345));
 INVxp67_ASAP7_75t_SL g15011 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_5348));
 NAND2xp5_ASAP7_75t_SL g15012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[18]),
    .B(n_17876),
    .Y(n_5349));
 INVxp67_ASAP7_75t_SL g15024 (.A(n_5368),
    .Y(n_5369));
 NAND2xp5_ASAP7_75t_SL g15025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[17]),
    .B(n_5332),
    .Y(n_5368));
 NAND2xp5_ASAP7_75t_SL g15027 (.A(n_5368),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_468),
    .Y(n_5371));
 OR2x2_ASAP7_75t_SL g15028 (.A(n_5369),
    .B(n_17936),
    .Y(n_5372));
 INVxp67_ASAP7_75t_SL g15031 (.A(n_5379),
    .Y(n_5380));
 NAND2xp5_ASAP7_75t_SL g15032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[17]),
    .B(n_17882),
    .Y(n_5379));
 OR2x2_ASAP7_75t_SL g15035 (.A(n_5380),
    .B(n_23932),
    .Y(n_5383));
 XNOR2xp5_ASAP7_75t_SL g15038 (.A(n_9659),
    .B(n_18831),
    .Y(n_5393));
 NAND2xp5_ASAP7_75t_SL g15059 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[15]),
    .B(n_5332),
    .Y(n_5426));
 OAI21xp33_ASAP7_75t_SL g15065 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .A2(n_5439),
    .B(n_5443),
    .Y(n_5444));
 NAND2xp33_ASAP7_75t_SL g15066 (.A(n_5438),
    .B(n_9988),
    .Y(n_5439));
 NAND2xp5_ASAP7_75t_SL g15067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[15]),
    .B(n_17876),
    .Y(n_5438));
 AOI21xp5_ASAP7_75t_SL g15068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .A2(n_5441),
    .B(n_5442),
    .Y(n_5443));
 NOR2xp33_ASAP7_75t_SL g15069 (.A(n_5440),
    .B(n_9988),
    .Y(n_5441));
 INVx1_ASAP7_75t_SL g15070 (.A(n_5438),
    .Y(n_5440));
 NOR2xp33_ASAP7_75t_SL g15071 (.A(n_5440),
    .B(n_17874),
    .Y(n_5442));
 AOI21x1_ASAP7_75t_SL g15074 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_483),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_442),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_407),
    .Y(n_5456));
 INVxp67_ASAP7_75t_SL g15081 (.A(n_13090),
    .Y(n_5471));
 NOR2xp67_ASAP7_75t_SL g15091 (.A(n_7343),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_271),
    .Y(n_5487));
 AND2x2_ASAP7_75t_SL g15094 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_740),
    .Y(n_5492));
 NAND2xp5_ASAP7_75t_SL g151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_175),
    .Y(n_19542));
 OAI21xp33_ASAP7_75t_SL g15103 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .A2(n_5505),
    .B(n_5509),
    .Y(n_5510));
 NAND2xp5_ASAP7_75t_SL g15104 (.A(n_5504),
    .B(n_9977),
    .Y(n_5505));
 AOI21xp5_ASAP7_75t_SL g15105 (.A1(n_5507),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .B(n_5508),
    .Y(n_5509));
 NOR2xp33_ASAP7_75t_SL g15106 (.A(n_5506),
    .B(n_9977),
    .Y(n_5507));
 INVxp67_ASAP7_75t_SL g15107 (.A(n_5504),
    .Y(n_5506));
 NOR2xp33_ASAP7_75t_SL g15108 (.A(n_5506),
    .B(n_23932),
    .Y(n_5508));
 NOR2xp67_ASAP7_75t_SL g15118 (.A(n_6191),
    .B(n_11418),
    .Y(n_5544));
 NOR2xp67_ASAP7_75t_SL g15119 (.A(n_12120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_46),
    .Y(n_5548));
 XNOR2xp5_ASAP7_75t_SL g15121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_89),
    .B(n_10916),
    .Y(n_5553));
 INVx1_ASAP7_75t_SL g15133 (.A(n_12303),
    .Y(n_5564));
 MAJx2_ASAP7_75t_SL g15143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_172),
    .Y(n_5575));
 NAND2x1_ASAP7_75t_L g15146 (.A(n_10094),
    .B(n_5583),
    .Y(n_5584));
 XNOR2x1_ASAP7_75t_SL g15147 (.B(n_5582),
    .Y(n_5583),
    .A(n_13330));
 NAND2x1p5_ASAP7_75t_SL g15168 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .B(n_4275),
    .Y(n_3806));
 AOI21xp5_ASAP7_75t_SL g15171 (.A1(n_22487),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_290),
    .B(n_5616),
    .Y(n_5617));
 NOR2xp67_ASAP7_75t_SL g15172 (.A(n_22489),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_271),
    .Y(n_5616));
 XNOR2x1_ASAP7_75t_SL g15179 (.B(n_14340),
    .Y(n_5627),
    .A(n_26049));
 NOR2xp67_ASAP7_75t_SL g15185 (.A(n_26222),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_271),
    .Y(n_5630));
 XNOR2xp5_ASAP7_75t_SL g15186 (.A(n_23835),
    .B(n_17413),
    .Y(n_5637));
 OAI22xp5_ASAP7_75t_SL g15192 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_99),
    .A2(n_5644),
    .B1(n_12622),
    .B2(n_5643),
    .Y(n_5645));
 INVx1_ASAP7_75t_SL g15193 (.A(n_5643),
    .Y(n_5644));
 MAJx2_ASAP7_75t_SL g15194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_71),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_34),
    .Y(n_5643));
 INVxp67_ASAP7_75t_SL g15197 (.A(n_15457),
    .Y(n_5649));
 HB1xp67_ASAP7_75t_SL g152 (.A(n_19958),
    .Y(n_6783));
 HB1xp67_ASAP7_75t_SL g15208 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_89),
    .Y(n_5664));
 NOR2x1p5_ASAP7_75t_SL g15216 (.A(n_5679),
    .B(n_5680),
    .Y(n_5681));
 INVxp67_ASAP7_75t_SL g15217 (.A(n_2158),
    .Y(n_5679));
 XNOR2xp5_ASAP7_75t_SL g15218 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_305),
    .B(n_7783),
    .Y(n_5680));
 INVx1_ASAP7_75t_SL g15219 (.A(n_5681),
    .Y(n_5683));
 INVx1_ASAP7_75t_SL g15231 (.A(n_18815),
    .Y(n_5697));
 XOR2xp5_ASAP7_75t_SL g15258 (.A(n_10346),
    .B(n_5743),
    .Y(n_5744));
 OAI22xp5_ASAP7_75t_SL g15259 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_78),
    .A2(n_5740),
    .B1(n_5741),
    .B2(n_5742),
    .Y(n_5743));
 NAND2xp5_ASAP7_75t_SL g15260 (.A(n_2831),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .Y(n_5740));
 INVx1_ASAP7_75t_SL g15261 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_78),
    .Y(n_5741));
 INVx1_ASAP7_75t_SL g15262 (.A(n_5740),
    .Y(n_5742));
 XNOR2xp5_ASAP7_75t_SL g15290 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_213),
    .B(n_26124),
    .Y(n_5780));
 XNOR2x1_ASAP7_75t_SL g15297 (.B(n_5783),
    .Y(n_5784),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_583));
 AND2x2_ASAP7_75t_SL g15298 (.A(n_2165),
    .B(n_22806),
    .Y(n_5783));
 NOR2xp33_ASAP7_75t_SL g153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_209),
    .Y(n_19539));
 AO21x1_ASAP7_75t_SL g15300 (.A1(n_5787),
    .A2(n_9821),
    .B(n_5792),
    .Y(n_5793));
 NAND2xp33_ASAP7_75t_SL g15301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_168),
    .Y(n_5787));
 NOR2xp33_ASAP7_75t_SL g15306 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_168),
    .Y(n_5792));
 AOI21x1_ASAP7_75t_SL g15308 (.A1(n_7981),
    .A2(n_5798),
    .B(n_5799),
    .Y(n_5800));
 INVx1_ASAP7_75t_SL g15310 (.A(n_5796),
    .Y(n_5794));
 NAND2xp5_ASAP7_75t_SL g15311 (.A(n_5796),
    .B(n_11241),
    .Y(n_5798));
 INVx1_ASAP7_75t_SL g15314 (.A(n_18577),
    .Y(n_5799));
 OAI22xp5_ASAP7_75t_SL g15316 (.A1(n_23824),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_77),
    .B1(n_23825),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_78),
    .Y(n_5804));
 AND2x2_ASAP7_75t_SL g15322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_656),
    .B(n_7595),
    .Y(n_5806));
 INVx1_ASAP7_75t_SL g15346 (.A(n_14643),
    .Y(n_5849));
 XNOR2xp5_ASAP7_75t_SL g15357 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_67),
    .B(n_13770),
    .Y(n_4231));
 NAND2xp33_ASAP7_75t_SL g15364 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_204),
    .B(n_22435),
    .Y(n_5880));
 INVx1_ASAP7_75t_SL g15365 (.A(n_2151),
    .Y(n_5881));
 XOR2xp5_ASAP7_75t_SL g15366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_88),
    .B(n_18850),
    .Y(n_5890));
 NAND2xp5_ASAP7_75t_SL g15369 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(n_14523),
    .Y(n_5886));
 OAI22xp5_ASAP7_75t_SL g15375 (.A1(n_5894),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_56),
    .B1(n_5895),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_55),
    .Y(n_5896));
 NAND2xp5_ASAP7_75t_SL g15376 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .Y(n_5894));
 OAI22xp5_ASAP7_75t_SL g15379 (.A1(n_5909),
    .A2(n_7189),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_24),
    .B2(n_19827),
    .Y(n_5910));
 INVxp67_ASAP7_75t_SL g15383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_95),
    .Y(n_5904));
 OAI22xp5_ASAP7_75t_SL g154 (.A1(n_26046),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_187),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_188),
    .B2(n_8344),
    .Y(n_8348));
 XOR2x1_ASAP7_75t_SL g15400 (.A(n_5929),
    .Y(n_5930),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_583));
 AND2x2_ASAP7_75t_SL g15401 (.A(n_19838),
    .B(n_22315),
    .Y(n_5929));
 NAND2x1_ASAP7_75t_SL g15402 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(n_11770),
    .Y(n_5948));
 MAJIxp5_ASAP7_75t_SL g15406 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_73),
    .Y(n_5955));
 INVxp67_ASAP7_75t_SL g15408 (.A(n_23665),
    .Y(n_5959));
 INVx1_ASAP7_75t_SL g15410 (.A(n_5955),
    .Y(n_5961));
 NAND2xp5_ASAP7_75t_SL g15434 (.A(n_11868),
    .B(n_9992),
    .Y(n_6008));
 AND2x2_ASAP7_75t_SL g15439 (.A(n_9992),
    .B(n_6016),
    .Y(n_6017));
 OAI211xp5_ASAP7_75t_SL g15440 (.A1(n_19928),
    .A2(n_6038),
    .B(n_19930),
    .C(n_6043),
    .Y(n_6044));
 NAND3xp33_ASAP7_75t_SL g15442 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .B(n_14152),
    .C(n_6037),
    .Y(n_6038));
 NAND2xp5_ASAP7_75t_SL g15443 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[17]),
    .B(n_17876),
    .Y(n_6037));
 INVx1_ASAP7_75t_SL g15446 (.A(n_6037),
    .Y(n_6039));
 NAND2xp5_ASAP7_75t_SL g15447 (.A(n_6037),
    .B(n_5351),
    .Y(n_6043));
 MAJx2_ASAP7_75t_SL g15457 (.A(n_10144),
    .B(n_22000),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_220),
    .Y(n_6063));
 INVxp67_ASAP7_75t_SL g15468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_737),
    .Y(n_6082));
 AOI21xp5_ASAP7_75t_SL g15478 (.A1(n_12888),
    .A2(n_14089),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_297),
    .Y(n_6102));
 INVxp67_ASAP7_75t_SL g15482 (.A(n_6102),
    .Y(n_6107));
 INVx1_ASAP7_75t_SL g15484 (.A(n_18820),
    .Y(n_6109));
 XNOR2xp5_ASAP7_75t_SL g15486 (.A(n_18729),
    .B(n_6116),
    .Y(n_6117));
 XNOR2x1_ASAP7_75t_SL g15488 (.B(n_6115),
    .Y(n_6116),
    .A(n_6113));
 XNOR2x1_ASAP7_75t_SL g15489 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_559),
    .Y(n_6113),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_783));
 INVx1_ASAP7_75t_SL g15490 (.A(n_6114),
    .Y(n_6115));
 AND2x2_ASAP7_75t_SL g15491 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_718),
    .Y(n_6114));
 MAJx2_ASAP7_75t_SL g15492 (.A(n_25996),
    .B(n_18729),
    .C(n_6116),
    .Y(n_6119));
 INVx1_ASAP7_75t_SL g155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_188));
 XNOR2xp5_ASAP7_75t_SL g15502 (.A(n_11726),
    .B(n_5641),
    .Y(n_6141));
 HB1xp67_ASAP7_75t_SL g15503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_303),
    .Y(n_6179));
 NAND2xp5_ASAP7_75t_SL g15504 (.A(n_6832),
    .B(n_12620),
    .Y(n_6189));
 NOR2xp67_ASAP7_75t_SL g15505 (.A(n_6832),
    .B(n_12620),
    .Y(n_6190));
 AOI21xp5_ASAP7_75t_SL g15506 (.A1(n_14723),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_243),
    .Y(n_6191));
 NAND2xp5_ASAP7_75t_SL g15512 (.A(n_10666),
    .B(n_10117),
    .Y(n_6194));
 AOI21x1_ASAP7_75t_SL g15513 (.A1(n_6198),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_319),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_313),
    .Y(n_6199));
 INVxp67_ASAP7_75t_SL g15514 (.A(n_9035),
    .Y(n_6198));
 NAND2xp5_ASAP7_75t_SL g15515 (.A(n_6200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_307),
    .Y(n_6201));
 HB1xp67_ASAP7_75t_SL g15516 (.A(n_10161),
    .Y(n_6200));
 OAI21xp5_ASAP7_75t_SL g15517 (.A1(n_6202),
    .A2(n_6199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_307),
    .Y(n_6203));
 INVxp67_ASAP7_75t_SL g15518 (.A(n_6200),
    .Y(n_6202));
 AOI21xp5_ASAP7_75t_SL g15519 (.A1(n_10162),
    .A2(n_6194),
    .B(n_5697),
    .Y(n_6204));
 AND2x2_ASAP7_75t_SL g15520 (.A(n_6194),
    .B(n_18815),
    .Y(n_6205));
 MAJx2_ASAP7_75t_SL g15524 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_132),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_152),
    .Y(n_6209));
 XNOR2x2_ASAP7_75t_SL g15525 (.A(n_6210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_182),
    .Y(n_6211));
 INVxp67_ASAP7_75t_SL g15526 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_157),
    .Y(n_6210));
 XOR2xp5_ASAP7_75t_SL g15530 (.A(n_22057),
    .B(n_6237),
    .Y(n_6238));
 OR2x2_ASAP7_75t_SL g15532 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_0),
    .Y(n_6237));
 MAJIxp5_ASAP7_75t_SL g15533 (.A(n_6125),
    .B(n_6240),
    .C(n_6241),
    .Y(n_6242));
 INVxp67_ASAP7_75t_SL g15534 (.A(n_6237),
    .Y(n_6240));
 INVxp67_ASAP7_75t_SL g15535 (.A(n_22057),
    .Y(n_6241));
 NAND2x1_ASAP7_75t_SL g15536 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_102),
    .B(n_6237),
    .Y(n_6243));
 INVx1_ASAP7_75t_SL g15537 (.A(n_15626),
    .Y(n_6251));
 MAJIxp5_ASAP7_75t_SL g15542 (.A(n_6255),
    .B(n_6256),
    .C(n_2439),
    .Y(n_6257));
 HB1xp67_ASAP7_75t_SL g15543 (.A(n_24200),
    .Y(n_6256));
 AOI21xp5_ASAP7_75t_SL g15550 (.A1(n_9801),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_309),
    .B(n_6264),
    .Y(n_6265));
 INVxp67_ASAP7_75t_SL g15551 (.A(n_8787),
    .Y(n_6264));
 INVx1_ASAP7_75t_SL g15553 (.A(n_8784),
    .Y(n_6266));
 AND2x2_ASAP7_75t_SL g15562 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .Y(n_6279));
 OAI22xp5_ASAP7_75t_SL g15569 (.A1(n_18933),
    .A2(n_17417),
    .B1(n_17416),
    .B2(n_6295),
    .Y(n_6296));
 OAI22x1_ASAP7_75t_SL g15570 (.A1(n_18933),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37),
    .B2(n_6295),
    .Y(n_2437));
 XNOR2x1_ASAP7_75t_SL g15572 (.B(n_6303),
    .Y(n_6304),
    .A(n_6302));
 XNOR2x1_ASAP7_75t_SL g15573 (.B(n_6301),
    .Y(n_6302),
    .A(n_6300));
 NAND2x1p5_ASAP7_75t_SL g15574 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(n_2335),
    .Y(n_6300));
 AND2x2_ASAP7_75t_SL g15575 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .B(n_6972),
    .Y(n_6301));
 INVx1_ASAP7_75t_SL g15576 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_27),
    .Y(n_6303));
 MAJIxp5_ASAP7_75t_SL g15577 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_27),
    .B(n_6300),
    .C(n_6301),
    .Y(n_6305));
 NAND2xp5_ASAP7_75t_SL g15586 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_270),
    .Y(n_6313));
 INVx1_ASAP7_75t_SL g15595 (.A(n_19790),
    .Y(n_6323));
 NOR2xp67_ASAP7_75t_SL g15600 (.A(n_6352),
    .B(n_6353),
    .Y(n_6354));
 MAJIxp5_ASAP7_75t_SL g15601 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_9),
    .C(n_5517),
    .Y(n_6352));
 XNOR2xp5_ASAP7_75t_SL g15602 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_11),
    .Y(n_6353));
 INVxp67_ASAP7_75t_SRAM g15606 (.A(n_14344),
    .Y(n_6365));
 OAI21xp5_ASAP7_75t_SL g15608 (.A1(n_6361),
    .A2(n_8520),
    .B(n_8519),
    .Y(n_6368));
 INVxp67_ASAP7_75t_SL g15609 (.A(n_6371),
    .Y(n_6372));
 XNOR2xp5_ASAP7_75t_SL g15610 (.A(n_6369),
    .B(n_6370),
    .Y(n_6371));
 MAJIxp5_ASAP7_75t_SL g15611 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_103),
    .Y(n_6369));
 OAI22xp33_ASAP7_75t_SL g15612 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_117),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_4),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_149),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_118),
    .Y(n_6370));
 MAJIxp5_ASAP7_75t_SL g15615 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_4),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_118),
    .C(n_6369),
    .Y(n_6377));
 NAND2xp33_ASAP7_75t_SL g15618 (.A(n_6381),
    .B(n_22614),
    .Y(n_6382));
 NAND2xp5_ASAP7_75t_SL g15619 (.A(n_17870),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[15]),
    .Y(n_6381));
 NOR2xp33_ASAP7_75t_SL g15623 (.A(n_6383),
    .B(n_22614),
    .Y(n_6384));
 INVxp67_ASAP7_75t_SL g15624 (.A(n_6381),
    .Y(n_6383));
 AND2x2_ASAP7_75t_SL g15625 (.A(n_17870),
    .B(n_6381),
    .Y(n_6385));
 XNOR2x1_ASAP7_75t_SL g15626 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_13),
    .Y(n_6411),
    .A(n_6410));
 MAJx2_ASAP7_75t_SL g15627 (.A(n_21136),
    .B(n_21135),
    .C(n_6409),
    .Y(n_6410));
 NAND2xp5_ASAP7_75t_SL g15630 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_716),
    .Y(n_6409));
 OAI21x1_ASAP7_75t_SL g15631 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_83),
    .A2(n_6410),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_86),
    .Y(n_3657));
 INVxp67_ASAP7_75t_SRAM g15640 (.A(n_20814),
    .Y(n_6420));
 HB1xp67_ASAP7_75t_SL g15641 (.A(n_20809),
    .Y(n_6421));
 HB1xp67_ASAP7_75t_SL g15650 (.A(n_12549),
    .Y(n_6430));
 INVx1_ASAP7_75t_SL g15651 (.A(n_24769),
    .Y(n_6431));
 XNOR2x1_ASAP7_75t_SL g15654 (.B(n_6438),
    .Y(n_6439),
    .A(n_19776));
 INVxp67_ASAP7_75t_SL g15656 (.A(n_6437),
    .Y(n_6438));
 NAND2xp5_ASAP7_75t_SL g15657 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(n_6437));
 MAJx2_ASAP7_75t_SL g15661 (.A(n_19774),
    .B(n_6437),
    .C(n_19775),
    .Y(n_6444));
 INVx1_ASAP7_75t_SL g15666 (.A(n_18863),
    .Y(n_6463));
 INVx1_ASAP7_75t_SL g15673 (.A(n_26101),
    .Y(n_6471));
 MAJIxp5_ASAP7_75t_SL g15674 (.A(n_19484),
    .B(n_19478),
    .C(n_18863),
    .Y(n_6474));
 NOR2x1p5_ASAP7_75t_SL g15675 (.A(n_10523),
    .B(n_6478),
    .Y(n_6479));
 XOR2x2_ASAP7_75t_SL g15676 (.A(n_6476),
    .B(n_6477),
    .Y(n_6478));
 XNOR2xp5_ASAP7_75t_SL g15677 (.A(n_18731),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_147),
    .Y(n_6476));
 XNOR2xp5_ASAP7_75t_SL g15679 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_8),
    .Y(n_6477));
 NAND2x1_ASAP7_75t_SL g15680 (.A(n_10523),
    .B(n_6478),
    .Y(n_6480));
 MAJIxp5_ASAP7_75t_SL g15681 (.A(n_6477),
    .B(n_6481),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_147),
    .Y(n_6483));
 INVxp67_ASAP7_75t_SL g15682 (.A(n_18731),
    .Y(n_6481));
 AND2x4_ASAP7_75t_SL g157 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(n_14523),
    .Y(n_20301));
 INVxp67_ASAP7_75t_SL g15723 (.A(n_11767),
    .Y(n_6546));
 MAJIxp5_ASAP7_75t_SL g15747 (.A(n_18865),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_146),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_207));
 MAJIxp5_ASAP7_75t_SL g15751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_112),
    .C(n_9810),
    .Y(n_6579));
 MAJIxp5_ASAP7_75t_SL g15757 (.A(n_9325),
    .B(n_9324),
    .C(n_6585),
    .Y(n_6586));
 MAJIxp5_ASAP7_75t_SL g15760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_75),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_79),
    .Y(n_6585));
 MAJIxp5_ASAP7_75t_SL g15761 (.A(n_19365),
    .B(n_6588),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_26),
    .Y(n_6589));
 INVxp67_ASAP7_75t_SL g15762 (.A(n_6586),
    .Y(n_6588));
 XOR2xp5_ASAP7_75t_SL g15763 (.A(n_6591),
    .B(n_9326),
    .Y(n_6592));
 INVxp67_ASAP7_75t_SL g15765 (.A(n_6585),
    .Y(n_6591));
 MAJx2_ASAP7_75t_SL g15768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_264),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_212),
    .C(n_23380),
    .Y(n_6593));
 MAJIxp5_ASAP7_75t_SL g15771 (.A(n_2620),
    .B(n_6599),
    .C(n_9963),
    .Y(n_6601));
 XNOR2xp5_ASAP7_75t_SL g15773 (.A(n_6866),
    .B(n_6604),
    .Y(n_6605));
 XNOR2x1_ASAP7_75t_SL g15774 (.B(n_6603),
    .Y(n_6604),
    .A(n_6602));
 NAND2xp5_ASAP7_75t_SL g15775 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .Y(n_6602));
 AND2x2_ASAP7_75t_SL g15776 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(n_15192),
    .Y(n_6603));
 MAJIxp5_ASAP7_75t_SL g15777 (.A(n_6866),
    .B(n_6603),
    .C(n_6602),
    .Y(n_6606));
 OAI21xp5_ASAP7_75t_SL g15778 (.A1(n_6610),
    .A2(n_6616),
    .B(n_6617),
    .Y(n_6618));
 INVx2_ASAP7_75t_SL g15779 (.A(n_18866),
    .Y(n_6610));
 NAND2xp5_ASAP7_75t_SL g15783 (.A(n_6614),
    .B(n_6615),
    .Y(n_6616));
 INVx1_ASAP7_75t_SL g15784 (.A(n_18867),
    .Y(n_6614));
 INVx1_ASAP7_75t_SL g15788 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_119),
    .Y(n_6615));
 NAND3xp33_ASAP7_75t_SL g15789 (.A(n_6610),
    .B(n_6615),
    .C(n_18867),
    .Y(n_6617));
 NAND2xp5_ASAP7_75t_SL g15790 (.A(n_6619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_119),
    .Y(n_6620));
 OAI22xp33_ASAP7_75t_SL g15791 (.A1(n_6610),
    .A2(n_6614),
    .B1(n_18867),
    .B2(n_18866),
    .Y(n_6619));
 XOR2xp5_ASAP7_75t_SL g158 (.A(n_12653),
    .B(n_26081),
    .Y(n_20101));
 NAND2xp5_ASAP7_75t_SL g15804 (.A(n_7573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_180),
    .Y(n_6639));
 OAI22xp5_ASAP7_75t_SL g15806 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_135),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_120),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_134),
    .Y(n_6635));
 HB1xp67_ASAP7_75t_SL g15815 (.A(n_5886),
    .Y(n_6646));
 AOI21xp5_ASAP7_75t_SL g15822 (.A1(n_6655),
    .A2(n_6656),
    .B(n_6657),
    .Y(n_6658));
 NAND2xp5_ASAP7_75t_SL g15823 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_214),
    .Y(n_6655));
 OAI21xp5_ASAP7_75t_SL g15824 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_198),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_201),
    .Y(n_6656));
 NOR2xp33_ASAP7_75t_SL g15825 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_214),
    .Y(n_6657));
 XOR2xp5_ASAP7_75t_SL g15826 (.A(n_13651),
    .B(n_6660),
    .Y(n_6661));
 HB1xp67_ASAP7_75t_SL g15827 (.A(n_6658),
    .Y(n_6660));
 XNOR2xp5_ASAP7_75t_SL g15828 (.A(n_6656),
    .B(n_19133),
    .Y(n_6666));
 AND2x2_ASAP7_75t_SL g15834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_672),
    .B(n_2160),
    .Y(n_6667));
 AND2x2_ASAP7_75t_SL g15835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_576),
    .B(n_2168),
    .Y(n_6668));
 MAJIxp5_ASAP7_75t_SL g15837 (.A(n_6667),
    .B(n_6668),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_737),
    .Y(n_6673));
 INVx2_ASAP7_75t_SL g15840 (.A(n_20673),
    .Y(n_6675));
 INVx1_ASAP7_75t_SL g15844 (.A(n_22892),
    .Y(n_6676));
 MAJIxp5_ASAP7_75t_SL g15850 (.A(n_6675),
    .B(n_2435),
    .C(n_15000),
    .Y(n_6687));
 MAJIxp5_ASAP7_75t_SL g15872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_101),
    .B(n_13769),
    .C(n_22622),
    .Y(n_6710));
 NAND2xp5_ASAP7_75t_SL g15886 (.A(n_16707),
    .B(n_10177),
    .Y(n_6730));
 INVx1_ASAP7_75t_SL g15891 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_320),
    .Y(n_6724));
 NAND2xp5_ASAP7_75t_SL g15892 (.A(n_11452),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_320),
    .Y(n_6727));
 INVxp67_ASAP7_75t_SL g15896 (.A(n_16705),
    .Y(n_6733));
 XNOR2x1_ASAP7_75t_SL g15899 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_182),
    .Y(n_6742),
    .A(n_6741));
 MAJIxp5_ASAP7_75t_SRAM g159 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_683),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_587),
    .C(n_7096),
    .Y(n_7097));
 XNOR2x1_ASAP7_75t_SL g15900 (.B(n_6740),
    .Y(n_6741),
    .A(n_6737));
 NAND2xp5_ASAP7_75t_SL g15901 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .B(n_12124),
    .Y(n_6737));
 OAI22xp5_ASAP7_75t_SL g15902 (.A1(n_13719),
    .A2(n_6738),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_107),
    .B2(n_6739),
    .Y(n_6740));
 INVx1_ASAP7_75t_SL g15903 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_107),
    .Y(n_6738));
 INVx1_ASAP7_75t_SL g15904 (.A(n_13719),
    .Y(n_6739));
 MAJIxp5_ASAP7_75t_SL g15909 (.A(n_6737),
    .B(n_6747),
    .C(n_6748),
    .Y(n_6749));
 INVxp67_ASAP7_75t_SL g15910 (.A(n_6738),
    .Y(n_6747));
 INVxp67_ASAP7_75t_SL g15911 (.A(n_6739),
    .Y(n_6748));
 INVx1_ASAP7_75t_SL g15916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_115),
    .Y(n_6751));
 XOR2x2_ASAP7_75t_SL g15917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_142),
    .B(n_6753),
    .Y(n_6754));
 INVx1_ASAP7_75t_SL g15918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_51),
    .Y(n_6753));
 MAJIxp5_ASAP7_75t_SL g15920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_236),
    .B(n_9541),
    .C(n_9544),
    .Y(n_6758));
 XNOR2x1_ASAP7_75t_SL g15925 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_182),
    .Y(n_6769),
    .A(n_18871));
 AND2x2_ASAP7_75t_SL g15931 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(n_12124),
    .Y(n_6766));
 MAJx2_ASAP7_75t_R g15932 (.A(n_18871),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_139),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_131),
    .Y(n_6771));
 AO21x1_ASAP7_75t_SL g15934 (.A1(n_6772),
    .A2(n_6766),
    .B(n_6773),
    .Y(n_6774));
 NAND2xp33_ASAP7_75t_SL g15935 (.A(n_13727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_107),
    .Y(n_6772));
 NOR2xp33_ASAP7_75t_SL g15936 (.A(n_13727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_107),
    .Y(n_6773));
 INVxp67_ASAP7_75t_SL g15944 (.A(n_6783),
    .Y(n_6784));
 NAND2xp33_ASAP7_75t_SL g15945 (.A(n_6783),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_307),
    .Y(n_5796));
 AND2x2_ASAP7_75t_SL g15946 (.A(n_8901),
    .B(n_6313),
    .Y(n_6787));
 AOI22xp33_ASAP7_75t_SL g15947 (.A1(n_8901),
    .A2(n_19959),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_270),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_274),
    .Y(n_6788));
 HB1xp67_ASAP7_75t_SL g15955 (.A(n_20844),
    .Y(n_6806));
 XNOR2xp5_ASAP7_75t_SL g15971 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_33),
    .B(n_15098),
    .Y(n_6824));
 INVx1_ASAP7_75t_SL g15975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_249),
    .Y(n_6830));
 AOI21xp5_ASAP7_75t_SL g15976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_239),
    .A2(n_6824),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_240),
    .Y(n_6832));
 INVx1_ASAP7_75t_SL g15980 (.A(n_21668),
    .Y(n_6836));
 NAND2x1_ASAP7_75t_SL g15999 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(n_2990),
    .Y(n_6853));
 NAND2xp33_ASAP7_75t_SL g16 (.A(n_13363),
    .B(n_8167),
    .Y(n_18003));
 INVxp67_ASAP7_75t_SL g160 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_213),
    .Y(n_10237));
 NAND2x1_ASAP7_75t_R g16004 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(n_6861),
    .Y(n_6862));
 MAJIxp5_ASAP7_75t_SL g16008 (.A(n_18710),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_49),
    .C(n_6862),
    .Y(n_6866));
 MAJIxp5_ASAP7_75t_SL g16013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_37),
    .Y(n_6871));
 OAI21xp5_ASAP7_75t_SL g16014 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_174),
    .Y(n_6872));
 XOR2xp5_ASAP7_75t_SL g16015 (.A(n_6871),
    .B(n_10520),
    .Y(n_6877));
 NAND2xp5_ASAP7_75t_SL g16018 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_740),
    .B(n_6879),
    .Y(n_6880));
 XOR2xp5_ASAP7_75t_SL g16024 (.A(n_21963),
    .B(n_10803),
    .Y(n_6888));
 MAJIxp5_ASAP7_75t_SL g16025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_207),
    .B(n_6895),
    .C(n_18719),
    .Y(n_6896));
 INVxp67_ASAP7_75t_SL g16026 (.A(n_6894),
    .Y(n_6895));
 XNOR2xp5_ASAP7_75t_SL g16027 (.A(n_6890),
    .B(n_26054),
    .Y(n_6894));
 AND2x2_ASAP7_75t_SL g16028 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(n_2359),
    .Y(n_6890));
 MAJIxp5_ASAP7_75t_SL g16034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_36),
    .B(n_6890),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_20),
    .Y(n_6902));
 NAND2x1p5_ASAP7_75t_L g16039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(n_19645),
    .Y(n_6903));
 AND2x2_ASAP7_75t_SL g16040 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(n_6904));
 NAND2xp5_ASAP7_75t_SL g16041 (.A(n_14975),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .Y(n_6905));
 XOR2xp5_ASAP7_75t_SL g16044 (.A(n_6904),
    .B(n_6903),
    .Y(n_6910));
 XOR2xp5_ASAP7_75t_SL g16045 (.A(n_6916),
    .B(n_10886),
    .Y(n_6917));
 XNOR2xp5_ASAP7_75t_SL g16046 (.A(n_26098),
    .B(n_26055),
    .Y(n_6916));
 XNOR2xp5_ASAP7_75t_SL g16054 (.A(n_6924),
    .B(n_6925),
    .Y(n_6926));
 MAJx2_ASAP7_75t_SL g16056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_88),
    .Y(n_6923));
 INVx1_ASAP7_75t_L g16058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_212),
    .Y(n_6925));
 INVxp67_ASAP7_75t_SL g16060 (.A(n_6923),
    .Y(n_6928));
 HB1xp67_ASAP7_75t_SL g16061 (.A(n_10471),
    .Y(n_6929));
 XNOR2xp5_ASAP7_75t_SL g16062 (.A(n_22005),
    .B(n_6939),
    .Y(n_6940));
 MAJIxp5_ASAP7_75t_SL g16063 (.A(n_6935),
    .B(n_6937),
    .C(n_6938),
    .Y(n_6939));
 HB1xp67_ASAP7_75t_SL g16064 (.A(n_10470),
    .Y(n_6935));
 INVxp67_ASAP7_75t_SL g16069 (.A(n_6936),
    .Y(n_6937));
 XNOR2xp5_ASAP7_75t_SL g16070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_80),
    .Y(n_6936));
 XNOR2x1_ASAP7_75t_SL g16071 (.B(n_24404),
    .Y(n_6938),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_20));
 NOR2xp33_ASAP7_75t_SL g16072 (.A(n_6939),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_205),
    .Y(n_6941));
 NAND2xp33_ASAP7_75t_SL g16073 (.A(n_6939),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_205),
    .Y(n_6942));
 XNOR2xp5_ASAP7_75t_SL g16074 (.A(n_6938),
    .B(n_6943),
    .Y(n_3279));
 XOR2xp5_ASAP7_75t_SL g16075 (.A(n_10470),
    .B(n_6936),
    .Y(n_6943));
 AND2x2_ASAP7_75t_SL g16079 (.A(n_9034),
    .B(n_9032),
    .Y(n_6949));
 MAJIxp5_ASAP7_75t_SL g16081 (.A(n_6950),
    .B(n_6954),
    .C(n_6957),
    .Y(n_6958));
 OAI21xp5_ASAP7_75t_SL g16082 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_179),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_180),
    .Y(n_6950));
 OAI22xp5_ASAP7_75t_SL g16085 (.A1(n_6955),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_157),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_162),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_158),
    .Y(n_6957));
 INVx1_ASAP7_75t_SL g16086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_162),
    .Y(n_6955));
 XOR2xp5_ASAP7_75t_SL g16089 (.A(n_10482),
    .B(n_6961),
    .Y(n_6962));
 HB1xp67_ASAP7_75t_SL g16090 (.A(n_6958),
    .Y(n_6961));
 XOR2xp5_ASAP7_75t_SL g16091 (.A(n_6950),
    .B(n_6963),
    .Y(n_6964));
 XOR2xp5_ASAP7_75t_SL g16092 (.A(n_6954),
    .B(n_6957),
    .Y(n_6963));
 BUFx6f_ASAP7_75t_SL g16093 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[3]),
    .Y(n_6965));
 MAJIxp5_ASAP7_75t_SL g16094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_73),
    .B(n_19341),
    .C(n_6967),
    .Y(n_6968));
 NAND2xp5_ASAP7_75t_SL g16095 (.A(n_6972),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .Y(n_6967));
 INVx1_ASAP7_75t_SL g16099 (.A(n_6967),
    .Y(n_6969));
 BUFx3_ASAP7_75t_SL g16101 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[3]),
    .Y(n_6973));
 NAND3xp33_ASAP7_75t_SL g16103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_268),
    .B(n_6974),
    .C(n_6975),
    .Y(n_6976));
 NAND2xp5_ASAP7_75t_SL g16104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_238),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_241),
    .Y(n_6974));
 NAND2xp5_ASAP7_75t_SL g16105 (.A(n_9404),
    .B(n_6368),
    .Y(n_6975));
 NAND2xp5_ASAP7_75t_SL g16109 (.A(n_6984),
    .B(n_6987),
    .Y(n_6988));
 INVxp67_ASAP7_75t_SL g16110 (.A(n_6368),
    .Y(n_6985));
 INVxp33_ASAP7_75t_SRAM g16111 (.A(n_9404),
    .Y(n_6986));
 NAND2xp5_ASAP7_75t_SL g16112 (.A(n_6989),
    .B(n_6974),
    .Y(n_6991));
 OAI21xp5_ASAP7_75t_SL g16113 (.A1(n_6992),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_279),
    .B(n_6987),
    .Y(n_6993));
 XNOR2x1_ASAP7_75t_SL g16115 (.B(n_6996),
    .Y(n_6997),
    .A(n_6995));
 INVx1_ASAP7_75t_SL g16116 (.A(n_6994),
    .Y(n_6995));
 AND2x2_ASAP7_75t_SL g16117 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .Y(n_6994));
 AOI22xp5_ASAP7_75t_SL g16118 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_34),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_19),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_33),
    .Y(n_6996));
 XNOR2xp5_ASAP7_75t_SL g16119 (.A(n_6997),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_188),
    .Y(n_6999));
 MAJIxp5_ASAP7_75t_SL g16120 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_34),
    .B(n_6994),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_19),
    .Y(n_7000));
 NOR2x1_ASAP7_75t_SL g16121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_240),
    .B(n_7006),
    .Y(n_7007));
 XNOR2x2_ASAP7_75t_SL g16123 (.A(n_8090),
    .B(n_9106),
    .Y(n_7006));
 NAND2xp5_ASAP7_75t_SL g16127 (.A(n_7006),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_240),
    .Y(n_7008));
 MAJIxp5_ASAP7_75t_SL g16128 (.A(n_7009),
    .B(n_7010),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_208),
    .Y(n_7011));
 INVx1_ASAP7_75t_SL g16129 (.A(n_8090),
    .Y(n_7009));
 NAND2x1_ASAP7_75t_SL g16132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_268),
    .B(n_7014),
    .Y(n_7015));
 AND2x2_ASAP7_75t_SL g16133 (.A(n_7012),
    .B(n_7013),
    .Y(n_7014));
 NAND2xp5_ASAP7_75t_SL g16134 (.A(n_21956),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_229),
    .Y(n_7012));
 NAND2xp5_ASAP7_75t_SL g16135 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_238),
    .B(n_13551),
    .Y(n_7013));
 AOI21x1_ASAP7_75t_SL g16136 (.A1(n_7014),
    .A2(n_13975),
    .B(n_7020),
    .Y(n_7021));
 OAI21xp5_ASAP7_75t_SL g16138 (.A1(n_7017),
    .A2(n_7018),
    .B(n_7019),
    .Y(n_7020));
 OR2x2_ASAP7_75t_SL g16139 (.A(n_21956),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_229),
    .Y(n_7017));
 INVx1_ASAP7_75t_SL g16140 (.A(n_7013),
    .Y(n_7018));
 OR2x2_ASAP7_75t_SL g16141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_238),
    .B(n_13551),
    .Y(n_7019));
 AOI21x1_ASAP7_75t_SL g16143 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_268),
    .A2(n_4769),
    .B(n_13975),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_279));
 NAND2xp33_ASAP7_75t_R g16144 (.A(n_7012),
    .B(n_7017),
    .Y(n_7025));
 NAND2xp5_ASAP7_75t_SL g16145 (.A(n_7013),
    .B(n_7019),
    .Y(n_7027));
 OAI21xp5_ASAP7_75t_SL g16147 (.A1(n_7028),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_279),
    .B(n_7017),
    .Y(n_7029));
 INVxp33_ASAP7_75t_R g16148 (.A(n_7012),
    .Y(n_7028));
 OAI22x1_ASAP7_75t_SL g16158 (.A1(n_18648),
    .A2(n_21144),
    .B1(n_21146),
    .B2(n_7040),
    .Y(n_7041));
 NOR2x1_ASAP7_75t_SL g16165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_252),
    .B(n_7071),
    .Y(n_7072));
 XOR2x2_ASAP7_75t_SL g16166 (.A(n_21010),
    .B(n_20845),
    .Y(n_7071));
 NAND2xp5_ASAP7_75t_SL g16173 (.A(n_7071),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_252),
    .Y(n_7073));
 MAJx2_ASAP7_75t_SL g16175 (.A(n_21010),
    .B(n_19989),
    .C(n_6806),
    .Y(n_7075));
 AND2x2_ASAP7_75t_SL g16177 (.A(n_8838),
    .B(n_8836),
    .Y(n_7082));
 INVxp67_ASAP7_75t_SL g16182 (.A(n_7079),
    .Y(n_7080));
 NAND2xp5_ASAP7_75t_SL g16183 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .Y(n_7079));
 INVx1_ASAP7_75t_SL g16195 (.A(n_9065),
    .Y(n_7096));
 XNOR2xp5_ASAP7_75t_SL g16196 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_274),
    .B(n_7105),
    .Y(n_7106));
 OAI21xp5_ASAP7_75t_SL g16197 (.A1(n_7100),
    .A2(n_7101),
    .B(n_7104),
    .Y(n_7105));
 INVxp67_ASAP7_75t_SL g16198 (.A(n_7098),
    .Y(n_7099));
 NOR2xp33_ASAP7_75t_SL g16199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_249),
    .Y(n_7098));
 XNOR2xp5_ASAP7_75t_SL g162 (.A(n_21687),
    .B(n_14354),
    .Y(n_14355));
 INVxp67_ASAP7_75t_SL g16200 (.A(n_22430),
    .Y(n_7101));
 AOI21xp33_ASAP7_75t_SL g16201 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_313),
    .A2(n_7099),
    .B(n_7103),
    .Y(n_7104));
 INVxp67_ASAP7_75t_SL g16202 (.A(n_7102),
    .Y(n_7103));
 NAND2xp5_ASAP7_75t_SL g16203 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_255),
    .Y(n_7102));
 NOR2xp33_ASAP7_75t_SL g16204 (.A(n_7103),
    .B(n_7098),
    .Y(n_7107));
 NAND2xp5_ASAP7_75t_SL g16206 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_265),
    .B(n_7099),
    .Y(n_7109));
 OA21x2_ASAP7_75t_SL g16208 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_264),
    .A2(n_7102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_263),
    .Y(n_7111));
 XNOR2xp5_ASAP7_75t_SL g16209 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_12),
    .B(n_17712),
    .Y(n_7116));
 MAJIxp5_ASAP7_75t_SL g16213 (.A(n_17712),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_174),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_185),
    .Y(n_7117));
 INVx1_ASAP7_75t_SL g16220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_611),
    .Y(n_7121));
 INVx1_ASAP7_75t_SL g16227 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_178),
    .Y(n_7128));
 XNOR2xp5_ASAP7_75t_SL g16251 (.A(n_7171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_250),
    .Y(n_7172));
 HB1xp67_ASAP7_75t_SL g16252 (.A(n_7170),
    .Y(n_7171));
 OAI21xp5_ASAP7_75t_SL g16253 (.A1(n_7167),
    .A2(n_20913),
    .B(n_7169),
    .Y(n_7170));
 NOR2xp33_ASAP7_75t_SL g16254 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_188),
    .B(n_21462),
    .Y(n_7167));
 NAND2xp5_ASAP7_75t_SL g16256 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_188),
    .B(n_21462),
    .Y(n_7169));
 XOR2xp5_ASAP7_75t_SL g16259 (.A(n_20914),
    .B(n_19142),
    .Y(n_7179));
 MAJx2_ASAP7_75t_SL g16271 (.A(n_20865),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_191),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_193),
    .Y(n_7188));
 MAJIxp5_ASAP7_75t_SL g16273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_148),
    .C(n_19834),
    .Y(n_7189));
 HB1xp67_ASAP7_75t_SL g16275 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_219),
    .Y(n_7190));
 OAI22xp5_ASAP7_75t_SL g16276 (.A1(n_7194),
    .A2(n_7195),
    .B1(n_21351),
    .B2(n_7196),
    .Y(n_7197));
 INVx1_ASAP7_75t_SL g16277 (.A(n_21351),
    .Y(n_7194));
 XNOR2xp5_ASAP7_75t_SL g16281 (.A(n_7754),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_179),
    .Y(n_7195));
 INVx1_ASAP7_75t_SL g16282 (.A(n_7195),
    .Y(n_7196));
 OAI22xp5_ASAP7_75t_SL g16284 (.A1(n_7199),
    .A2(n_21351),
    .B1(n_7194),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_219),
    .Y(n_7200));
 INVx1_ASAP7_75t_SL g16285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_219),
    .Y(n_7199));
 XNOR2xp5_ASAP7_75t_SL g16299 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_124),
    .Y(n_7212));
 INVxp67_ASAP7_75t_SL g16300 (.A(n_7213),
    .Y(n_7214));
 MAJIxp5_ASAP7_75t_SL g16301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_103),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_78),
    .Y(n_7213));
 XNOR2xp5_ASAP7_75t_SL g16302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_20),
    .Y(n_7215));
 XOR2xp5_ASAP7_75t_SL g16305 (.A(n_7215),
    .B(n_7213),
    .Y(n_7222));
 MAJIxp5_ASAP7_75t_SL g16306 (.A(n_13294),
    .B(n_7553),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_185),
    .Y(n_7227));
 XNOR2xp5_ASAP7_75t_SL g16310 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_12),
    .B(n_13294),
    .Y(n_7228));
 INVxp67_ASAP7_75t_SL g16314 (.A(n_7236),
    .Y(n_7237));
 XOR2xp5_ASAP7_75t_SL g16315 (.A(n_7232),
    .B(n_7235),
    .Y(n_7236));
 INVxp67_ASAP7_75t_SL g16316 (.A(n_7231),
    .Y(n_7232));
 AND2x2_ASAP7_75t_SL g16317 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_53),
    .Y(n_7231));
 OAI22xp5_ASAP7_75t_SL g16318 (.A1(n_7233),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_80),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_89),
    .B2(n_7234),
    .Y(n_7235));
 INVx1_ASAP7_75t_SL g16319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_89),
    .Y(n_7233));
 INVx1_ASAP7_75t_SL g16320 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_80),
    .Y(n_7234));
 XNOR2xp5_ASAP7_75t_SL g16321 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_174),
    .B(n_7236),
    .Y(n_7239));
 XOR2x2_ASAP7_75t_SL g16333 (.A(n_18819),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_42),
    .Y(n_7249));
 XNOR2x2_ASAP7_75t_SL g16335 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_63),
    .B(n_21912),
    .Y(n_7250));
 MAJIxp5_ASAP7_75t_SL g16337 (.A(n_7249),
    .B(n_7250),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_155),
    .Y(n_7255));
 AND2x2_ASAP7_75t_SL g16340 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_4826),
    .Y(n_7256));
 NAND2xp5_ASAP7_75t_SL g16341 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .Y(n_7257));
 INVx1_ASAP7_75t_SL g16344 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_146));
 INVx1_ASAP7_75t_SL g16346 (.A(n_19144),
    .Y(n_7263));
 AOI21xp33_ASAP7_75t_SL g16347 (.A1(n_4826),
    .A2(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_7257),
    .Y(n_7265));
 AND2x2_ASAP7_75t_SL g16354 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(n_18031),
    .Y(n_7269));
 NAND2xp5_ASAP7_75t_SL g16357 (.A(n_22296),
    .B(n_10104),
    .Y(n_7282));
 NOR2xp67_ASAP7_75t_SL g16365 (.A(n_10104),
    .B(n_22296),
    .Y(n_7283));
 HB1xp67_ASAP7_75t_SL g16367 (.A(n_9634),
    .Y(n_7284));
 XNOR2x1_ASAP7_75t_SL g16386 (.B(n_14763),
    .Y(n_7309),
    .A(n_7307));
 MAJx2_ASAP7_75t_SL g16387 (.A(n_6880),
    .B(n_21963),
    .C(n_10803),
    .Y(n_7307));
 MAJIxp5_ASAP7_75t_SL g16389 (.A(n_14763),
    .B(n_7307),
    .C(n_12571),
    .Y(n_7311));
 XNOR2x1_ASAP7_75t_SL g16393 (.B(n_7317),
    .Y(n_7318),
    .A(n_7314));
 INVx1_ASAP7_75t_SL g16394 (.A(n_7313),
    .Y(n_7314));
 AND2x2_ASAP7_75t_SL g16395 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_53),
    .Y(n_7313));
 OAI22xp5_ASAP7_75t_SL g16396 (.A1(n_7315),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_80),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_89),
    .B2(n_7316),
    .Y(n_7317));
 INVx1_ASAP7_75t_SL g16397 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_80),
    .Y(n_7316));
 MAJIxp5_ASAP7_75t_SL g164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_81),
    .C(n_6279),
    .Y(n_6284));
 XOR2xp5_ASAP7_75t_SL g16402 (.A(n_7334),
    .B(n_10334),
    .Y(n_7332));
 NAND2xp5_ASAP7_75t_SL g16406 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(n_14183),
    .Y(n_7326));
 INVx1_ASAP7_75t_SL g16407 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_75),
    .Y(n_7327));
 AND2x2_ASAP7_75t_SL g16408 (.A(n_14179),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .Y(n_7328));
 INVxp67_ASAP7_75t_SL g16409 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_67),
    .Y(n_7330));
 MAJIxp5_ASAP7_75t_SL g16410 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_216),
    .B(n_7333),
    .C(n_7334),
    .Y(n_7335));
 HB1xp67_ASAP7_75t_SL g16411 (.A(n_10334),
    .Y(n_7333));
 MAJIxp5_ASAP7_75t_SL g16413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_75),
    .C(n_7326),
    .Y(n_7336));
 NOR2xp67_ASAP7_75t_SL g16418 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_258),
    .B(n_9841),
    .Y(n_7342));
 AOI21xp5_ASAP7_75t_SL g16419 (.A1(n_9840),
    .A2(n_20199),
    .B(n_20198),
    .Y(n_7343));
 AOI221xp5_ASAP7_75t_SL g16420 (.A1(n_18885),
    .A2(n_18886),
    .B1(n_7350),
    .B2(n_7351),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_119),
    .Y(n_7352));
 INVx2_ASAP7_75t_SL g16427 (.A(n_18885),
    .Y(n_7350));
 INVx1_ASAP7_75t_SL g16428 (.A(n_18886),
    .Y(n_7351));
 NAND2xp5_ASAP7_75t_SL g16429 (.A(n_7353),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_119),
    .Y(n_7354));
 OAI22xp5_ASAP7_75t_SL g16430 (.A1(n_18886),
    .A2(n_18885),
    .B1(n_7350),
    .B2(n_7351),
    .Y(n_7353));
 HB1xp67_ASAP7_75t_SL g16433 (.A(n_22631),
    .Y(n_7356));
 OAI21xp5_ASAP7_75t_SL g16434 (.A1(n_7360),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .B(n_7361),
    .Y(n_7362));
 NOR2xp67_ASAP7_75t_SL g16435 (.A(n_11544),
    .B(n_10393),
    .Y(n_7360));
 NAND2xp5_ASAP7_75t_SL g16437 (.A(n_11544),
    .B(n_10393),
    .Y(n_7361));
 NAND2xp5_ASAP7_75t_SL g16438 (.A(n_7361),
    .B(n_7363),
    .Y(n_7364));
 INVxp67_ASAP7_75t_SRAM g16439 (.A(n_7360),
    .Y(n_7363));
 XNOR2x2_ASAP7_75t_SL g16443 (.A(n_7381),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_6),
    .Y(n_7382));
 INVxp67_ASAP7_75t_SL g16444 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_65),
    .Y(n_7381));
 MAJIxp5_ASAP7_75t_SL g16445 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_75),
    .Y(n_7383));
 XNOR2xp5_ASAP7_75t_SL g16450 (.A(n_7382),
    .B(n_12934),
    .Y(n_7389));
 INVx1_ASAP7_75t_SL g16451 (.A(n_7383),
    .Y(n_7390));
 MAJx2_ASAP7_75t_SL g16455 (.A(n_7394),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_58),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_40),
    .Y(n_7397));
 INVx1_ASAP7_75t_SL g16456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_44),
    .Y(n_7394));
 INVx2_ASAP7_75t_SL g16457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_58));
 NOR2x1_ASAP7_75t_SL g16461 (.A(n_18738),
    .B(n_7406),
    .Y(n_7407));
 HB1xp67_ASAP7_75t_SL g16463 (.A(n_21439),
    .Y(n_7402));
 XNOR2xp5_ASAP7_75t_SL g16464 (.A(n_22896),
    .B(n_22055),
    .Y(n_7405));
 NAND2xp5_ASAP7_75t_SL g16465 (.A(n_7406),
    .B(n_18738),
    .Y(n_7408));
 MAJIxp5_ASAP7_75t_SL g16466 (.A(n_7409),
    .B(n_22896),
    .C(n_7403),
    .Y(n_7410));
 XOR2xp5_ASAP7_75t_SL g16499 (.A(n_7450),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_209),
    .Y(n_7451));
 XNOR2xp5_ASAP7_75t_SL g165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_81),
    .B(n_6279),
    .Y(n_6280));
 XNOR2xp5_ASAP7_75t_SL g16500 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_2),
    .B(n_18889),
    .Y(n_7450));
 NAND2xp5_ASAP7_75t_SL g16503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_121),
    .Y(n_7447));
 MAJIxp5_ASAP7_75t_SL g16505 (.A(n_7450),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_178),
    .C(n_6749),
    .Y(n_7452));
 MAJIxp5_ASAP7_75t_SL g16506 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_2),
    .B(n_7447),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_50),
    .Y(n_7453));
 OAI22xp33_ASAP7_75t_SL g16507 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_205),
    .A2(n_7457),
    .B1(n_7458),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_206),
    .Y(n_7459));
 XNOR2xp5_ASAP7_75t_SL g16508 (.A(n_7455),
    .B(n_7456),
    .Y(n_7457));
 INVxp67_ASAP7_75t_SL g16509 (.A(n_7454),
    .Y(n_7455));
 MAJIxp5_ASAP7_75t_SL g16510 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_103),
    .Y(n_7454));
 OAI22xp33_ASAP7_75t_SL g16511 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_117),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_4),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_149),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_118),
    .Y(n_7456));
 INVx1_ASAP7_75t_SL g16512 (.A(n_7457),
    .Y(n_7458));
 HB1xp67_ASAP7_75t_SL g16514 (.A(n_7457),
    .Y(n_7460));
 MAJIxp5_ASAP7_75t_SL g16515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_4),
    .B(n_7454),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_118),
    .Y(n_7462));
 XOR2xp5_ASAP7_75t_SL g16516 (.A(n_7898),
    .B(n_7468),
    .Y(n_7469));
 XOR2xp5_ASAP7_75t_SL g16517 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_67),
    .B(n_7467),
    .Y(n_7468));
 OAI22xp5_ASAP7_75t_SL g16518 (.A1(n_7463),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_75),
    .B1(n_7464),
    .B2(n_18739),
    .Y(n_7467));
 NAND2xp5_ASAP7_75t_SL g16519 (.A(n_22865),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .Y(n_7463));
 INVx1_ASAP7_75t_SL g16520 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_75),
    .Y(n_7464));
 MAJIxp5_ASAP7_75t_SL g16523 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_216),
    .B(n_7470),
    .C(n_7898),
    .Y(n_7471));
 HB1xp67_ASAP7_75t_SL g16524 (.A(n_7468),
    .Y(n_7470));
 NOR2x1p5_ASAP7_75t_SL g16526 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_180),
    .B(n_7477),
    .Y(n_7478));
 XNOR2x1_ASAP7_75t_SL g16527 (.B(n_7476),
    .Y(n_7477),
    .A(n_7474));
 XNOR2x1_ASAP7_75t_SL g16528 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_8),
    .Y(n_7474),
    .A(n_7473));
 INVx1_ASAP7_75t_SL g16529 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_106),
    .Y(n_7473));
 XNOR2x1_ASAP7_75t_SL g16530 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_147),
    .Y(n_7476),
    .A(n_18740));
 NAND2xp5_ASAP7_75t_SL g16532 (.A(n_7477),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_180),
    .Y(n_7479));
 INVx1_ASAP7_75t_SL g16534 (.A(n_7474),
    .Y(n_7480));
 HB1xp67_ASAP7_75t_SL g16535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_147),
    .Y(n_7481));
 INVxp67_ASAP7_75t_SL g16536 (.A(n_18740),
    .Y(n_7482));
 MAJIxp5_ASAP7_75t_SL g16538 (.A(n_7485),
    .B(n_13321),
    .C(n_7488),
    .Y(n_7489));
 XOR2x2_ASAP7_75t_SL g16539 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_11),
    .B(n_22257),
    .Y(n_7485));
 XNOR2x2_ASAP7_75t_SL g16542 (.A(n_7487),
    .B(n_19522),
    .Y(n_7488));
 NOR2x1_ASAP7_75t_SL g16543 (.A(n_7489),
    .B(n_11120),
    .Y(n_7491));
 XNOR2x1_ASAP7_75t_SL g16544 (.B(n_7492),
    .Y(n_7493),
    .A(n_7485));
 XNOR2x1_ASAP7_75t_SL g16545 (.B(n_13321),
    .Y(n_7492),
    .A(n_7488));
 NAND2xp5_ASAP7_75t_SL g16548 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_6973),
    .Y(n_7494));
 INVx1_ASAP7_75t_SL g16549 (.A(n_7495),
    .Y(n_7496));
 NAND2xp5_ASAP7_75t_SL g16550 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(n_7495));
 NAND2xp5_ASAP7_75t_SL g16551 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(n_2325),
    .Y(n_7497));
 XOR2xp5_ASAP7_75t_SL g16555 (.A(n_7494),
    .B(n_7497),
    .Y(n_7502));
 INVxp67_ASAP7_75t_SL g16560 (.A(n_7506),
    .Y(n_7507));
 OR2x2_ASAP7_75t_SL g16561 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_228),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_219),
    .Y(n_7506));
 NAND2xp5_ASAP7_75t_SL g16562 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_228),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_219),
    .Y(n_7508));
 INVxp67_ASAP7_75t_SL g16567 (.A(n_7514),
    .Y(n_7515));
 NOR2xp33_ASAP7_75t_SL g16568 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_232),
    .B(n_7507),
    .Y(n_7514));
 INVxp67_ASAP7_75t_SL g16569 (.A(n_7516),
    .Y(n_7517));
 OAI21xp33_ASAP7_75t_SL g16570 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_232),
    .A2(n_7508),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_236),
    .Y(n_7516));
 XOR2xp5_ASAP7_75t_SL g16573 (.A(n_7521),
    .B(n_20689),
    .Y(n_7523));
 XNOR2xp5_ASAP7_75t_SL g16574 (.A(n_7520),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_11),
    .Y(n_7521));
 HB1xp67_ASAP7_75t_SL g16575 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_32),
    .Y(n_7520));
 NOR2xp33_ASAP7_75t_SL g16578 (.A(n_7521),
    .B(n_20689),
    .Y(n_7526));
 NAND2xp33_ASAP7_75t_L g16579 (.A(n_20689),
    .B(n_7521),
    .Y(n_7527));
 NOR2xp67_ASAP7_75t_SL g16580 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_260),
    .B(n_7543),
    .Y(n_7531));
 NOR2xp33_ASAP7_75t_SL g16586 (.A(n_7539),
    .B(n_5277),
    .Y(n_7540));
 MAJIxp5_ASAP7_75t_SL g16587 (.A(n_7534),
    .B(n_7536),
    .C(n_7538),
    .Y(n_7539));
 XOR2xp5_ASAP7_75t_SL g16589 (.A(n_7534),
    .B(n_7542),
    .Y(n_7543));
 AND2x2_ASAP7_75t_SL g16594 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_121),
    .Y(n_7544));
 OAI22xp5_ASAP7_75t_SL g16595 (.A1(n_7546),
    .A2(n_13538),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_50),
    .B2(n_7547),
    .Y(n_7548));
 INVx1_ASAP7_75t_SL g16596 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_50),
    .Y(n_7546));
 INVx1_ASAP7_75t_SL g16597 (.A(n_13538),
    .Y(n_7547));
 MAJx2_ASAP7_75t_SL g16599 (.A(n_7547),
    .B(n_7546),
    .C(n_7544),
    .Y(n_7553));
 AND2x2_ASAP7_75t_SL g16602 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(n_3713),
    .Y(n_7558));
 MAJIxp5_ASAP7_75t_SL g16605 (.A(n_7571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_135),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_121),
    .Y(n_7572));
 XNOR2x1_ASAP7_75t_SL g16607 (.B(n_7569),
    .Y(n_7570),
    .A(n_7565));
 NAND2xp5_ASAP7_75t_SL g16608 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(n_14186),
    .Y(n_7565));
 OAI22x1_ASAP7_75t_SL g16609 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_87),
    .A2(n_7566),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_88),
    .B2(n_7568),
    .Y(n_7569));
 INVxp67_ASAP7_75t_SL g16610 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_104),
    .Y(n_7566));
 INVx2_ASAP7_75t_SL g16611 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_88));
 BUFx2_ASAP7_75t_SL g16612 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_104),
    .Y(n_7568));
 XNOR2x1_ASAP7_75t_SL g16613 (.B(n_7570),
    .Y(n_7573),
    .A(n_6635));
 MAJIxp5_ASAP7_75t_SL g16614 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_88),
    .B(n_7568),
    .C(n_7565),
    .Y(n_7334));
 XNOR2xp5_ASAP7_75t_SL g16616 (.A(n_7575),
    .B(n_7576),
    .Y(n_7577));
 XNOR2xp5_ASAP7_75t_SL g16617 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_4),
    .Y(n_7575));
 AOI22xp5_ASAP7_75t_SL g16618 (.A1(n_11090),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_140),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_156),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_3),
    .Y(n_7576));
 XNOR2xp5_ASAP7_75t_SL g16619 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_12),
    .B(n_7577),
    .Y(n_7579));
 OAI21xp5_ASAP7_75t_SL g16621 (.A1(n_7587),
    .A2(n_13640),
    .B(n_13641),
    .Y(n_7588));
 MAJIxp5_ASAP7_75t_SL g16622 (.A(n_7581),
    .B(n_7585),
    .C(n_7586),
    .Y(n_7587));
 OAI21xp5_ASAP7_75t_SL g16623 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_174),
    .Y(n_7581));
 MAJIxp5_ASAP7_75t_SL g16624 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_116),
    .B(n_7583),
    .C(n_7584),
    .Y(n_7585));
 HB1xp67_ASAP7_75t_SL g16626 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_35),
    .Y(n_7583));
 XNOR2xp5_ASAP7_75t_SL g16627 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_151),
    .Y(n_7586));
 XOR2xp5_ASAP7_75t_SL g16629 (.A(n_7590),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_231),
    .Y(n_7591));
 HB1xp67_ASAP7_75t_SL g16630 (.A(n_7587),
    .Y(n_7590));
 XOR2xp5_ASAP7_75t_SL g16631 (.A(n_7592),
    .B(n_7581),
    .Y(n_7593));
 XOR2xp5_ASAP7_75t_SL g16632 (.A(n_7585),
    .B(n_7586),
    .Y(n_7592));
 AND3x2_ASAP7_75t_SL g16634 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[4]),
    .Y(n_7595));
 OAI21x1_ASAP7_75t_SL g16636 (.A1(n_7596),
    .A2(n_7597),
    .B(n_7595),
    .Y(n_7598));
 AND2x2_ASAP7_75t_SL g16637 (.A(n_8180),
    .B(n_8298),
    .Y(n_7596));
 NOR2xp67_ASAP7_75t_SL g16638 (.A(n_8180),
    .B(n_8298),
    .Y(n_7597));
 OA21x2_ASAP7_75t_SL g16641 (.A1(n_7597),
    .A2(n_7596),
    .B(n_7595),
    .Y(n_7601));
 INVx1_ASAP7_75t_SL g16644 (.A(n_6836),
    .Y(n_7604));
 XOR2xp5_ASAP7_75t_SL g16645 (.A(n_18891),
    .B(n_7609),
    .Y(n_7610));
 INVx1_ASAP7_75t_SL g16649 (.A(n_7608),
    .Y(n_7609));
 OAI21xp5_ASAP7_75t_SL g16650 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .A2(n_11105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(n_7608));
 INVx1_ASAP7_75t_SL g16655 (.A(n_20124),
    .Y(n_7615));
 NOR2xp33_ASAP7_75t_SL g16673 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_257),
    .B(n_19532),
    .Y(n_7637));
 INVx2_ASAP7_75t_SL g16674 (.A(n_19531),
    .Y(n_7638));
 OAI21xp5_ASAP7_75t_SL g16680 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_257),
    .A2(n_19534),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_260),
    .Y(n_7644));
 XNOR2x1_ASAP7_75t_SL g16692 (.B(n_7656),
    .Y(n_7657),
    .A(n_7655));
 NAND2x1_ASAP7_75t_L g16693 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(n_3214),
    .Y(n_7655));
 NAND2xp5_ASAP7_75t_SL g16694 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .Y(n_7656));
 XNOR2x1_ASAP7_75t_SL g16699 (.B(n_19796),
    .Y(n_7665),
    .A(n_7661));
 OAI21xp5_ASAP7_75t_SL g167 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_51),
    .A2(n_22954),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .Y(n_9908));
 AO22x1_ASAP7_75t_SL g16700 (.A1(n_4965),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_22),
    .B1(n_20878),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_153),
    .Y(n_7661));
 MAJx2_ASAP7_75t_SL g16705 (.A(n_21036),
    .B(n_7669),
    .C(n_3915),
    .Y(n_7670));
 INVxp67_ASAP7_75t_SL g16706 (.A(n_7665),
    .Y(n_7669));
 NOR2xp33_ASAP7_75t_SL g16710 (.A(n_19146),
    .B(n_7675),
    .Y(n_7676));
 XNOR2xp5_ASAP7_75t_SL g16713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_137),
    .Y(n_7675));
 NAND2xp5_ASAP7_75t_SL g16714 (.A(n_19146),
    .B(n_7675),
    .Y(n_7677));
 AO22x1_ASAP7_75t_SL g16719 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_34),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_33),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_19),
    .Y(n_7681));
 AND2x2_ASAP7_75t_SL g16720 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32),
    .Y(n_7682));
 XNOR2xp5_ASAP7_75t_SL g16721 (.A(n_19358),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_188),
    .Y(n_7685));
 MAJIxp5_ASAP7_75t_SL g16722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_34),
    .B(n_7682),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_19),
    .Y(n_7686));
 NAND2xp5_ASAP7_75t_SL g16736 (.A(n_10774),
    .B(n_19605),
    .Y(n_7697));
 NAND2xp5_ASAP7_75t_SL g16737 (.A(n_9614),
    .B(n_19909),
    .Y(n_7698));
 AOI21x1_ASAP7_75t_SL g16738 (.A1(n_7702),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_319),
    .B(n_6107),
    .Y(n_7703));
 INVxp67_ASAP7_75t_SL g16739 (.A(n_12892),
    .Y(n_7702));
 AND2x2_ASAP7_75t_SRAM g16740 (.A(n_7697),
    .B(n_6109),
    .Y(n_7704));
 AOI21xp5_ASAP7_75t_SL g16741 (.A1(n_9616),
    .A2(n_7697),
    .B(n_18820),
    .Y(n_7705));
 OAI21xp5_ASAP7_75t_SL g16742 (.A1(n_7707),
    .A2(n_7703),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_307),
    .Y(n_7708));
 INVxp67_ASAP7_75t_SL g16743 (.A(n_7706),
    .Y(n_7707));
 HB1xp67_ASAP7_75t_SL g16744 (.A(n_7698),
    .Y(n_7706));
 NAND2xp5_ASAP7_75t_SL g16745 (.A(n_7706),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_307),
    .Y(n_7709));
 XOR2x2_ASAP7_75t_SL g16748 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_277),
    .B(n_10274),
    .Y(n_7710));
 NOR2x1p5_ASAP7_75t_SL g16752 (.A(n_10395),
    .B(n_23092),
    .Y(n_7716));
 XNOR2x1_ASAP7_75t_SL g16756 (.B(n_7720),
    .Y(n_7721),
    .A(n_7719));
 NAND2xp5_ASAP7_75t_SL g16757 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(n_3275),
    .Y(n_7719));
 XNOR2x2_ASAP7_75t_SL g16758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_65),
    .Y(n_7720));
 MAJIxp5_ASAP7_75t_SL g16762 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_78),
    .C(n_7719),
    .Y(n_7726));
 MAJx2_ASAP7_75t_SL g16763 (.A(n_9143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_29),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_9),
    .Y(n_7727));
 XNOR2xp5_ASAP7_75t_SL g16773 (.A(n_7742),
    .B(n_21205),
    .Y(n_7746));
 INVxp67_ASAP7_75t_SL g16774 (.A(n_21061),
    .Y(n_7742));
 AOI21xp5_ASAP7_75t_SL g16779 (.A1(n_7748),
    .A2(n_7527),
    .B(n_7526),
    .Y(n_7749));
 INVx1_ASAP7_75t_SL g16780 (.A(n_7746),
    .Y(n_7748));
 MAJIxp5_ASAP7_75t_SL g16783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_80),
    .B(n_20510),
    .C(n_7753),
    .Y(n_7754));
 NAND2xp5_ASAP7_75t_R g16784 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .Y(n_7753));
 INVxp67_ASAP7_75t_SL g168 (.A(n_9905),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_51));
 OAI21xp5_ASAP7_75t_SL g16805 (.A1(n_7782),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_285),
    .B(n_5047),
    .Y(n_7783));
 INVx1_ASAP7_75t_SL g16806 (.A(n_7781),
    .Y(n_7782));
 OAI21x1_ASAP7_75t_SL g16807 (.A1(n_7776),
    .A2(n_7779),
    .B(n_7780),
    .Y(n_7781));
 INVx2_ASAP7_75t_SL g16808 (.A(n_7775),
    .Y(n_7776));
 AO21x2_ASAP7_75t_SL g16809 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_266),
    .A2(n_13655),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_264),
    .Y(n_7775));
 INVx1_ASAP7_75t_SL g16810 (.A(n_7778),
    .Y(n_7779));
 HB1xp67_ASAP7_75t_SL g16811 (.A(n_7227),
    .Y(n_7777));
 XNOR2xp5_ASAP7_75t_SL g16813 (.A(n_7786),
    .B(n_7787),
    .Y(n_7788));
 INVxp67_ASAP7_75t_SL g16814 (.A(n_7776),
    .Y(n_7786));
 NAND2xp5_ASAP7_75t_SL g16815 (.A(n_7778),
    .B(n_7780),
    .Y(n_7787));
 XNOR2xp5_ASAP7_75t_SL g16822 (.A(n_7798),
    .B(n_7799),
    .Y(n_7800));
 NAND2xp5_ASAP7_75t_SL g16823 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(n_7798));
 NOR2x1_ASAP7_75t_SL g16824 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_43),
    .B(n_3107),
    .Y(n_7799));
 INVx1_ASAP7_75t_SL g16825 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_126),
    .Y(n_7801));
 AO21x1_ASAP7_75t_SL g16826 (.A1(n_7803),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_126),
    .B(n_7804),
    .Y(n_7805));
 NAND2xp33_ASAP7_75t_SL g16827 (.A(n_7799),
    .B(n_7798),
    .Y(n_7803));
 NOR2xp33_ASAP7_75t_SL g16828 (.A(n_7798),
    .B(n_7799),
    .Y(n_7804));
 XNOR2x1_ASAP7_75t_SL g16841 (.B(n_7820),
    .Y(n_7821),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_709));
 XNOR2x1_ASAP7_75t_SL g16842 (.B(n_7819),
    .Y(n_7820),
    .A(n_14339));
 AND2x2_ASAP7_75t_SL g16844 (.A(n_2163),
    .B(n_21662),
    .Y(n_7819));
 NOR2xp67_ASAP7_75t_SL g16870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_217),
    .B(n_7854),
    .Y(n_7855));
 XOR2x2_ASAP7_75t_SL g16871 (.A(n_13332),
    .B(n_21796),
    .Y(n_7854));
 NAND2xp5_ASAP7_75t_SL g16879 (.A(n_7854),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_217),
    .Y(n_7858));
 INVx1_ASAP7_75t_SL g16881 (.A(n_13332),
    .Y(n_7859));
 NAND2xp5_ASAP7_75t_SL g16885 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .Y(n_7862));
 AND2x2_ASAP7_75t_SL g16886 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(n_7863));
 XNOR2xp5_ASAP7_75t_SL g16889 (.A(n_13767),
    .B(n_7868),
    .Y(n_7869));
 NAND2xp33_ASAP7_75t_SL g16891 (.A(n_14674),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .Y(n_7868));
 OAI21xp5_ASAP7_75t_SL g16892 (.A1(n_6569),
    .A2(n_7872),
    .B(n_7873),
    .Y(n_7874));
 NOR2xp33_ASAP7_75t_SL g16893 (.A(n_13767),
    .B(n_7871),
    .Y(n_7872));
 NAND2xp5_ASAP7_75t_SL g16894 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(n_14674),
    .Y(n_7871));
 NAND2xp5_ASAP7_75t_SL g16895 (.A(n_13767),
    .B(n_7871),
    .Y(n_7873));
 MAJx2_ASAP7_75t_SL g16898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_207),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_156),
    .C(n_21679),
    .Y(n_7876));
 XNOR2xp5_ASAP7_75t_SL g169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_111),
    .B(n_5841),
    .Y(n_5842));
 AOI22xp5_ASAP7_75t_SL g16900 (.A1(n_7877),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_239),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_238),
    .B2(n_10307),
    .Y(n_7879));
 INVx1_ASAP7_75t_SL g16901 (.A(n_10307),
    .Y(n_7877));
 MAJx2_ASAP7_75t_SL g16905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_239),
    .B(n_7876),
    .C(n_10307),
    .Y(n_7884));
 INVxp67_ASAP7_75t_SL g16908 (.A(n_7885),
    .Y(n_7886));
 NOR2xp33_ASAP7_75t_SL g16909 (.A(n_14372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_46),
    .Y(n_7885));
 NAND2xp5_ASAP7_75t_SL g16916 (.A(n_3468),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .Y(n_7893));
 NAND2xp5_ASAP7_75t_SL g16918 (.A(n_2927),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .Y(n_7894));
 MAJIxp5_ASAP7_75t_SL g16919 (.A(n_6523),
    .B(n_7894),
    .C(n_22997),
    .Y(n_7898));
 OAI21xp5_ASAP7_75t_SL g16924 (.A1(n_9904),
    .A2(n_7904),
    .B(n_7905),
    .Y(n_7906));
 OR2x2_ASAP7_75t_SL g16925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_264),
    .B(n_9896),
    .Y(n_7904));
 OA21x2_ASAP7_75t_SL g16926 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_264),
    .A2(n_9900),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_263),
    .Y(n_7905));
 NOR2xp33_ASAP7_75t_SL g16928 (.A(n_7908),
    .B(n_9896),
    .Y(n_7909));
 INVx1_ASAP7_75t_SL g16929 (.A(n_9900),
    .Y(n_7908));
 MAJx2_ASAP7_75t_SL g16945 (.A(n_7925),
    .B(n_3907),
    .C(n_7926),
    .Y(n_7927));
 NAND2xp5_ASAP7_75t_SL g16955 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_610),
    .B(n_2179),
    .Y(n_7932));
 INVx1_ASAP7_75t_SL g16959 (.A(n_7932),
    .Y(n_7938));
 NAND2xp5_ASAP7_75t_SL g16961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_258),
    .B(n_23169),
    .Y(n_7947));
 XNOR2xp5_ASAP7_75t_SL g16983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_6),
    .Y(n_7963));
 INVx1_ASAP7_75t_SL g16985 (.A(n_24754),
    .Y(n_7964));
 INVx1_ASAP7_75t_SL g16986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154),
    .Y(n_7965));
 OAI22xp33_ASAP7_75t_SL g16988 (.A1(n_7973),
    .A2(n_2848),
    .B1(n_7963),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154),
    .Y(n_7974));
 AND3x1_ASAP7_75t_SL g16989 (.A(n_7971),
    .B(n_7972),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154),
    .Y(n_7973));
 OR2x2_ASAP7_75t_SL g16990 (.A(n_7970),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_6),
    .Y(n_7971));
 INVx1_ASAP7_75t_SL g16991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_119),
    .Y(n_7970));
 NAND2xp33_ASAP7_75t_SL g16992 (.A(n_7970),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_6),
    .Y(n_7972));
 OAI21xp5_ASAP7_75t_SL g16993 (.A1(n_6784),
    .A2(n_7979),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_307),
    .Y(n_7980));
 INVx1_ASAP7_75t_SL g16994 (.A(n_11241),
    .Y(n_7979));
 NAND2xp5_ASAP7_75t_SL g16999 (.A(n_7979),
    .B(n_5794),
    .Y(n_7981));
 XOR2xp5_ASAP7_75t_SL g17 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_8),
    .Y(n_25921));
 OAI22xp5_ASAP7_75t_SL g170 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_69),
    .A2(n_13724),
    .B1(n_4026),
    .B2(n_5840),
    .Y(n_5841));
 XNOR2x1_ASAP7_75t_SL g17007 (.B(n_7399),
    .Y(n_7994),
    .A(n_7992));
 XOR2xp5_ASAP7_75t_SL g17008 (.A(n_7990),
    .B(n_7991),
    .Y(n_7992));
 MAJx2_ASAP7_75t_SL g17009 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_65),
    .B(n_7655),
    .C(n_7656),
    .Y(n_7991));
 INVx1_ASAP7_75t_SL g17010 (.A(n_7397),
    .Y(n_7399));
 INVxp67_ASAP7_75t_SL g17012 (.A(n_7991),
    .Y(n_7996));
 HB1xp67_ASAP7_75t_SL g17013 (.A(n_7990),
    .Y(n_7997));
 XNOR2xp5_ASAP7_75t_SL g17015 (.A(n_8000),
    .B(n_8002),
    .Y(n_8003));
 INVx1_ASAP7_75t_SL g17016 (.A(n_7999),
    .Y(n_8000));
 MAJIxp5_ASAP7_75t_SL g17017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_45),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_95),
    .C(n_14725),
    .Y(n_7999));
 XOR2xp5_ASAP7_75t_SL g17018 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_123),
    .B(n_8001),
    .Y(n_8002));
 INVx1_ASAP7_75t_SL g17019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_98),
    .Y(n_8001));
 MAJIxp5_ASAP7_75t_SL g17020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_171),
    .B(n_7999),
    .C(n_8005),
    .Y(n_8006));
 HB1xp67_ASAP7_75t_SL g17021 (.A(n_8002),
    .Y(n_8005));
 AND2x2_ASAP7_75t_SL g17026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_98),
    .Y(n_8007));
 OR2x2_ASAP7_75t_SL g17030 (.A(n_16557),
    .B(n_9182),
    .Y(n_8014));
 XNOR2xp5_ASAP7_75t_SL g17031 (.A(n_9182),
    .B(n_16557),
    .Y(n_8016));
 OAI21x1_ASAP7_75t_SL g17032 (.A1(n_8017),
    .A2(n_8007),
    .B(n_8018),
    .Y(n_8019));
 NOR2xp33_ASAP7_75t_SL g17033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_73),
    .Y(n_8017));
 NAND2xp5_ASAP7_75t_SL g17034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_73),
    .Y(n_8018));
 INVxp67_ASAP7_75t_SL g17040 (.A(n_19143),
    .Y(n_8022));
 HB1xp67_ASAP7_75t_SL g17043 (.A(n_8862),
    .Y(n_8027));
 XNOR2x1_ASAP7_75t_SL g17046 (.B(n_8031),
    .Y(n_8032),
    .A(n_8030));
 NAND2x1_ASAP7_75t_SL g17047 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(n_2335),
    .Y(n_8030));
 AND2x2_ASAP7_75t_SL g17048 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .B(n_6972),
    .Y(n_8031));
 MAJIxp5_ASAP7_75t_SL g17050 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_27),
    .B(n_8030),
    .C(n_8031),
    .Y(n_8035));
 MAJx2_ASAP7_75t_SL g17067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_705),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_769),
    .C(n_21519),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117));
 AOI22xp5_ASAP7_75t_SL g17070 (.A1(n_18157),
    .A2(n_8053),
    .B1(n_9246),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .Y(n_8057));
 XOR2xp5_ASAP7_75t_SL g17079 (.A(n_8067),
    .B(n_8068),
    .Y(n_8069));
 XNOR2xp5_ASAP7_75t_SL g17080 (.A(n_8066),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_8),
    .Y(n_8067));
 INVx1_ASAP7_75t_SL g17081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_156),
    .Y(n_8066));
 MAJIxp5_ASAP7_75t_SL g17082 (.A(n_7212),
    .B(n_7214),
    .C(n_7215),
    .Y(n_8068));
 XNOR2x1_ASAP7_75t_SL g17098 (.B(n_8089),
    .Y(n_8090),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_158));
 XOR2x1_ASAP7_75t_SL g17099 (.A(n_23403),
    .Y(n_8089),
    .B(n_8088));
 INVxp67_ASAP7_75t_SL g171 (.A(n_13724),
    .Y(n_5840));
 XNOR2x2_ASAP7_75t_SL g17102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_6),
    .Y(n_8088));
 INVxp67_ASAP7_75t_SL g17103 (.A(n_8091),
    .Y(n_8092));
 MAJIxp5_ASAP7_75t_SL g17104 (.A(n_23403),
    .B(n_8088),
    .C(n_4951),
    .Y(n_8091));
 MAJIxp5_ASAP7_75t_SL g17124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_17),
    .B(n_9750),
    .C(n_8130),
    .Y(n_8131));
 INVx1_ASAP7_75t_SL g17125 (.A(n_8129),
    .Y(n_8130));
 XNOR2xp5_ASAP7_75t_SL g17126 (.A(n_8125),
    .B(n_18901),
    .Y(n_8129));
 NAND2xp5_ASAP7_75t_SL g17127 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_6965),
    .Y(n_8125));
 MAJIxp5_ASAP7_75t_SL g17133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_71),
    .C(n_8125),
    .Y(n_8134));
 INVx1_ASAP7_75t_SL g17136 (.A(n_13596),
    .Y(n_8137));
 INVx1_ASAP7_75t_SL g17138 (.A(n_21971),
    .Y(n_8135));
 MAJIxp5_ASAP7_75t_SL g17139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_188),
    .B(n_22594),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_115),
    .Y(n_8140));
 INVx1_ASAP7_75t_SL g17142 (.A(n_8140),
    .Y(n_8141));
 MAJIxp5_ASAP7_75t_SL g17143 (.A(n_13596),
    .B(n_8141),
    .C(n_8144),
    .Y(n_8145));
 INVx1_ASAP7_75t_SL g17144 (.A(n_21686),
    .Y(n_8144));
 XNOR2xp5_ASAP7_75t_SL g17146 (.A(n_8146),
    .B(n_19646),
    .Y(n_8148));
 NAND2x1_ASAP7_75t_SL g17147 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_14987),
    .Y(n_8146));
 MAJIxp5_ASAP7_75t_SL g17149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_91),
    .B(n_19646),
    .C(n_8146),
    .Y(n_8150));
 NOR2x1_ASAP7_75t_SL g17157 (.A(n_11021),
    .B(n_8158),
    .Y(n_8159));
 XNOR2x1_ASAP7_75t_SL g17159 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_221),
    .Y(n_8158),
    .A(n_22123));
 NOR2xp67_ASAP7_75t_SL g17160 (.A(n_8159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_262),
    .Y(n_8161));
 INVxp67_ASAP7_75t_SL g17168 (.A(n_8166),
    .Y(n_8167));
 AND2x2_ASAP7_75t_SL g17171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_247),
    .Y(n_8170));
 INVx1_ASAP7_75t_SL g17172 (.A(n_8299),
    .Y(n_8178));
 NOR2xp33_ASAP7_75t_SL g17174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_262),
    .B(n_8166),
    .Y(n_8174));
 OAI21xp5_ASAP7_75t_SL g17175 (.A1(n_8175),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_262),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_261),
    .Y(n_8176));
 INVx1_ASAP7_75t_SL g17176 (.A(n_8170),
    .Y(n_8175));
 NOR2xp33_ASAP7_75t_SL g17178 (.A(n_8170),
    .B(n_8166),
    .Y(n_8180));
 XNOR2xp5_ASAP7_75t_SL g17179 (.A(n_9756),
    .B(n_10376),
    .Y(n_8185));
 XNOR2xp5_ASAP7_75t_SL g17185 (.A(n_9751),
    .B(n_8187),
    .Y(n_8188));
 XOR2xp5_ASAP7_75t_SL g17186 (.A(n_9753),
    .B(n_9752),
    .Y(n_8187));
 INVxp67_ASAP7_75t_SL g17191 (.A(n_19600),
    .Y(n_8194));
 MAJIxp5_ASAP7_75t_SL g172 (.A(n_19623),
    .B(n_3827),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_88),
    .Y(n_10029));
 MAJIxp5_ASAP7_75t_SL g17204 (.A(n_22949),
    .B(n_8213),
    .C(n_14106),
    .Y(n_8214));
 MAJIxp5_ASAP7_75t_SL g17215 (.A(n_8227),
    .B(n_8225),
    .C(n_8224),
    .Y(n_8228));
 NAND2x1_ASAP7_75t_SL g17216 (.A(n_2335),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .Y(n_8224));
 NAND2x1_ASAP7_75t_SL g17217 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .B(n_6973),
    .Y(n_8225));
 INVx1_ASAP7_75t_SL g17218 (.A(n_8226),
    .Y(n_8227));
 NAND2xp5_ASAP7_75t_SL g17219 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .Y(n_8226));
 XOR2xp5_ASAP7_75t_SL g17222 (.A(n_8226),
    .B(n_8232),
    .Y(n_8233));
 XNOR2xp5_ASAP7_75t_SL g17223 (.A(n_8225),
    .B(n_8224),
    .Y(n_8232));
 MAJx2_ASAP7_75t_SL g17225 (.A(n_8235),
    .B(n_8238),
    .C(n_8240),
    .Y(n_8241));
 NAND2xp5_ASAP7_75t_SL g17226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_748),
    .B(n_2154),
    .Y(n_8235));
 INVxp67_ASAP7_75t_SL g17228 (.A(n_8237),
    .Y(n_8238));
 INVx2_ASAP7_75t_SL g17229 (.A(n_9925),
    .Y(n_8237));
 NAND2x1p5_ASAP7_75t_SL g17231 (.A(n_8239),
    .B(n_11970),
    .Y(n_8240));
 HB1xp67_ASAP7_75t_SL g17232 (.A(n_2165),
    .Y(n_8239));
 AOI22x1_ASAP7_75t_SL g17235 (.A1(n_8244),
    .A2(n_8237),
    .B1(n_8240),
    .B2(n_9925),
    .Y(n_8245));
 INVx1_ASAP7_75t_SL g17236 (.A(n_8240),
    .Y(n_8244));
 MAJIxp5_ASAP7_75t_SL g17238 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_159),
    .C(n_11200),
    .Y(n_8248));
 NAND2xp5_ASAP7_75t_SL g17247 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(n_8255));
 NAND2xp5_ASAP7_75t_SL g17248 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(n_2325),
    .Y(n_8256));
 MAJIxp5_ASAP7_75t_SL g17249 (.A(n_9545),
    .B(n_8259),
    .C(n_8256),
    .Y(n_8260));
 INVx1_ASAP7_75t_SL g17250 (.A(n_8255),
    .Y(n_8259));
 NAND2xp5_ASAP7_75t_SL g17251 (.A(n_13126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_180),
    .Y(n_8265));
 OAI22xp5_ASAP7_75t_SL g17253 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_135),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_120),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_134),
    .Y(n_8261));
 NAND3xp33_ASAP7_75t_SL g17279 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_268),
    .B(n_15173),
    .C(n_15187),
    .Y(n_8290));
 AND2x2_ASAP7_75t_SL g17283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_302),
    .B(n_12272),
    .Y(n_8292));
 AOI21xp5_ASAP7_75t_SL g17284 (.A1(n_8167),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_311),
    .B(n_8170),
    .Y(n_8295));
 AOI21xp33_ASAP7_75t_SL g17285 (.A1(n_8292),
    .A2(n_13363),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_311),
    .Y(n_8298));
 A2O1A1O1Ixp25_ASAP7_75t_SL g17286 (.A1(n_13363),
    .A2(n_8292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_311),
    .C(n_8174),
    .D(n_8176),
    .Y(n_8299));
 OAI21xp5_ASAP7_75t_SL g17287 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_252),
    .A2(n_8303),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_254),
    .Y(n_8304));
 AOI21xp5_ASAP7_75t_SL g17288 (.A1(n_8300),
    .A2(n_10796),
    .B(n_8302),
    .Y(n_8303));
 NAND2xp5_ASAP7_75t_SL g17289 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_214),
    .Y(n_8300));
 NOR2xp33_ASAP7_75t_SL g17291 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_214),
    .Y(n_8302));
 XOR2xp5_ASAP7_75t_SL g17292 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_262),
    .B(n_8305),
    .Y(n_8306));
 HB1xp67_ASAP7_75t_SL g17293 (.A(n_8303),
    .Y(n_8305));
 XNOR2xp5_ASAP7_75t_SL g17294 (.A(n_10797),
    .B(n_8310),
    .Y(n_8311));
 NAND2xp5_ASAP7_75t_SL g17295 (.A(n_8300),
    .B(n_8309),
    .Y(n_8310));
 NAND2xp5_ASAP7_75t_SL g17296 (.A(n_8307),
    .B(n_8308),
    .Y(n_8309));
 INVx1_ASAP7_75t_SL g17297 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_181),
    .Y(n_8307));
 INVxp67_ASAP7_75t_SRAM g17298 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_214),
    .Y(n_8308));
 NAND2xp5_ASAP7_75t_SL g173 (.A(n_12748),
    .B(n_7638),
    .Y(n_22287));
 INVxp67_ASAP7_75t_SL g17301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_100),
    .Y(n_8312));
 INVx1_ASAP7_75t_SL g17305 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_54),
    .Y(n_8315));
 AND2x2_ASAP7_75t_SL g17309 (.A(n_22218),
    .B(n_22216),
    .Y(n_8321));
 OAI21xp5_ASAP7_75t_SL g17311 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_23),
    .A2(n_13247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_27),
    .Y(n_8322));
 INVx1_ASAP7_75t_SL g17314 (.A(n_17486),
    .Y(n_8329));
 AOI221xp5_ASAP7_75t_SL g17329 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_187),
    .A2(n_26046),
    .B1(n_8344),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_188),
    .C(n_8346),
    .Y(n_8347));
 INVx1_ASAP7_75t_SL g17330 (.A(n_26046),
    .Y(n_8344));
 MAJIxp5_ASAP7_75t_SL g17331 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_115),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_108),
    .Y(n_8346));
 NAND2xp5_ASAP7_75t_SL g17332 (.A(n_8348),
    .B(n_8346),
    .Y(n_8349));
 NAND2xp5_ASAP7_75t_SL g17334 (.A(n_8349),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_222),
    .Y(n_8352));
 AOI22xp33_ASAP7_75t_SL g17346 (.A1(n_19729),
    .A2(n_8367),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_270),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_274),
    .Y(n_8368));
 NOR2xp67_ASAP7_75t_SL g17347 (.A(n_8365),
    .B(n_12666),
    .Y(n_8367));
 MAJIxp5_ASAP7_75t_SL g17348 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_234),
    .B(n_2962),
    .C(n_3552),
    .Y(n_8365));
 INVxp67_ASAP7_75t_SL g17351 (.A(n_8367),
    .Y(n_8369));
 XNOR2xp5_ASAP7_75t_SL g17354 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_148),
    .B(n_8375),
    .Y(n_8376));
 XOR2xp5_ASAP7_75t_SL g17355 (.A(n_8373),
    .B(n_8374),
    .Y(n_8375));
 MAJIxp5_ASAP7_75t_SL g17356 (.A(n_6905),
    .B(n_6904),
    .C(n_6903),
    .Y(n_8373));
 MAJIxp5_ASAP7_75t_SL g17357 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_39),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_21),
    .Y(n_8374));
 NAND2xp33_ASAP7_75t_SL g17359 (.A(n_8374),
    .B(n_8373),
    .Y(n_8377));
 NOR2xp33_ASAP7_75t_SL g17360 (.A(n_8373),
    .B(n_8374),
    .Y(n_8378));
 MAJx2_ASAP7_75t_SL g17363 (.A(n_21002),
    .B(n_21007),
    .C(n_21004),
    .Y(n_8380));
 MAJx2_ASAP7_75t_SL g17367 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_239),
    .B(n_8380),
    .C(n_9292),
    .Y(n_8387));
 NOR2xp33_ASAP7_75t_SL g17368 (.A(n_8390),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_290),
    .Y(n_8391));
 NOR2xp67_ASAP7_75t_SL g17369 (.A(n_8388),
    .B(n_21637),
    .Y(n_8390));
 XNOR2xp5_ASAP7_75t_SL g17370 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_232),
    .Y(n_8388));
 NAND2xp5_ASAP7_75t_SL g17373 (.A(n_8388),
    .B(n_21637),
    .Y(n_8392));
 INVxp67_ASAP7_75t_SL g17387 (.A(n_10311),
    .Y(n_8406));
 XNOR2xp5_ASAP7_75t_SL g17392 (.A(n_12520),
    .B(n_12518),
    .Y(n_8418));
 OAI22xp5_ASAP7_75t_SL g17394 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_87),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_41),
    .B1(n_8412),
    .B2(n_8413),
    .Y(n_8414));
 INVx1_ASAP7_75t_SL g17395 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_87),
    .Y(n_8412));
 INVx1_ASAP7_75t_SL g17396 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_41),
    .Y(n_8413));
 INVx1_ASAP7_75t_SL g17397 (.A(n_8415),
    .Y(n_8416));
 NAND2xp5_ASAP7_75t_SL g17398 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_61),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_91),
    .Y(n_8415));
 AND2x2_ASAP7_75t_SL g17402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_41),
    .Y(n_8421));
 NAND2xp5_ASAP7_75t_SL g17403 (.A(n_8412),
    .B(n_8413),
    .Y(n_8422));
 AOI22xp5_ASAP7_75t_SL g17408 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_152),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_110),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_22),
    .Y(n_8428));
 XNOR2x1_ASAP7_75t_SL g17412 (.B(n_8441),
    .Y(n_8442),
    .A(n_8440));
 AOI22xp5_ASAP7_75t_SL g17413 (.A1(n_8437),
    .A2(n_8439),
    .B1(n_8436),
    .B2(n_8438),
    .Y(n_8440));
 INVx1_ASAP7_75t_SL g17414 (.A(n_8436),
    .Y(n_8437));
 XNOR2x1_ASAP7_75t_SL g17415 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_2),
    .Y(n_8436),
    .A(n_22056));
 INVx1_ASAP7_75t_SL g17416 (.A(n_8438),
    .Y(n_8439));
 XNOR2x2_ASAP7_75t_SL g17417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_101),
    .Y(n_8438));
 HB1xp67_ASAP7_75t_SL g17437 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30),
    .Y(n_8461));
 OAI21xp5_ASAP7_75t_SL g17447 (.A1(n_19868),
    .A2(n_8473),
    .B(n_19792),
    .Y(n_8474));
 AOI21xp5_ASAP7_75t_SL g17448 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .A2(n_19792),
    .B(n_8473),
    .Y(n_8476));
 XOR2xp5_ASAP7_75t_SL g17451 (.A(n_8478),
    .B(n_11036),
    .Y(n_8481));
 OR2x2_ASAP7_75t_SL g17452 (.A(n_14382),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_274),
    .Y(n_8478));
 XNOR2xp5_ASAP7_75t_SL g17459 (.A(n_8486),
    .B(n_8489),
    .Y(n_8490));
 NAND2xp5_ASAP7_75t_SL g17460 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_746),
    .Y(n_8486));
 AOI22xp5_ASAP7_75t_SL g17461 (.A1(n_24230),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_683),
    .B1(n_8488),
    .B2(n_24231),
    .Y(n_8489));
 INVx1_ASAP7_75t_SL g17463 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_683),
    .Y(n_8488));
 INVxp67_ASAP7_75t_SL g17465 (.A(n_8490),
    .Y(n_8492));
 MAJIxp5_ASAP7_75t_SL g17466 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_683),
    .B(n_24231),
    .C(n_8494),
    .Y(n_8495));
 INVx1_ASAP7_75t_SL g17467 (.A(n_8486),
    .Y(n_8494));
 MAJx2_ASAP7_75t_SL g17468 (.A(n_10686),
    .B(n_8496),
    .C(n_8500),
    .Y(n_8501));
 HB1xp67_ASAP7_75t_SL g17469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_29),
    .Y(n_8496));
 XOR2x2_ASAP7_75t_SL g17470 (.A(n_8497),
    .B(n_8499),
    .Y(n_8500));
 OAI22xp5_ASAP7_75t_SL g17471 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_172),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_186),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_173),
    .Y(n_8497));
 HB1xp67_ASAP7_75t_SL g17472 (.A(n_8498),
    .Y(n_8499));
 MAJIxp5_ASAP7_75t_SL g17473 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_157),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_4),
    .Y(n_8498));
 MAJx2_ASAP7_75t_SL g17479 (.A(n_21370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_212),
    .C(n_5627),
    .Y(n_8505));
 HB1xp67_ASAP7_75t_SL g17484 (.A(n_21250),
    .Y(n_8512));
 NAND2xp33_ASAP7_75t_SRAM g17491 (.A(n_19719),
    .B(n_11533),
    .Y(n_8519));
 NOR2xp33_ASAP7_75t_SRAM g17492 (.A(n_11533),
    .B(n_19719),
    .Y(n_8520));
 AND2x2_ASAP7_75t_SL g17496 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_740),
    .Y(n_8522));
 INVxp67_ASAP7_75t_SL g17498 (.A(n_22104),
    .Y(n_8525));
 AND2x2_ASAP7_75t_SL g17500 (.A(n_4645),
    .B(n_22290),
    .Y(n_8527));
 OR2x2_ASAP7_75t_SL g17501 (.A(n_4645),
    .B(n_22290),
    .Y(n_8528));
 MAJx2_ASAP7_75t_SL g17503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_26),
    .Y(n_8530));
 INVx1_ASAP7_75t_SL g17504 (.A(n_8531),
    .Y(n_8532));
 NOR2xp33_ASAP7_75t_SL g17505 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_90),
    .Y(n_8531));
 INVx1_ASAP7_75t_SL g17532 (.A(n_8567),
    .Y(n_8568));
 XNOR2xp5_ASAP7_75t_SL g17533 (.A(n_8563),
    .B(n_8573),
    .Y(n_8567));
 INVxp67_ASAP7_75t_SL g17538 (.A(n_8575),
    .Y(n_8576));
 NAND2x1_ASAP7_75t_SL g17539 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(n_3868),
    .Y(n_8575));
 MAJIxp5_ASAP7_75t_SL g17541 (.A(n_8580),
    .B(n_3206),
    .C(n_2805),
    .Y(n_8581));
 INVx1_ASAP7_75t_SL g17542 (.A(n_20054),
    .Y(n_8580));
 MAJIxp5_ASAP7_75t_SL g17543 (.A(n_25988),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_52),
    .C(n_8575),
    .Y(n_8582));
 XNOR2x1_ASAP7_75t_SL g17545 (.B(n_8585),
    .Y(n_8586),
    .A(n_18069));
 XNOR2x2_ASAP7_75t_SL g17547 (.A(n_6117),
    .B(n_25996),
    .Y(n_8585));
 XNOR2x1_ASAP7_75t_SL g17549 (.B(n_8587),
    .Y(n_8588),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_277));
 INVxp67_ASAP7_75t_SL g17550 (.A(n_10505),
    .Y(n_8587));
 MAJIxp5_ASAP7_75t_SL g17556 (.A(n_19029),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_22),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_111),
    .Y(n_8594));
 XNOR2x1_ASAP7_75t_SL g17559 (.B(n_8595),
    .Y(n_8596),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_210));
 INVxp67_ASAP7_75t_SL g17560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_187),
    .Y(n_8595));
 MAJIxp5_ASAP7_75t_SL g17568 (.A(n_8490),
    .B(n_21141),
    .C(n_22178),
    .Y(n_8605));
 INVx1_ASAP7_75t_SL g17570 (.A(n_3657),
    .Y(n_8606));
 INVx1_ASAP7_75t_SL g17573 (.A(n_12632),
    .Y(n_8612));
 XNOR2xp5_ASAP7_75t_SL g17575 (.A(n_8613),
    .B(n_8614),
    .Y(n_8615));
 XNOR2x1_ASAP7_75t_SL g17576 (.B(n_14702),
    .Y(n_8613),
    .A(n_8525));
 XNOR2xp5_ASAP7_75t_SL g17577 (.A(n_22716),
    .B(n_20355),
    .Y(n_8614));
 INVxp67_ASAP7_75t_SL g17590 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_719),
    .Y(n_8646));
 XNOR2xp5_ASAP7_75t_SL g17593 (.A(n_8653),
    .B(n_19625),
    .Y(n_8657));
 XOR2xp5_ASAP7_75t_SL g17594 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_170),
    .B(n_8652),
    .Y(n_8653));
 INVx1_ASAP7_75t_SL g17595 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_134),
    .Y(n_8652));
 AOI31xp33_ASAP7_75t_SL g17599 (.A1(n_8661),
    .A2(n_8662),
    .A3(n_8663),
    .B(n_8665),
    .Y(n_8666));
 MAJIxp5_ASAP7_75t_SL g176 (.A(n_12653),
    .B(n_3659),
    .C(n_21492),
    .Y(n_11246));
 INVxp67_ASAP7_75t_SRAM g1760 (.A(n_7540),
    .Y(n_5300));
 OAI21xp5_ASAP7_75t_SL g17600 (.A1(n_8658),
    .A2(n_18666),
    .B(n_8660),
    .Y(n_8661));
 NAND2xp33_ASAP7_75t_SL g17602 (.A(n_7677),
    .B(n_7676),
    .Y(n_8662));
 NAND2xp33_ASAP7_75t_SL g17603 (.A(n_7677),
    .B(n_22980),
    .Y(n_8663));
 NOR3xp33_ASAP7_75t_SL g17604 (.A(n_8658),
    .B(n_18666),
    .C(n_8660),
    .Y(n_8665));
 OAI21xp33_ASAP7_75t_SL g17607 (.A1(n_22980),
    .A2(n_7676),
    .B(n_7677),
    .Y(n_2634));
 AND2x2_ASAP7_75t_SL g17609 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_746),
    .Y(n_8670));
 NAND2xp5_ASAP7_75t_SL g17610 (.A(n_10478),
    .B(n_2162),
    .Y(n_8672));
 INVx1_ASAP7_75t_SL g17619 (.A(n_11818),
    .Y(n_8688));
 NAND2xp5_ASAP7_75t_SL g17623 (.A(n_12051),
    .B(n_14709),
    .Y(n_8690));
 AND2x2_ASAP7_75t_SL g17627 (.A(n_12050),
    .B(n_18704),
    .Y(n_8694));
 INVxp33_ASAP7_75t_R g17628 (.A(n_8696),
    .Y(n_8697));
 NOR2x1_ASAP7_75t_SL g17629 (.A(n_14709),
    .B(n_12051),
    .Y(n_8696));
 AND2x2_ASAP7_75t_SL g17635 (.A(n_20825),
    .B(n_26057),
    .Y(n_8702));
 NAND2xp5_ASAP7_75t_SL g17651 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .Y(n_8719));
 NAND2xp5_ASAP7_75t_SL g17652 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_11770),
    .Y(n_8722));
 NAND2xp5_ASAP7_75t_SL g17655 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_11770),
    .Y(n_8725));
 XNOR2x2_ASAP7_75t_SL g17664 (.A(n_8731),
    .B(n_6280),
    .Y(n_8732));
 INVxp67_ASAP7_75t_SL g17665 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_56),
    .Y(n_8731));
 NAND2x1_ASAP7_75t_SL g17666 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(n_22743),
    .Y(n_8738));
 OA21x2_ASAP7_75t_SL g17669 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_115),
    .Y(n_8739));
 MAJIxp5_ASAP7_75t_SL g17677 (.A(n_8748),
    .B(n_8752),
    .C(n_8759),
    .Y(n_8760));
 OAI21xp5_ASAP7_75t_SL g17678 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_174),
    .Y(n_8748));
 MAJIxp5_ASAP7_75t_SL g17679 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_37),
    .Y(n_8752));
 XNOR2x1_ASAP7_75t_SL g17682 (.B(n_8758),
    .Y(n_8759),
    .A(n_18916));
 INVx2_ASAP7_75t_SL g17686 (.A(n_8757),
    .Y(n_8758));
 XOR2xp5_ASAP7_75t_SL g17687 (.A(n_8756),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_124),
    .Y(n_8757));
 INVxp67_ASAP7_75t_SL g17688 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_85),
    .Y(n_8756));
 XOR2x2_ASAP7_75t_SL g17689 (.A(n_12251),
    .B(n_8768),
    .Y(n_8770));
 XOR2xp5_ASAP7_75t_SL g1769 (.A(n_5276),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_247),
    .Y(n_5277));
 MAJIxp5_ASAP7_75t_SL g17696 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_737),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_68),
    .Y(n_8768));
 INVxp67_ASAP7_75t_SL g17704 (.A(n_8776),
    .Y(n_8777));
 MAJIxp5_ASAP7_75t_SL g17705 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_74),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_72),
    .Y(n_8776));
 NAND2xp5_ASAP7_75t_SL g17727 (.A(n_10033),
    .B(n_7579),
    .Y(n_8821));
 NOR2xp67_ASAP7_75t_SL g17729 (.A(n_10033),
    .B(n_7579),
    .Y(n_8823));
 AND2x2_ASAP7_75t_SL g17731 (.A(n_26250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_275),
    .Y(n_8826));
 XNOR2xp5_ASAP7_75t_SL g17738 (.A(n_9271),
    .B(n_8839),
    .Y(n_8840));
 XOR2xp5_ASAP7_75t_SL g17740 (.A(n_8837),
    .B(n_8838),
    .Y(n_8839));
 INVx1_ASAP7_75t_SL g17741 (.A(n_8836),
    .Y(n_8837));
 MAJIxp5_ASAP7_75t_SL g17742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_84),
    .Y(n_8836));
 XNOR2x2_ASAP7_75t_SL g17743 (.A(n_7080),
    .B(n_18874),
    .Y(n_8838));
 MAJIxp5_ASAP7_75t_SL g17746 (.A(n_19915),
    .B(n_8732),
    .C(n_19363),
    .Y(n_8841));
 XNOR2x1_ASAP7_75t_SL g17750 (.B(n_8851),
    .Y(n_8852),
    .A(n_8849));
 XNOR2xp5_ASAP7_75t_SL g17751 (.A(n_8847),
    .B(n_8848),
    .Y(n_8849));
 NAND2x1_ASAP7_75t_SL g17752 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_582),
    .Y(n_8847));
 NAND2xp5_ASAP7_75t_SL g17753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_678),
    .B(n_2162),
    .Y(n_8848));
 INVx1_ASAP7_75t_SL g17754 (.A(n_8850),
    .Y(n_8851));
 AND2x2_ASAP7_75t_SL g17755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_742),
    .B(n_2174),
    .Y(n_8850));
 INVxp67_ASAP7_75t_SL g17756 (.A(n_8848),
    .Y(n_8853));
 NOR2xp67_ASAP7_75t_SL g17758 (.A(n_8855),
    .B(n_20222),
    .Y(n_8861));
 MAJIxp5_ASAP7_75t_SL g17759 (.A(n_18885),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_71),
    .C(n_7356),
    .Y(n_8855));
 XNOR2xp5_ASAP7_75t_L g17768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_15),
    .Y(n_8864));
 INVxp67_ASAP7_75t_SL g17769 (.A(n_8865),
    .Y(n_8866));
 INVxp67_ASAP7_75t_SL g1777 (.A(n_23195),
    .Y(n_5276));
 MAJIxp5_ASAP7_75t_SL g17770 (.A(n_13776),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_101),
    .C(n_22620),
    .Y(n_8865));
 OAI22xp5_ASAP7_75t_SL g17774 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_81),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_19),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_82),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_132),
    .Y(n_8871));
 XNOR2xp5_ASAP7_75t_SL g17776 (.A(n_8873),
    .B(n_18919),
    .Y(n_8878));
 NAND2xp5_ASAP7_75t_SL g17777 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .B(n_2544),
    .Y(n_8872));
 HB1xp67_ASAP7_75t_SL g17782 (.A(n_14111),
    .Y(n_8882));
 INVx2_ASAP7_75t_SL g17786 (.A(n_8886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41));
 XNOR2x1_ASAP7_75t_SL g17787 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_737),
    .Y(n_8886),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_4));
 OR2x2_ASAP7_75t_SL g17789 (.A(n_17416),
    .B(n_26202),
    .Y(n_8888));
 NAND2xp5_ASAP7_75t_SL g17798 (.A(n_19958),
    .B(n_8901),
    .Y(n_8902));
 NAND2xp5_ASAP7_75t_SL g17799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_269),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_273),
    .Y(n_8901));
 AOI211xp5_ASAP7_75t_SL g178 (.A1(n_22141),
    .A2(n_22142),
    .B(n_18767),
    .C(n_22143),
    .Y(n_22147));
 XNOR2xp5_ASAP7_75t_SL g17812 (.A(n_19149),
    .B(n_8927),
    .Y(n_8928));
 OAI22xp5_ASAP7_75t_SL g17814 (.A1(n_8924),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .B1(n_8925),
    .B2(n_8926),
    .Y(n_8927));
 OAI22xp5_ASAP7_75t_SL g17815 (.A1(n_8919),
    .A2(n_8923),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_n_757),
    .B2(n_19150),
    .Y(n_8924));
 INVx1_ASAP7_75t_SL g17816 (.A(n_19150),
    .Y(n_8923));
 INVxp67_ASAP7_75t_SL g17818 (.A(n_8924),
    .Y(n_8925));
 XNOR2x1_ASAP7_75t_SL g17830 (.B(n_8947),
    .Y(n_8948),
    .A(n_21944));
 NAND2xp5_ASAP7_75t_SL g17832 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .Y(n_8943));
 INVxp67_ASAP7_75t_SL g17834 (.A(n_8943),
    .Y(n_8945));
 HB1xp67_ASAP7_75t_SL g17835 (.A(n_4856),
    .Y(n_8947));
 OAI21x1_ASAP7_75t_SL g17838 (.A1(n_11760),
    .A2(n_11058),
    .B(n_11056),
    .Y(n_8951));
 MAJx2_ASAP7_75t_SL g17841 (.A(n_8955),
    .B(n_8957),
    .C(n_11456),
    .Y(n_8959));
 INVx1_ASAP7_75t_SL g17842 (.A(n_8954),
    .Y(n_8955));
 XNOR2xp5_ASAP7_75t_SL g17843 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_18),
    .Y(n_8954));
 INVxp67_ASAP7_75t_SL g17844 (.A(n_8956),
    .Y(n_8957));
 MAJIxp5_ASAP7_75t_SL g17845 (.A(n_18793),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_655),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_623),
    .Y(n_8956));
 INVxp67_ASAP7_75t_SL g17849 (.A(n_21250),
    .Y(n_8962));
 NOR2x1_ASAP7_75t_SL g17861 (.A(n_8973),
    .B(n_8974),
    .Y(n_8975));
 NOR2x1_ASAP7_75t_SL g17862 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_72),
    .Y(n_8973));
 NOR2x1_ASAP7_75t_SL g17863 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_113),
    .Y(n_8974));
 OAI21xp5_ASAP7_75t_SL g17865 (.A1(n_8985),
    .A2(n_8989),
    .B(n_8990),
    .Y(n_8991));
 NOR2xp33_ASAP7_75t_SL g17866 (.A(n_8981),
    .B(n_8984),
    .Y(n_8985));
 INVxp67_ASAP7_75t_SL g17867 (.A(n_8980),
    .Y(n_8981));
 MAJIxp5_ASAP7_75t_SL g17868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_45),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_29),
    .Y(n_8980));
 AOI22xp5_ASAP7_75t_SL g17871 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_158),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_162),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_157),
    .B2(n_8983),
    .Y(n_8984));
 INVx1_ASAP7_75t_SL g17873 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_162),
    .Y(n_8983));
 AO21x1_ASAP7_75t_L g17874 (.A1(n_18695),
    .A2(n_18749),
    .B(n_8988),
    .Y(n_8989));
 INVx1_ASAP7_75t_SL g17876 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_180),
    .Y(n_8988));
 NAND2xp5_ASAP7_75t_SL g17877 (.A(n_8981),
    .B(n_8984),
    .Y(n_8990));
 INVx1_ASAP7_75t_SL g17878 (.A(n_8984),
    .Y(n_8993));
 NAND2xp5_ASAP7_75t_SL g17889 (.A(n_10416),
    .B(n_26208),
    .Y(n_9008));
 XOR2x1_ASAP7_75t_SL g17895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_743),
    .Y(n_9009),
    .B(n_18839));
 HB1xp67_ASAP7_75t_SL g179 (.A(n_8474),
    .Y(n_6079));
 XNOR2xp5_ASAP7_75t_SL g17907 (.A(n_9031),
    .B(n_9032),
    .Y(n_9033));
 NAND2xp5_ASAP7_75t_SL g17908 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .Y(n_9031));
 NAND2xp5_ASAP7_75t_SL g17909 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .Y(n_9032));
 INVxp67_ASAP7_75t_SL g17910 (.A(n_9031),
    .Y(n_9034));
 NOR2xp67_ASAP7_75t_SL g17911 (.A(n_9035),
    .B(n_9036),
    .Y(n_9037));
 NAND2xp5_ASAP7_75t_SL g17912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_290),
    .B(n_22488),
    .Y(n_9035));
 NAND2xp5_ASAP7_75t_SL g17913 (.A(n_10161),
    .B(n_6194),
    .Y(n_9036));
 MAJIxp5_ASAP7_75t_SL g17914 (.A(n_9739),
    .B(n_9740),
    .C(n_9041),
    .Y(n_9042));
 INVx1_ASAP7_75t_SL g17916 (.A(n_15585),
    .Y(n_9038));
 MAJx2_ASAP7_75t_SL g17918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_5),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_127),
    .C(n_24405),
    .Y(n_9041));
 HB1xp67_ASAP7_75t_SL g17926 (.A(n_22618),
    .Y(n_9048));
 NOR2xp67_ASAP7_75t_L g17930 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_647),
    .B(n_22097),
    .Y(n_9053));
 NAND2xp5_ASAP7_75t_SL g17931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_647),
    .B(n_22097),
    .Y(n_9054));
 NAND2xp5_ASAP7_75t_SL g17934 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .Y(n_9059));
 INVxp67_ASAP7_75t_SL g17937 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_95),
    .Y(n_9061));
 NAND2xp5_ASAP7_75t_SL g17941 (.A(n_2154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_746),
    .Y(n_9065));
 MAJx2_ASAP7_75t_SL g17943 (.A(n_9069),
    .B(n_9070),
    .C(n_5826),
    .Y(n_9074));
 NAND2x1_ASAP7_75t_SL g17944 (.A(n_2181),
    .B(n_11341),
    .Y(n_9069));
 NAND2xp5_ASAP7_75t_SL g17945 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_716),
    .Y(n_9070));
 NAND2xp5_ASAP7_75t_SL g17947 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_780),
    .B(n_21789),
    .Y(n_5826));
 INVx1_ASAP7_75t_SL g17948 (.A(n_9070),
    .Y(n_9076));
 XNOR2xp5_ASAP7_75t_SL g17949 (.A(n_9077),
    .B(n_9078),
    .Y(n_9079));
 NAND2xp5_ASAP7_75t_SL g17950 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .Y(n_9077));
 NAND2xp5_ASAP7_75t_SL g17951 (.A(n_3479),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .Y(n_9078));
 INVx1_ASAP7_75t_SL g17952 (.A(n_9078),
    .Y(n_9080));
 XNOR2x1_ASAP7_75t_SL g17961 (.B(n_11829),
    .Y(n_9094),
    .A(n_9091));
 MAJx2_ASAP7_75t_SL g17962 (.A(n_13724),
    .B(n_4026),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_111),
    .Y(n_9091));
 INVx1_ASAP7_75t_SL g17964 (.A(n_6094),
    .Y(n_9092));
 XNOR2xp5_ASAP7_75t_SL g17972 (.A(n_9104),
    .B(n_9105),
    .Y(n_9106));
 INVx1_ASAP7_75t_SL g17973 (.A(n_7010),
    .Y(n_9104));
 XNOR2xp5_ASAP7_75t_SL g17974 (.A(n_7000),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_8),
    .Y(n_7010));
 MAJIxp5_ASAP7_75t_SL g17976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_148),
    .B(n_6997),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_128),
    .Y(n_9105));
 XNOR2x1_ASAP7_75t_SL g17977 (.B(n_26071),
    .Y(n_9111),
    .A(n_9107));
 XNOR2xp5_ASAP7_75t_SL g17978 (.A(n_9009),
    .B(n_14301),
    .Y(n_9107));
 MAJIxp5_ASAP7_75t_SL g17982_dup (.A(n_12252),
    .B(n_26175),
    .C(n_12254),
    .Y(n_12257));
 MAJIxp5_ASAP7_75t_SL g17991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_109),
    .C(n_13721),
    .Y(n_9120));
 INVx1_ASAP7_75t_SL g17992 (.A(n_9120),
    .Y(n_9123));
 OAI21xp5_ASAP7_75t_SL g17994 (.A1(n_7620),
    .A2(n_9124),
    .B(n_9125),
    .Y(n_9126));
 AND2x2_ASAP7_75t_SL g17995 (.A(n_19910),
    .B(n_20124),
    .Y(n_9124));
 OR2x2_ASAP7_75t_SL g17996 (.A(n_20124),
    .B(n_19910),
    .Y(n_9125));
 MAJIxp5_ASAP7_75t_SL g180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_188),
    .B(n_19660),
    .C(n_5133),
    .Y(n_19661));
 AOI22xp5_ASAP7_75t_SL g18004 (.A1(n_9136),
    .A2(n_9138),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_151),
    .B2(n_9140),
    .Y(n_9141));
 INVxp67_ASAP7_75t_SL g18005 (.A(n_8461),
    .Y(n_9136));
 INVx1_ASAP7_75t_SL g18008 (.A(n_11350),
    .Y(n_9140));
 OAI22xp33_ASAP7_75t_SL g18009 (.A1(n_11346),
    .A2(n_8461),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_152),
    .B2(n_11350),
    .Y(n_9143));
 BUFx12f_ASAP7_75t_SL g18019 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[46]),
    .Y(n_9154));
 NAND2xp33_ASAP7_75t_SL g18021 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .Y(n_9155));
 AND2x2_ASAP7_75t_SRAM g18022 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[47]),
    .Y(n_9156));
 XNOR2xp5_ASAP7_75t_SL g18023 (.A(n_3088),
    .B(n_10360),
    .Y(n_9162));
 MAJIxp5_ASAP7_75t_SL g18024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_16),
    .C(n_19436),
    .Y(n_3088));
 INVx1_ASAP7_75t_SL g18027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_80),
    .Y(n_9160));
 NAND2x1_ASAP7_75t_SL g18038 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_14987),
    .Y(n_9172));
 MAJx2_ASAP7_75t_SL g18044 (.A(n_9179),
    .B(n_9180),
    .C(n_9181),
    .Y(n_9182));
 AOI22xp5_ASAP7_75t_SL g18045 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_98),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_58),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_97),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_59),
    .Y(n_9179));
 NAND2xp5_ASAP7_75t_SL g18046 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B(n_3709),
    .Y(n_9180));
 NAND2xp5_ASAP7_75t_SL g18047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_52),
    .Y(n_9181));
 INVx1_ASAP7_75t_SL g18048 (.A(n_9181),
    .Y(n_9183));
 INVx1_ASAP7_75t_SL g18066 (.A(n_9214),
    .Y(n_9215));
 XNOR2xp5_ASAP7_75t_SL g18067 (.A(n_8852),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_21),
    .Y(n_9214));
 AOI22xp5_ASAP7_75t_SL g18070 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_155),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_140),
    .B1(n_26173),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_156),
    .Y(n_9218));
 XNOR2xp5_ASAP7_75t_SL g18079 (.A(n_12565),
    .B(n_26258),
    .Y(n_9234));
 XOR2xp5_ASAP7_75t_SL g18083 (.A(n_21646),
    .B(n_9237),
    .Y(n_9238));
 MAJIxp5_ASAP7_75t_SL g18084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .C(n_6119),
    .Y(n_9237));
 XNOR2x2_ASAP7_75t_SL g18090 (.A(n_9244),
    .B(n_18851),
    .Y(n_9246));
 AND2x2_ASAP7_75t_SL g18091 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_736),
    .Y(n_9244));
 AOI21xp5_ASAP7_75t_SL g18096 (.A1(n_9252),
    .A2(n_9253),
    .B(n_9254),
    .Y(n_9255));
 OAI21xp5_ASAP7_75t_SL g18097 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_199),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_201),
    .Y(n_9252));
 NAND2xp5_ASAP7_75t_SL g18098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_181),
    .B(n_6769),
    .Y(n_9253));
 NOR2x1_ASAP7_75t_SL g18099 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_181),
    .B(n_6769),
    .Y(n_9254));
 OAI21xp5_ASAP7_75t_SL g181 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_207),
    .A2(n_10731),
    .B(n_10732),
    .Y(n_19662));
 XNOR2xp5_ASAP7_75t_SL g18101 (.A(n_18865),
    .B(n_9258),
    .Y(n_9259));
 AOI22xp5_ASAP7_75t_SL g18103 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_126),
    .A2(n_6710),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_146),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_127),
    .Y(n_9258));
 AOI22xp33_ASAP7_75t_SL g18106 (.A1(n_12111),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_110),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_152),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109),
    .Y(n_9261));
 OR2x2_ASAP7_75t_SL g18109 (.A(n_22218),
    .B(n_22216),
    .Y(n_9263));
 XNOR2x1_ASAP7_75t_SL g18111 (.B(n_9270),
    .Y(n_9271),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_131));
 OAI22xp5_ASAP7_75t_SL g18112 (.A1(n_9267),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_76),
    .B1(n_9269),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_77),
    .Y(n_9270));
 NAND2xp5_ASAP7_75t_SL g18113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_105),
    .B(n_13699),
    .Y(n_9267));
 BUFx12f_ASAP7_75t_SL g18116 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[39]),
    .Y(n_9273));
 NAND2xp5_ASAP7_75t_SL g18118 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[39]),
    .Y(n_9274));
 XNOR2xp5_ASAP7_75t_SL g18120 (.A(n_23113),
    .B(n_14877),
    .Y(n_9281));
 INVx1_ASAP7_75t_SL g18124 (.A(n_26137),
    .Y(n_9279));
 XNOR2xp5_ASAP7_75t_SL g18133 (.A(n_9293),
    .B(n_20900),
    .Y(n_9295));
 INVx1_ASAP7_75t_SL g18134 (.A(n_9292),
    .Y(n_9293));
 MAJIxp5_ASAP7_75t_SL g18135 (.A(n_20842),
    .B(n_19390),
    .C(n_21988),
    .Y(n_9292));
 XOR2xp5_ASAP7_75t_SL g18138 (.A(n_9297),
    .B(n_9298),
    .Y(n_9299));
 XOR2xp5_ASAP7_75t_SL g18139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_8),
    .B(n_9296),
    .Y(n_9297));
 INVx1_ASAP7_75t_SL g18140 (.A(n_10915),
    .Y(n_9296));
 MAJIxp5_ASAP7_75t_SL g18141 (.A(n_5553),
    .B(n_15210),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_126),
    .Y(n_9298));
 AND2x4_ASAP7_75t_SL g18146 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_pvld[7]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_pvld[7]),
    .Y(n_9301));
 NOR2xp33_ASAP7_75t_SL g18149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[11]),
    .B(n_9301),
    .Y(n_9305));
 XNOR2xp5_ASAP7_75t_SL g18154 (.A(n_26008),
    .B(n_18926),
    .Y(n_9316));
 NAND2x1p5_ASAP7_75t_SL g18158 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B(n_19391),
    .Y(n_9313));
 XOR2xp5_ASAP7_75t_SL g18159 (.A(n_9317),
    .B(n_19360),
    .Y(n_9321));
 XOR2xp5_ASAP7_75t_SL g18160 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_8),
    .Y(n_9317));
 XNOR2xp5_ASAP7_75t_SL g18165 (.A(n_9324),
    .B(n_9325),
    .Y(n_9326));
 XNOR2x2_ASAP7_75t_SL g18166 (.A(n_9323),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_6),
    .Y(n_9324));
 INVxp67_ASAP7_75t_SL g18167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_65),
    .Y(n_9323));
 XNOR2xp5_ASAP7_75t_SL g18168 (.A(n_9274),
    .B(n_13327),
    .Y(n_9325));
 NAND2xp5_ASAP7_75t_SL g18172 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(n_9327));
 AOI21x1_ASAP7_75t_SL g18174 (.A1(n_9333),
    .A2(n_9335),
    .B(n_9337),
    .Y(n_9338));
 INVx1_ASAP7_75t_SL g18175 (.A(n_21508),
    .Y(n_9333));
 HB1xp67_ASAP7_75t_SL g18177 (.A(n_9334),
    .Y(n_9335));
 NOR2xp67_ASAP7_75t_SL g18178 (.A(n_7072),
    .B(n_11965),
    .Y(n_9334));
 HB1xp67_ASAP7_75t_SL g18179 (.A(n_9336),
    .Y(n_9337));
 OAI21x1_ASAP7_75t_SL g18180 (.A1(n_11967),
    .A2(n_7072),
    .B(n_7073),
    .Y(n_9336));
 MAJIxp5_ASAP7_75t_SL g18183 (.A(n_9339),
    .B(n_9340),
    .C(n_9341),
    .Y(n_9342));
 INVxp67_ASAP7_75t_SL g18184 (.A(n_22621),
    .Y(n_9339));
 INVx1_ASAP7_75t_SL g18185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_101),
    .Y(n_9340));
 INVx2_ASAP7_75t_SL g18186 (.A(n_13788),
    .Y(n_9341));
 XNOR2xp5_ASAP7_75t_SL g18188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_20),
    .Y(n_9344));
 NAND2xp5_ASAP7_75t_SL g18196 (.A(n_2180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_642),
    .Y(n_9354));
 OAI321xp33_ASAP7_75t_SL g182 (.A1(n_21392),
    .A2(n_13009),
    .A3(n_13012),
    .B1(n_13014),
    .B2(n_21392),
    .C(n_21393),
    .Y(n_13521));
 INVx1_ASAP7_75t_SL g18203 (.A(n_4902),
    .Y(n_9359));
 AOI21xp5_ASAP7_75t_SL g18205 (.A1(n_2852),
    .A2(n_21479),
    .B(n_21480),
    .Y(n_9367));
 NOR2xp67_ASAP7_75t_SL g18207 (.A(n_10841),
    .B(n_19445),
    .Y(n_2852));
 XNOR2x1_ASAP7_75t_SL g18209 (.B(n_9368),
    .Y(n_9370),
    .A(n_11932));
 NAND2x1p5_ASAP7_75t_SL g18210 (.A(n_2161),
    .B(n_12642),
    .Y(n_9368));
 INVx1_ASAP7_75t_SL g18215 (.A(n_13241),
    .Y(n_9373));
 INVxp67_ASAP7_75t_SL g18217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106),
    .Y(n_9376));
 OAI22xp5_ASAP7_75t_SL g18218 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106),
    .A2(n_9373),
    .B1(n_9376),
    .B2(n_13241),
    .Y(n_9379));
 NAND2xp5_ASAP7_75t_SL g18226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_282),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_8),
    .Y(n_9385));
 INVx1_ASAP7_75t_SL g18227 (.A(n_21364),
    .Y(n_9388));
 MAJx2_ASAP7_75t_SL g18229 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_39),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_21),
    .Y(n_9389));
 NOR2x1_ASAP7_75t_SL g18232 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_282),
    .B(n_25983),
    .Y(n_9392));
 XNOR2xp5_ASAP7_75t_SL g18240 (.A(n_9402),
    .B(n_22736),
    .Y(n_9404));
 HB1xp67_ASAP7_75t_SL g18241 (.A(n_12218),
    .Y(n_9402));
 AND2x2_ASAP7_75t_SL g18245 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_653),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_621),
    .Y(n_9405));
 OR2x2_ASAP7_75t_SL g18246 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_653),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_621),
    .Y(n_9406));
 OAI21xp5_ASAP7_75t_SL g18247 (.A1(n_9405),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_133),
    .B(n_9406),
    .Y(n_9410));
 INVx1_ASAP7_75t_SL g18256 (.A(n_9419),
    .Y(n_9420));
 XNOR2xp5_ASAP7_75t_SL g18262 (.A(n_21311),
    .B(n_10623),
    .Y(n_9430));
 NAND2xp5_ASAP7_75t_SL g18268 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .Y(n_9432));
 NAND2x1_ASAP7_75t_SL g18269 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(n_14523),
    .Y(n_9434));
 NAND2xp5_ASAP7_75t_SL g18276 (.A(n_2985),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .Y(n_9441));
 INVx1_ASAP7_75t_SL g18279 (.A(n_11249),
    .Y(n_9447));
 XOR2xp5_ASAP7_75t_SL g18281 (.A(n_9449),
    .B(n_9450),
    .Y(n_9451));
 MAJIxp5_ASAP7_75t_SL g18282 (.A(n_7462),
    .B(n_13577),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_186),
    .Y(n_9449));
 XOR2x2_ASAP7_75t_SL g18283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_188),
    .B(n_13576),
    .Y(n_9450));
 INVx1_ASAP7_75t_SL g18285 (.A(n_9449),
    .Y(n_9453));
 NOR2xp67_ASAP7_75t_SL g18286 (.A(n_12892),
    .B(n_9455),
    .Y(n_9456));
 NAND2xp5_ASAP7_75t_SL g18288 (.A(n_7697),
    .B(n_7698),
    .Y(n_9455));
 OAI22xp5_ASAP7_75t_SL g18289 (.A1(n_18927),
    .A2(n_9464),
    .B1(n_5513),
    .B2(n_5514),
    .Y(n_9467));
 OAI21x1_ASAP7_75t_SL g18293 (.A1(n_9462),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_71),
    .B(n_9463),
    .Y(n_9464));
 AND2x2_ASAP7_75t_SL g18294 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_70),
    .Y(n_9462));
 OR2x2_ASAP7_75t_SL g18295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_54),
    .Y(n_9463));
 XNOR2x1_ASAP7_75t_SL g18298 (.B(n_9470),
    .Y(n_9471),
    .A(n_18754));
 XOR2xp5_ASAP7_75t_SL g183 (.A(n_21423),
    .B(n_18938),
    .Y(n_21424));
 AND2x2_ASAP7_75t_SL g18300 (.A(n_3468),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .Y(n_9470));
 XNOR2xp5_ASAP7_75t_SL g18303 (.A(n_18928),
    .B(n_9479),
    .Y(n_9480));
 INVx1_ASAP7_75t_SL g18307 (.A(n_20233),
    .Y(n_9479));
 NOR2xp67_ASAP7_75t_SL g18311 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_14),
    .Y(n_9481));
 NAND2xp5_ASAP7_75t_SL g18313 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_14),
    .Y(n_9483));
 NOR2xp67_ASAP7_75t_SL g18324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_362),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_400),
    .Y(n_9494));
 NAND2xp5_ASAP7_75t_SL g18327 (.A(n_5793),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_243),
    .Y(n_9498));
 NAND2xp5_ASAP7_75t_SL g18328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_240),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_255),
    .Y(n_9503));
 XNOR2xp5_ASAP7_75t_SL g18330 (.A(n_14443),
    .B(n_13359),
    .Y(n_9510));
 NOR2xp33_ASAP7_75t_SL g18333 (.A(n_22037),
    .B(n_10419),
    .Y(n_9513));
 NOR2x1_ASAP7_75t_SL g18338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_46),
    .B(n_12120),
    .Y(n_9514));
 AOI22xp5_ASAP7_75t_SL g18339 (.A1(n_13710),
    .A2(n_15156),
    .B1(n_15157),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_95),
    .Y(n_9516));
 OR2x2_ASAP7_75t_SL g18340 (.A(n_12639),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_276),
    .Y(n_9518));
 MAJIxp5_ASAP7_75t_SL g18348 (.A(n_6339),
    .B(n_6342),
    .C(n_6343),
    .Y(n_9525));
 NAND2x1_ASAP7_75t_SL g18354 (.A(n_2825),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .Y(n_9534));
 MAJIxp5_ASAP7_75t_SL g18358 (.A(n_6431),
    .B(n_6430),
    .C(n_2277),
    .Y(n_9536));
 XNOR2x1_ASAP7_75t_SL g18362 (.B(n_6754),
    .Y(n_9541),
    .A(n_19208));
 INVx1_ASAP7_75t_SL g18365 (.A(n_10713),
    .Y(n_9544));
 XOR2xp5_ASAP7_75t_SL g18366 (.A(n_9548),
    .B(n_8256),
    .Y(n_9549));
 AOI22xp5_ASAP7_75t_SL g18367 (.A1(n_9546),
    .A2(n_8255),
    .B1(n_9545),
    .B2(n_8259),
    .Y(n_9548));
 INVx1_ASAP7_75t_SL g18368 (.A(n_9545),
    .Y(n_9546));
 NAND2x1_ASAP7_75t_SL g18369 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(n_3275),
    .Y(n_9545));
 AND2x2_ASAP7_75t_SL g18387 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .Y(n_9570));
 MAJIxp5_ASAP7_75t_SL g18388 (.A(n_9574),
    .B(n_9575),
    .C(n_9576),
    .Y(n_9577));
 INVx1_ASAP7_75t_SL g18389 (.A(n_9573),
    .Y(n_9574));
 NAND2x1_ASAP7_75t_SL g18390 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(n_19645),
    .Y(n_9573));
 AND2x2_ASAP7_75t_SL g18391 (.A(n_14975),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .Y(n_9575));
 NAND2x1_ASAP7_75t_SL g18392 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(n_9576));
 AOI21x1_ASAP7_75t_SL g184 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_309),
    .A2(n_14800),
    .B(n_6546),
    .Y(n_14802));
 XNOR2x1_ASAP7_75t_SL g18400 (.B(n_20729),
    .Y(n_9591),
    .A(n_18757));
 XOR2xp5_ASAP7_75t_SL g18416 (.A(n_9603),
    .B(n_9604),
    .Y(n_9605));
 XNOR2x2_ASAP7_75t_SL g18417 (.A(n_26242),
    .B(n_18811),
    .Y(n_9603));
 MAJx2_ASAP7_75t_SL g18419 (.A(n_8948),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_172),
    .Y(n_9604));
 NOR2xp67_ASAP7_75t_SL g18428 (.A(n_9614),
    .B(n_19909),
    .Y(n_9616));
 OAI22xp5_ASAP7_75t_SL g18431 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_329),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_54),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_311),
    .B2(n_4102),
    .Y(n_9617));
 XNOR2xp5_ASAP7_75t_SL g18432 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_23),
    .Y(n_9618));
 NOR2xp33_ASAP7_75t_SL g18437 (.A(n_9625),
    .B(n_10090),
    .Y(n_9627));
 MAJIxp5_ASAP7_75t_SL g18438 (.A(n_13201),
    .B(n_9624),
    .C(n_2283),
    .Y(n_9625));
 AND2x2_ASAP7_75t_SL g18442 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(n_3309),
    .Y(n_9628));
 MAJIxp5_ASAP7_75t_SL g18444 (.A(n_9631),
    .B(n_9632),
    .C(n_9633),
    .Y(n_9634));
 MAJx2_ASAP7_75t_SL g18445 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_116),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_142),
    .Y(n_9631));
 XNOR2x1_ASAP7_75t_SL g18446 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_0),
    .Y(n_9633),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_4));
 XNOR2xp5_ASAP7_75t_SL g18447 (.A(n_9635),
    .B(n_9636),
    .Y(n_9637));
 NAND2x1_ASAP7_75t_SL g18448 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_22019),
    .Y(n_9635));
 NOR2x1_ASAP7_75t_SL g18449 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_43),
    .B(n_4550),
    .Y(n_9636));
 INVx1_ASAP7_75t_SL g18450 (.A(n_9635),
    .Y(n_9638));
 INVx1_ASAP7_75t_SL g18451 (.A(n_9636),
    .Y(n_9639));
 XOR2xp5_ASAP7_75t_SL g18452 (.A(n_19270),
    .B(n_22465),
    .Y(n_9642));
 AND2x2_ASAP7_75t_SL g18465 (.A(n_2159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_588),
    .Y(n_9650));
 INVx1_ASAP7_75t_SL g18466 (.A(n_9652),
    .Y(n_9653));
 AND2x2_ASAP7_75t_SL g18467 (.A(n_2162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_684),
    .Y(n_9652));
 AND2x2_ASAP7_75t_SL g18470 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_554),
    .B(n_2182),
    .Y(n_9657));
 AND2x2_ASAP7_75t_SL g18471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_778),
    .B(n_24102),
    .Y(n_9658));
 AND2x2_ASAP7_75t_SL g18472 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_714),
    .B(n_19370),
    .Y(n_9659));
 BUFx3_ASAP7_75t_L g18473 (.A(n_2177),
    .Y(n_9661));
 BUFx3_ASAP7_75t_L g18474 (.A(n_2155),
    .Y(n_9662));
 MAJIxp5_ASAP7_75t_SL g18480 (.A(n_22104),
    .B(n_9669),
    .C(n_14701),
    .Y(n_9671));
 MAJx2_ASAP7_75t_SL g18482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_583),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_743),
    .C(n_5783),
    .Y(n_9669));
 XOR2xp5_ASAP7_75t_SL g18484 (.A(n_9672),
    .B(n_21572),
    .Y(n_9677));
 INVxp67_ASAP7_75t_SL g18485 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_100),
    .Y(n_9672));
 INVx1_ASAP7_75t_SL g18488 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_54),
    .Y(n_9675));
 XNOR2x1_ASAP7_75t_SL g18489 (.B(n_18934),
    .Y(n_9682),
    .A(n_20054));
 XNOR2xp5_ASAP7_75t_SL g18494 (.A(n_24680),
    .B(n_9685),
    .Y(n_9686));
 XNOR2xp5_ASAP7_75t_SL g18496 (.A(n_9684),
    .B(n_26060),
    .Y(n_9685));
 INVx1_ASAP7_75t_SL g18497 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_80),
    .Y(n_9684));
 INVx1_ASAP7_75t_SL g185 (.A(n_23386),
    .Y(n_6186));
 XOR2xp5_ASAP7_75t_SL g18503 (.A(n_9693),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_87),
    .Y(n_9694));
 XNOR2xp5_ASAP7_75t_SL g18504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_104),
    .B(n_9692),
    .Y(n_9693));
 NAND2x1_ASAP7_75t_SL g18505 (.A(n_22865),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .Y(n_9692));
 NOR2xp67_ASAP7_75t_SL g18507 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_284),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_290),
    .Y(n_9695));
 INVxp67_ASAP7_75t_SL g18509 (.A(n_9697),
    .Y(n_9698));
 OAI21xp5_ASAP7_75t_SL g18510 (.A1(n_8390),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_291),
    .B(n_8392),
    .Y(n_9697));
 XOR2x2_ASAP7_75t_SL g18512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_44),
    .Y(n_9700));
 XNOR2xp5_ASAP7_75t_SL g18519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_9),
    .B(n_6439),
    .Y(n_9708));
 MAJx2_ASAP7_75t_SL g18520 (.A(n_6377),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_172),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_186),
    .Y(n_9709));
 INVx1_ASAP7_75t_SL g18521 (.A(n_9708),
    .Y(n_9711));
 XOR2xp5_ASAP7_75t_SL g18524 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_29),
    .B(n_13148),
    .Y(n_9713));
 XOR2xp5_ASAP7_75t_SL g18535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_559),
    .B(n_9725),
    .Y(n_9726));
 NAND2xp5_ASAP7_75t_SL g18536 (.A(n_20825),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_718),
    .Y(n_9725));
 INVxp67_ASAP7_75t_SL g18537 (.A(n_9725),
    .Y(n_9728));
 XNOR2xp5_ASAP7_75t_SL g18549 (.A(n_9038),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_135),
    .Y(n_9739));
 XNOR2x1_ASAP7_75t_SL g18550 (.B(n_7801),
    .Y(n_9740),
    .A(n_7800));
 AOI21x1_ASAP7_75t_SL g18551 (.A1(n_20078),
    .A2(n_9744),
    .B(n_9745),
    .Y(n_9746));
 NAND2x1p5_ASAP7_75t_SL g18553 (.A(n_9743),
    .B(n_4193),
    .Y(n_9744));
 HB1xp67_ASAP7_75t_SL g18554 (.A(n_21293),
    .Y(n_9743));
 AND2x2_ASAP7_75t_SL g18555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_249),
    .Y(n_9745));
 XNOR2x1_ASAP7_75t_SL g18556 (.B(n_19160),
    .Y(n_9750),
    .A(n_9747));
 AND2x2_ASAP7_75t_SL g18557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_46),
    .Y(n_9747));
 OAI21x1_ASAP7_75t_SL g18560 (.A1(n_9751),
    .A2(n_9754),
    .B(n_9755),
    .Y(n_9756));
 NAND2xp67_ASAP7_75t_SL g18561 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_53),
    .Y(n_9751));
 AND2x2_ASAP7_75t_SL g18562 (.A(n_9752),
    .B(n_9753),
    .Y(n_9754));
 NAND2xp5_ASAP7_75t_L g18563 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .Y(n_9752));
 NAND2x1_ASAP7_75t_SL g18564 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_2392),
    .Y(n_9753));
 OR2x2_ASAP7_75t_SL g18565 (.A(n_9752),
    .B(n_9753),
    .Y(n_9755));
 NAND2xp5_ASAP7_75t_SL g18567 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .B(n_3528),
    .Y(n_9757));
 INVxp67_ASAP7_75t_SL g18569 (.A(n_9759),
    .Y(n_4044));
 NAND2xp5_ASAP7_75t_SL g18570 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .Y(n_9759));
 NAND2x1p5_ASAP7_75t_SL g18572 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .B(n_2825),
    .Y(n_9762));
 AND2x2_ASAP7_75t_SL g18573 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .Y(n_9763));
 XNOR2x1_ASAP7_75t_SL g18598 (.B(n_9793),
    .Y(n_9794),
    .A(n_9792));
 NAND2x1_ASAP7_75t_SL g18599 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_648),
    .B(n_2180),
    .Y(n_9792));
 AND2x2_ASAP7_75t_SL g18600 (.A(n_2176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_616),
    .Y(n_9793));
 NAND2x1p5_ASAP7_75t_SL g18603 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113));
 MAJIxp5_ASAP7_75t_SL g18604 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_0),
    .Y(n_9797));
 INVx1_ASAP7_75t_SL g18605 (.A(n_9797),
    .Y(n_9799));
 AO21x1_ASAP7_75t_SL g18608 (.A1(n_7778),
    .A2(n_7775),
    .B(n_7784),
    .Y(n_9801));
 AOI21xp5_ASAP7_75t_SL g18611 (.A1(n_9806),
    .A2(n_9805),
    .B(n_9807),
    .Y(n_9808));
 OAI21x1_ASAP7_75t_SL g18612 (.A1(n_7109),
    .A2(n_22431),
    .B(n_7111),
    .Y(n_9805));
 NAND2xp5_ASAP7_75t_SL g18613 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_191),
    .Y(n_9806));
 NOR2xp33_ASAP7_75t_SL g18614 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_191),
    .Y(n_9807));
 NAND2xp5_ASAP7_75t_SL g18615 (.A(n_4275),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .Y(n_9810));
 AND2x2_ASAP7_75t_SL g18619 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_674),
    .B(n_2160),
    .Y(n_9811));
 INVx1_ASAP7_75t_SL g18620 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_579),
    .Y(n_9813));
 INVx1_ASAP7_75t_SL g18624 (.A(n_19408),
    .Y(n_9818));
 XNOR2xp5_ASAP7_75t_SL g18625 (.A(n_9819),
    .B(n_9820),
    .Y(n_9821));
 AND2x2_ASAP7_75t_SL g18626 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_54),
    .Y(n_9819));
 OAI22xp5_ASAP7_75t_SL g18627 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_76),
    .A2(n_3239),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_77),
    .Y(n_9820));
 MAJIxp5_ASAP7_75t_SL g18635 (.A(n_9828),
    .B(n_9829),
    .C(n_9830),
    .Y(n_9831));
 INVx1_ASAP7_75t_SL g18636 (.A(n_21134),
    .Y(n_9828));
 INVxp67_ASAP7_75t_SL g18637 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .Y(n_9829));
 INVxp67_ASAP7_75t_SL g18638 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_291),
    .Y(n_9830));
 INVx1_ASAP7_75t_SL g18640 (.A(n_9827),
    .Y(n_9833));
 XNOR2xp5_ASAP7_75t_SL g18643 (.A(n_22950),
    .B(n_9840),
    .Y(n_9841));
 XNOR2xp5_ASAP7_75t_SL g18645 (.A(n_7338),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_13),
    .Y(n_9840));
 NAND2xp5_ASAP7_75t_SL g18648 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .Y(n_9842));
 INVx1_ASAP7_75t_SL g18652 (.A(n_14781),
    .Y(n_9848));
 OAI22xp5_ASAP7_75t_SL g18654 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_110),
    .A2(n_14783),
    .B1(n_14786),
    .B2(n_14784),
    .Y(n_9849));
 XNOR2x1_ASAP7_75t_SL g18663 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_4),
    .Y(n_9860),
    .A(n_9859));
 BUFx2_ASAP7_75t_SL g18664 (.A(n_22617),
    .Y(n_9859));
 XNOR2x1_ASAP7_75t_SL g18665 (.B(n_18760),
    .Y(n_9862),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_133));
 NOR2xp67_ASAP7_75t_SL g18669 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_247),
    .Y(n_9865));
 NAND2xp5_ASAP7_75t_SL g18670 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_247),
    .Y(n_9866));
 INVx1_ASAP7_75t_SL g18677 (.A(n_12786),
    .Y(n_9874));
 OAI21xp5_ASAP7_75t_SL g18678 (.A1(n_19282),
    .A2(n_15079),
    .B(n_9879),
    .Y(n_9880));
 OAI21xp5_ASAP7_75t_SL g18684 (.A1(n_9881),
    .A2(n_9882),
    .B(n_9883),
    .Y(n_9884));
 NOR2xp33_ASAP7_75t_SL g18685 (.A(n_22040),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_198),
    .Y(n_9881));
 OAI21xp5_ASAP7_75t_SL g18686 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_181),
    .A2(n_21210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_201),
    .Y(n_9882));
 NAND2xp5_ASAP7_75t_SL g18687 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_181),
    .B(n_21210),
    .Y(n_9883));
 XOR2xp5_ASAP7_75t_SL g18694 (.A(n_20164),
    .B(n_9892),
    .Y(n_9893));
 NAND2xp5_ASAP7_75t_SL g18696 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_648),
    .B(n_9662),
    .Y(n_9892));
 OAI21xp5_ASAP7_75t_SL g18699 (.A1(n_9898),
    .A2(n_9899),
    .B(n_9902),
    .Y(n_9903));
 INVx1_ASAP7_75t_SL g187 (.A(n_22252),
    .Y(n_21419));
 NAND2xp5_ASAP7_75t_SL g18700 (.A(n_9897),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_310),
    .Y(n_9898));
 INVxp67_ASAP7_75t_SL g18701 (.A(n_9896),
    .Y(n_9897));
 NOR2xp33_ASAP7_75t_SL g18702 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_249),
    .Y(n_9896));
 INVxp67_ASAP7_75t_SL g18703 (.A(n_20347),
    .Y(n_9899));
 AOI21xp33_ASAP7_75t_SL g18704 (.A1(n_23032),
    .A2(n_9897),
    .B(n_7908),
    .Y(n_9902));
 NAND2xp5_ASAP7_75t_SL g18706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_249),
    .Y(n_9900));
 AOI21xp5_ASAP7_75t_SL g18707 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_310),
    .A2(n_20347),
    .B(n_23032),
    .Y(n_9904));
 OAI22xp5_ASAP7_75t_SL g18708 (.A1(n_9908),
    .A2(n_3873),
    .B1(n_9905),
    .B2(n_22953),
    .Y(n_3450));
 NAND2xp5_ASAP7_75t_SL g18709 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .Y(n_9905));
 INVx1_ASAP7_75t_SL g18711 (.A(n_3868),
    .Y(n_3873));
 NAND2xp5_ASAP7_75t_SL g18713 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(n_3868),
    .Y(n_9912));
 OAI21x1_ASAP7_75t_SL g18722 (.A1(n_9922),
    .A2(n_9923),
    .B(n_12748),
    .Y(n_9925));
 NOR2xp33_ASAP7_75t_SL g18723 (.A(n_18761),
    .B(n_21476),
    .Y(n_9922));
 AND2x2_ASAP7_75t_SL g18725 (.A(n_21476),
    .B(n_18761),
    .Y(n_9923));
 XNOR2xp5_ASAP7_75t_SL g18727 (.A(n_9927),
    .B(n_9928),
    .Y(n_9929));
 INVxp67_ASAP7_75t_SL g18728 (.A(n_9926),
    .Y(n_9927));
 NOR2xp67_ASAP7_75t_SL g18729 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_46),
    .B(n_12120),
    .Y(n_9926));
 AOI22xp5_ASAP7_75t_SL g18730 (.A1(n_13711),
    .A2(n_5423),
    .B1(n_5422),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_95),
    .Y(n_9928));
 INVx1_ASAP7_75t_SL g18753 (.A(n_9776),
    .Y(n_9950));
 AOI21xp5_ASAP7_75t_SL g18756 (.A1(n_22429),
    .A2(n_9695),
    .B(n_9698),
    .Y(n_9957));
 NOR2x1_ASAP7_75t_SL g18758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_268),
    .B(n_14417),
    .Y(n_9959));
 NAND2xp5_ASAP7_75t_SL g18760 (.A(n_14417),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_268),
    .Y(n_9961));
 INVxp67_ASAP7_75t_SRAM g18761 (.A(n_13061),
    .Y(n_9963));
 XNOR2xp5_ASAP7_75t_SL g18770 (.A(n_9971),
    .B(n_19599),
    .Y(n_9972));
 XOR2x2_ASAP7_75t_SL g18771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_265),
    .Y(n_9971));
 MAJIxp5_ASAP7_75t_SL g18772 (.A(n_9971),
    .B(n_8191),
    .C(n_8194),
    .Y(n_9973));
 NAND2xp5_ASAP7_75t_SL g18774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_399),
    .B(n_20111),
    .Y(n_9974));
 NAND2xp33_ASAP7_75t_SL g18776 (.A(n_9974),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_430),
    .Y(n_9977));
 NAND2xp5_ASAP7_75t_SL g18783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .B(n_9985),
    .Y(n_9986));
 NAND2xp5_ASAP7_75t_SL g18784 (.A(n_14122),
    .B(n_10091),
    .Y(n_9985));
 OAI21xp5_ASAP7_75t_SL g18785 (.A1(n_9627),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .B(n_9985),
    .Y(n_9987));
 NAND2xp33_ASAP7_75t_R g18786 (.A(n_9985),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_430),
    .Y(n_9988));
 AND2x2_ASAP7_75t_SL g18787 (.A(n_9990),
    .B(n_11611),
    .Y(n_9991));
 XNOR2xp5_ASAP7_75t_SL g18788 (.A(n_9989),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_247),
    .Y(n_9990));
 INVx1_ASAP7_75t_SL g18789 (.A(n_20134),
    .Y(n_9989));
 OR2x2_ASAP7_75t_SL g18790 (.A(n_11611),
    .B(n_9990),
    .Y(n_9992));
 XNOR2x1_ASAP7_75t_SL g18796 (.B(n_15077),
    .Y(n_9997),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_65));
 XNOR2xp5_ASAP7_75t_SL g188 (.A(n_11537),
    .B(n_11538),
    .Y(n_11539));
 HB1xp67_ASAP7_75t_SL g18803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_37),
    .Y(n_10005));
 XNOR2xp5_ASAP7_75t_SL g18804 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_137),
    .B(n_18941),
    .Y(n_10009));
 MAJIxp5_ASAP7_75t_SL g18808 (.A(n_10012),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_164),
    .Y(n_10013));
 XOR2xp5_ASAP7_75t_SL g18812 (.A(n_10012),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_195),
    .Y(n_10014));
 MAJIxp5_ASAP7_75t_SL g18827 (.A(n_8653),
    .B(n_10029),
    .C(n_10032),
    .Y(n_10033));
 OAI21xp33_ASAP7_75t_SL g18833 (.A1(n_22955),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_282),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_291),
    .Y(n_10038));
 XOR2xp5_ASAP7_75t_L g18836 (.A(n_22955),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_297),
    .Y(n_10039));
 XNOR2xp5_ASAP7_75t_SL g18839 (.A(n_12038),
    .B(n_3652),
    .Y(n_10044));
 XOR2xp5_ASAP7_75t_SL g18842 (.A(n_14117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_56),
    .Y(n_10046));
 AOI21xp5_ASAP7_75t_SL g18850 (.A1(n_10912),
    .A2(n_17869),
    .B(n_10053),
    .Y(n_10054));
 AND2x2_ASAP7_75t_SL g18851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[16]),
    .B(n_17870),
    .Y(n_10053));
 OAI21xp5_ASAP7_75t_SL g18852 (.A1(n_4084),
    .A2(n_10055),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_277),
    .Y(n_10056));
 AOI21xp5_ASAP7_75t_SL g18853 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_278),
    .A2(n_21401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_281),
    .Y(n_10055));
 XOR2xp5_ASAP7_75t_L g18854 (.A(n_10055),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_285),
    .Y(n_10057));
 XOR2xp5_ASAP7_75t_SL g18865 (.A(n_10068),
    .B(n_3450),
    .Y(n_10069));
 XNOR2xp5_ASAP7_75t_SL g18866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_108),
    .B(n_25337),
    .Y(n_10068));
 MAJIxp5_ASAP7_75t_SL g18867 (.A(n_19964),
    .B(n_3450),
    .C(n_10070),
    .Y(n_10071));
 HB1xp67_ASAP7_75t_SL g18868 (.A(n_10068),
    .Y(n_10070));
 NAND2x1p5_ASAP7_75t_SL g18871 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_63),
    .Y(n_10073));
 MAJIxp5_ASAP7_75t_SL g18873 (.A(n_19718),
    .B(n_10073),
    .C(n_19714),
    .Y(n_10078));
 OAI21xp5_ASAP7_75t_SL g18878 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_206),
    .A2(n_10082),
    .B(n_10084),
    .Y(n_10085));
 XOR2xp5_ASAP7_75t_SL g18879 (.A(n_10081),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_182),
    .Y(n_10082));
 INVxp67_ASAP7_75t_SL g18880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_157),
    .Y(n_10081));
 NAND2xp5_ASAP7_75t_SL g18881 (.A(n_10083),
    .B(n_10082),
    .Y(n_10084));
 INVxp67_ASAP7_75t_SL g18882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_205),
    .Y(n_10083));
 INVxp67_ASAP7_75t_SL g18884 (.A(n_10082),
    .Y(n_10086));
 XNOR2xp5_ASAP7_75t_SL g18885 (.A(n_22540),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_350),
    .Y(n_10090));
 MAJIxp5_ASAP7_75t_SL g18888 (.A(n_22540),
    .B(n_20357),
    .C(n_20719),
    .Y(n_10091));
 MAJIxp5_ASAP7_75t_SL g18889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_228),
    .B(n_10093),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_174),
    .Y(n_10094));
 HB1xp67_ASAP7_75t_SL g18890 (.A(n_10092),
    .Y(n_10093));
 XNOR2xp5_ASAP7_75t_SL g18891 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_127),
    .Y(n_10092));
 OAI22xp5_ASAP7_75t_SL g18894 (.A1(n_10097),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_48),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_47),
    .B2(n_10098),
    .Y(n_10099));
 NAND2xp5_ASAP7_75t_SL g18895 (.A(n_4826),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .Y(n_10097));
 INVx1_ASAP7_75t_SL g18896 (.A(n_10097),
    .Y(n_10098));
 MAJIxp5_ASAP7_75t_SL g18897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_49),
    .C(n_10097),
    .Y(n_10100));
 XNOR2xp5_ASAP7_75t_SL g18898 (.A(n_22825),
    .B(n_7994),
    .Y(n_10102));
 XOR2x1_ASAP7_75t_SL g188_0 (.A(n_6667),
    .Y(n_6669),
    .B(n_6668));
 INVxp67_ASAP7_75t_SL g18900 (.A(n_22825),
    .Y(n_10103));
 XOR2xp5_ASAP7_75t_SL g18901 (.A(n_14732),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_257),
    .Y(n_10106));
 XNOR2xp5_ASAP7_75t_SL g18910 (.A(n_10114),
    .B(n_10116),
    .Y(n_10117));
 INVx1_ASAP7_75t_SL g18911 (.A(n_11072),
    .Y(n_10114));
 XNOR2xp5_ASAP7_75t_SL g18912 (.A(n_10115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_36),
    .Y(n_10116));
 INVx1_ASAP7_75t_SL g18913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_190),
    .Y(n_10115));
 AND2x2_ASAP7_75t_SL g18919 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .Y(n_10122));
 INVxp67_ASAP7_75t_SL g18923 (.A(n_10122),
    .Y(n_10125));
 XNOR2xp5_ASAP7_75t_SL g18924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_204),
    .B(n_10128),
    .Y(n_10129));
 MAJIxp5_ASAP7_75t_SL g18925 (.A(n_7575),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_156),
    .Y(n_10128));
 NOR2xp33_ASAP7_75t_SL g18926 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_205),
    .B(n_10128),
    .Y(n_10130));
 NAND2xp33_ASAP7_75t_SL g18927 (.A(n_10128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_205),
    .Y(n_10131));
 A2O1A1Ixp33_ASAP7_75t_SL g18932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_259),
    .A2(n_10136),
    .B(n_10137),
    .C(n_10138),
    .Y(n_10139));
 OR2x2_ASAP7_75t_SL g18934 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_261),
    .Y(n_10137));
 OR2x2_ASAP7_75t_SL g18935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_189),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_183),
    .Y(n_10138));
 OAI22xp5_ASAP7_75t_SL g18936 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_257),
    .A2(n_10136),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_258),
    .B2(n_16564),
    .Y(n_10141));
 INVx2_ASAP7_75t_SL g18937 (.A(n_16564),
    .Y(n_10136));
 XNOR2xp5_ASAP7_75t_SL g18938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_126),
    .B(n_10142),
    .Y(n_10143));
 XNOR2xp5_ASAP7_75t_SL g18939 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_717),
    .B(n_18581),
    .Y(n_10142));
 MAJIxp5_ASAP7_75t_SL g18940 (.A(n_10142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_126),
    .C(n_11295),
    .Y(n_10144));
 MAJIxp5_ASAP7_75t_SL g18947 (.A(n_21869),
    .B(n_21864),
    .C(n_21862),
    .Y(n_10153));
 XOR2xp5_ASAP7_75t_SL g18955 (.A(n_10157),
    .B(n_20076),
    .Y(n_10159));
 NAND2xp5_ASAP7_75t_SL g18956 (.A(n_22482),
    .B(n_19575),
    .Y(n_10161));
 NOR2xp67_ASAP7_75t_SL g18958 (.A(n_22482),
    .B(n_19575),
    .Y(n_10162));
 NAND2x1_ASAP7_75t_SL g18960 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(n_9349),
    .Y(n_10163));
 XOR2xp5_ASAP7_75t_SL g18964 (.A(n_11374),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_240),
    .Y(n_10171));
 INVx1_ASAP7_75t_SL g18966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .Y(n_10169));
 MAJx2_ASAP7_75t_SL g18967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_32),
    .B(n_10172),
    .C(n_10176),
    .Y(n_10177));
 HB1xp67_ASAP7_75t_SL g18968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .Y(n_10172));
 OAI22xp5_ASAP7_75t_SL g18969 (.A1(n_10173),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_240),
    .B1(n_10174),
    .B2(n_10175),
    .Y(n_10176));
 INVx1_ASAP7_75t_SL g18970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_240),
    .Y(n_10175));
 OAI21xp5_ASAP7_75t_SL g18973 (.A1(n_10180),
    .A2(n_10182),
    .B(n_23066),
    .Y(n_10185));
 INVx2_ASAP7_75t_SL g18974 (.A(n_14689),
    .Y(n_10180));
 NAND2xp5_ASAP7_75t_SL g18975 (.A(n_10181),
    .B(n_23054),
    .Y(n_10182));
 INVxp67_ASAP7_75t_SL g18976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_273),
    .Y(n_10181));
 INVx1_ASAP7_75t_SL g18978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_274));
 NOR2xp33_ASAP7_75t_SL g18980 (.A(n_10187),
    .B(n_20501),
    .Y(n_10188));
 NOR2x1_ASAP7_75t_SL g18981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_264),
    .B(n_8214),
    .Y(n_10187));
 AOI21x1_ASAP7_75t_SL g18988 (.A1(n_10195),
    .A2(n_18948),
    .B(n_18797),
    .Y(n_10200));
 NAND2xp5_ASAP7_75t_SL g18989 (.A(n_9617),
    .B(n_9618),
    .Y(n_10195));
 NAND3xp33_ASAP7_75t_SL g18995 (.A(n_18797),
    .B(n_18948),
    .C(n_10195),
    .Y(n_10202));
 OAI21xp5_ASAP7_75t_SL g18996 (.A1(n_16156),
    .A2(n_16155),
    .B(n_18954),
    .Y(n_10205));
 OAI21x1_ASAP7_75t_SL g19 (.A1(n_10762),
    .A2(n_21962),
    .B(n_2160),
    .Y(n_21963));
 XNOR2x1_ASAP7_75t_SL g190 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_192),
    .Y(n_6097),
    .A(n_9094));
 HB1xp67_ASAP7_75t_SL g19001 (.A(n_22881),
    .Y(n_10208));
 XNOR2xp5_ASAP7_75t_SL g19002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_137),
    .B(n_18949),
    .Y(n_10212));
 XNOR2xp5_ASAP7_75t_SL g19010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_238),
    .B(n_19663),
    .Y(n_10220));
 MAJIxp5_ASAP7_75t_SL g19015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_149),
    .B(n_12528),
    .C(n_10224),
    .Y(n_10225));
 XNOR2x1_ASAP7_75t_SL g19018 (.B(n_15795),
    .Y(n_10224),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_6));
 OAI21x1_ASAP7_75t_SL g19027 (.A1(n_23564),
    .A2(n_10234),
    .B(n_23566),
    .Y(n_10235));
 XNOR2x1_ASAP7_75t_SL g19028 (.B(n_21143),
    .Y(n_10234),
    .A(n_7041));
 XNOR2xp5_ASAP7_75t_SL g19029 (.A(n_23568),
    .B(n_10234),
    .Y(n_10236));
 INVxp67_ASAP7_75t_SL g19031 (.A(n_10239),
    .Y(n_10240));
 NOR2xp33_ASAP7_75t_SL g19032 (.A(n_10238),
    .B(n_12108),
    .Y(n_10239));
 NAND2xp5_ASAP7_75t_SL g19033 (.A(n_2173),
    .B(n_10237),
    .Y(n_10238));
 AOI21xp33_ASAP7_75t_SL g19034 (.A1(n_10241),
    .A2(n_10239),
    .B(n_10242),
    .Y(n_10243));
 INVxp67_ASAP7_75t_SL g19035 (.A(n_12107),
    .Y(n_10241));
 NOR2xp33_ASAP7_75t_SL g19036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_211),
    .B(n_10238),
    .Y(n_10242));
 NOR2xp33_ASAP7_75t_R g19040 (.A(n_16326),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_235),
    .Y(n_10248));
 OAI22xp5_ASAP7_75t_SL g19046 (.A1(n_10256),
    .A2(n_10260),
    .B1(n_22596),
    .B2(n_10261),
    .Y(n_10262));
 NAND2xp5_ASAP7_75t_SL g19047 (.A(n_2182),
    .B(n_10255),
    .Y(n_10256));
 INVxp67_ASAP7_75t_SL g19048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_213),
    .Y(n_10255));
 AOI21xp5_ASAP7_75t_SL g19049 (.A1(n_10257),
    .A2(n_10258),
    .B(n_18763),
    .Y(n_10260));
 INVxp67_ASAP7_75t_SL g19050 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_298),
    .Y(n_10257));
 INVx1_ASAP7_75t_SL g19051 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_301),
    .Y(n_10258));
 XNOR2xp5_ASAP7_75t_SL g19052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_357),
    .B(n_10263),
    .Y(n_10264));
 XOR2x1_ASAP7_75t_SL g19053 (.A(n_24770),
    .Y(n_10263),
    .B(n_9215));
 OAI21xp5_ASAP7_75t_SL g19054 (.A1(n_10263),
    .A2(n_10265),
    .B(n_10266),
    .Y(n_10267));
 NOR2xp33_ASAP7_75t_SL g19055 (.A(n_11246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_257),
    .Y(n_10265));
 NAND2xp33_ASAP7_75t_L g19056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_257),
    .B(n_11246),
    .Y(n_10266));
 XNOR2xp5_ASAP7_75t_SL g19057 (.A(n_18764),
    .B(n_20988),
    .Y(n_10271));
 OAI21x1_ASAP7_75t_SL g19061 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_188),
    .A2(n_10272),
    .B(n_11808),
    .Y(n_10274));
 NOR2xp33_ASAP7_75t_SL g19062 (.A(n_18764),
    .B(n_20988),
    .Y(n_10272));
 MAJIxp5_ASAP7_75t_SL g19064 (.A(n_18144),
    .B(n_10276),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_174),
    .Y(n_10278));
 XOR2xp5_ASAP7_75t_SL g19066 (.A(n_25999),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_127),
    .Y(n_10276));
 XNOR2xp5_ASAP7_75t_SL g19068 (.A(n_10279),
    .B(n_10276),
    .Y(n_10280));
 INVx1_ASAP7_75t_SL g19069 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_174),
    .Y(n_10279));
 XNOR2xp5_ASAP7_75t_SL g19071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_106),
    .B(n_13242),
    .Y(n_10281));
 XNOR2xp5_ASAP7_75t_SL g19072 (.A(n_10281),
    .B(n_4904),
    .Y(n_10283));
 MAJIxp5_ASAP7_75t_SL g19074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_305),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .Y(n_10284));
 INVx1_ASAP7_75t_SL g19076 (.A(n_10284),
    .Y(n_10286));
 NAND2xp5_ASAP7_75t_SL g19077 (.A(n_12283),
    .B(n_10286),
    .Y(n_10290));
 OAI211xp5_ASAP7_75t_SL g19080 (.A1(n_9238),
    .A2(n_11891),
    .B(n_12284),
    .C(n_10284),
    .Y(n_10291));
 XOR2xp5_ASAP7_75t_SL g19083 (.A(n_9162),
    .B(n_18942),
    .Y(n_10294));
 MAJIxp5_ASAP7_75t_SL g19084 (.A(n_24751),
    .B(n_24752),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_35),
    .Y(n_10295));
 INVxp67_ASAP7_75t_SL g19086 (.A(n_10295),
    .Y(n_10298));
 AOI22xp5_ASAP7_75t_SL g19089 (.A1(n_9389),
    .A2(n_10301),
    .B1(n_10302),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_163),
    .Y(n_10303));
 INVx1_ASAP7_75t_SL g19090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_163),
    .Y(n_10301));
 MAJIxp5_ASAP7_75t_SL g19092 (.A(n_10305),
    .B(n_4248),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_115),
    .Y(n_10307));
 XOR2xp5_ASAP7_75t_SL g19094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_142),
    .Y(n_10305));
 OAI21xp5_ASAP7_75t_SL g19096 (.A1(n_10309),
    .A2(n_21361),
    .B(n_15886),
    .Y(n_10311));
 OAI22xp5_ASAP7_75t_SL g191 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_286),
    .A2(n_22797),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_287),
    .B2(n_22796),
    .Y(n_22806));
 OAI22xp5_ASAP7_75t_SL g19104 (.A1(n_10325),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_149),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_4),
    .B2(n_10324),
    .Y(n_10326));
 INVx1_ASAP7_75t_SL g19105 (.A(n_10324),
    .Y(n_10325));
 NOR2x1_ASAP7_75t_SL g19106 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_64),
    .Y(n_10324));
 MAJIxp5_ASAP7_75t_SL g19107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_4),
    .B(n_10325),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_157),
    .Y(n_10327));
 AOI21xp5_ASAP7_75t_SL g19108 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_n_186),
    .A2(n_23932),
    .B(n_10328),
    .Y(n_10329));
 AND2x2_ASAP7_75t_SL g19109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[16]),
    .B(n_17882),
    .Y(n_10328));
 XNOR2xp5_ASAP7_75t_SL g19113 (.A(n_7330),
    .B(n_10333),
    .Y(n_10334));
 OAI22xp5_ASAP7_75t_SL g19114 (.A1(n_7328),
    .A2(n_7327),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_75),
    .B2(n_7326),
    .Y(n_10333));
 NAND2xp5_ASAP7_75t_SL g19119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_400),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_362),
    .Y(n_10338));
 INVxp67_ASAP7_75t_SL g19122 (.A(n_10338),
    .Y(n_10340));
 NAND2xp5_ASAP7_75t_SL g19125 (.A(n_16757),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .Y(n_10344));
 MAJIxp5_ASAP7_75t_SL g19126 (.A(n_10344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_49),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_40),
    .Y(n_10346));
 AND2x2_ASAP7_75t_SL g19127 (.A(n_13448),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_265),
    .Y(n_10348));
 NOR2xp67_ASAP7_75t_SL g19129 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_265),
    .B(n_13448),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_290));
 NAND2x1_ASAP7_75t_SL g19131 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_100),
    .Y(n_10350));
 MAJIxp5_ASAP7_75t_SL g19133 (.A(n_7726),
    .B(n_10350),
    .C(n_10719),
    .Y(n_10355));
 MAJx2_ASAP7_75t_SL g19136 (.A(n_7997),
    .B(n_7996),
    .C(n_7399),
    .Y(n_10356));
 XNOR2xp5_ASAP7_75t_SL g19138 (.A(n_9160),
    .B(n_10359),
    .Y(n_10360));
 AOI22xp5_ASAP7_75t_SL g19139 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_101),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_93),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_102),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_94),
    .Y(n_10359));
 XOR2xp5_ASAP7_75t_SL g19147 (.A(n_21541),
    .B(n_10368),
    .Y(n_10369));
 INVxp67_ASAP7_75t_SL g19148 (.A(n_21826),
    .Y(n_10368));
 OAI22xp5_ASAP7_75t_SL g19150 (.A1(n_9042),
    .A2(n_2940),
    .B1(n_22463),
    .B2(n_3548),
    .Y(n_10370));
 OAI22xp33_ASAP7_75t_SL g19153 (.A1(n_23555),
    .A2(n_10374),
    .B1(n_10375),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_171),
    .Y(n_10376));
 INVxp67_ASAP7_75t_SL g19154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_171),
    .Y(n_10374));
 INVx1_ASAP7_75t_SL g19155 (.A(n_23555),
    .Y(n_10375));
 AO21x1_ASAP7_75t_SRAM g19156 (.A1(n_23000),
    .A2(n_6527),
    .B(n_6528),
    .Y(n_10378));
 XNOR2xp5_ASAP7_75t_SL g19158 (.A(n_6519),
    .B(n_23000),
    .Y(n_10379));
 INVxp67_ASAP7_75t_SL g19169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_5),
    .Y(n_10389));
 XOR2xp5_ASAP7_75t_SL g19170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_34),
    .B(n_26074),
    .Y(n_10393));
 MAJx2_ASAP7_75t_SL g19173 (.A(n_2901),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .C(n_10394),
    .Y(n_10395));
 INVx1_ASAP7_75t_SL g19174 (.A(n_26074),
    .Y(n_10394));
 MAJIxp5_ASAP7_75t_SL g19188 (.A(n_6327),
    .B(n_6331),
    .C(n_6329),
    .Y(n_10408));
 INVxp67_ASAP7_75t_SL g19191 (.A(n_10408),
    .Y(n_10411));
 XNOR2xp5_ASAP7_75t_SL g19192 (.A(n_18766),
    .B(n_20141),
    .Y(n_10416));
 INVx1_ASAP7_75t_SL g19195 (.A(n_19131),
    .Y(n_10414));
 XOR2x2_ASAP7_75t_SL g19197 (.A(n_26169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_265),
    .Y(n_10417));
 XNOR2xp5_ASAP7_75t_SL g19198 (.A(n_10417),
    .B(n_22977),
    .Y(n_10419));
 MAJIxp5_ASAP7_75t_SL g192 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_192),
    .B(n_6098),
    .C(n_6099),
    .Y(n_6100));
 NAND2xp5_ASAP7_75t_SL g19201 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .Y(n_10421));
 XNOR2xp5_ASAP7_75t_SL g19202 (.A(n_10421),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_37),
    .Y(n_10423));
 NOR2xp67_ASAP7_75t_SL g19207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_262),
    .B(n_13487),
    .Y(n_10427));
 AOI21xp5_ASAP7_75t_SL g19208 (.A1(n_10427),
    .A2(n_21364),
    .B(n_18753),
    .Y(n_10429));
 NOR2xp33_ASAP7_75t_SRAM g19221 (.A(n_10442),
    .B(n_9776),
    .Y(n_10443));
 NOR2xp33_ASAP7_75t_SL g19222 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_236),
    .B(n_11388),
    .Y(n_10442));
 OA21x2_ASAP7_75t_SL g19223 (.A1(n_10444),
    .A2(n_11124),
    .B(n_11126),
    .Y(n_10445));
 INVxp67_ASAP7_75t_SL g19224 (.A(n_10442),
    .Y(n_10444));
 HB1xp67_ASAP7_75t_SL g19226 (.A(n_10444),
    .Y(n_10446));
 AOI21xp5_ASAP7_75t_SL g19233 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .A2(n_16319),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_475),
    .Y(n_10455));
 INVx1_ASAP7_75t_SL g19237 (.A(n_8492),
    .Y(n_10456));
 INVxp67_ASAP7_75t_SL g19244 (.A(n_10465),
    .Y(n_10466));
 XNOR2xp5_ASAP7_75t_SL g19245 (.A(n_9183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_164),
    .Y(n_10465));
 MAJIxp5_ASAP7_75t_SL g19247 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_77),
    .B(n_10469),
    .C(n_6932),
    .Y(n_10470));
 OR2x2_ASAP7_75t_SL g19248 (.A(n_14372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_46),
    .Y(n_10469));
 XOR2x2_ASAP7_75t_SL g19249 (.A(n_10469),
    .B(n_18812),
    .Y(n_10471));
 XNOR2xp5_ASAP7_75t_SL g19251 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_234),
    .B(n_10370),
    .Y(n_10472));
 XNOR2xp5_ASAP7_75t_SL g19253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_300),
    .B(n_10477),
    .Y(n_10478));
 AOI21x1_ASAP7_75t_SL g19254 (.A1(n_13603),
    .A2(n_10475),
    .B(n_10476),
    .Y(n_10477));
 HB1xp67_ASAP7_75t_SL g19256 (.A(n_15816),
    .Y(n_10476));
 OAI21xp33_ASAP7_75t_SL g19257 (.A1(n_10477),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_297),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_295),
    .Y(n_10479));
 OAI21xp5_ASAP7_75t_SL g19258 (.A1(n_6958),
    .A2(n_10480),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_229),
    .Y(n_10481));
 NOR2xp33_ASAP7_75t_SL g19259 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_216),
    .Y(n_10480));
 OAI21xp33_ASAP7_75t_SL g19260 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_216),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_229),
    .Y(n_10482));
 XOR2x2_ASAP7_75t_SL g19262 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_265),
    .Y(n_10483));
 XNOR2xp5_ASAP7_75t_SL g19277 (.A(n_10500),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_240),
    .Y(n_10501));
 XNOR2x2_ASAP7_75t_SL g19278 (.A(n_10499),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_3),
    .Y(n_10500));
 INVxp67_ASAP7_75t_SL g19279 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_753),
    .Y(n_10499));
 OAI22xp5_ASAP7_75t_SL g19280 (.A1(n_19170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_195),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_145),
    .B2(n_10500),
    .Y(n_10505));
 NAND2xp5_ASAP7_75t_SL g19283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_753),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_3),
    .Y(n_10503));
 NAND2xp5_ASAP7_75t_SL g19286 (.A(n_2176),
    .B(n_9808),
    .Y(n_10506));
 XOR2x2_ASAP7_75t_SL g19289 (.A(n_19869),
    .B(n_18157),
    .Y(n_10509));
 MAJIxp5_ASAP7_75t_SL g19290 (.A(n_10509),
    .B(n_23392),
    .C(n_6079),
    .Y(n_10512));
 XNOR2xp5_ASAP7_75t_SL g19292 (.A(n_7604),
    .B(n_7610),
    .Y(n_10513));
 NOR2xp67_ASAP7_75t_SL g19293 (.A(n_6833),
    .B(n_10513),
    .Y(n_10515));
 XOR2xp5_ASAP7_75t_SL g19295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_85),
    .Y(n_10516));
 AO21x2_ASAP7_75t_SL g19299 (.A1(n_10516),
    .A2(n_10521),
    .B(n_10522),
    .Y(n_10523));
 INVxp67_ASAP7_75t_SL g193 (.A(n_9091),
    .Y(n_6098));
 NAND2xp33_ASAP7_75t_SL g19300 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_108),
    .Y(n_10521));
 NOR2xp33_ASAP7_75t_SL g19301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_115),
    .Y(n_10522));
 INVx1_ASAP7_75t_SL g19307 (.A(n_8959),
    .Y(n_10527));
 MAJIxp5_ASAP7_75t_SL g19311 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_237),
    .B(n_10532),
    .C(n_7460),
    .Y(n_10533));
 HB1xp67_ASAP7_75t_SL g19312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_206),
    .Y(n_10532));
 XNOR2xp5_ASAP7_75t_SL g19314 (.A(n_10537),
    .B(n_5473),
    .Y(n_10538));
 NOR2xp33_ASAP7_75t_SL g19315 (.A(n_10536),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_303),
    .Y(n_10537));
 HB1xp67_ASAP7_75t_SL g19316 (.A(n_7618),
    .Y(n_10536));
 XOR2xp5_ASAP7_75t_SL g19319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_262),
    .B(n_10542),
    .Y(n_10543));
 HB1xp67_ASAP7_75t_SL g19320 (.A(n_10541),
    .Y(n_10542));
 AOI21xp5_ASAP7_75t_SL g19321 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_230),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_228),
    .Y(n_10541));
 OAI21xp5_ASAP7_75t_SL g19322 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_252),
    .A2(n_10541),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_254),
    .Y(n_10544));
 NOR2x1_ASAP7_75t_SL g19334 (.A(n_10557),
    .B(n_10560),
    .Y(n_10561));
 INVxp67_ASAP7_75t_SL g19335 (.A(n_11324),
    .Y(n_10557));
 AOI22xp5_ASAP7_75t_SL g19336 (.A1(n_10558),
    .A2(n_11788),
    .B1(n_23450),
    .B2(n_11789),
    .Y(n_10560));
 INVx1_ASAP7_75t_L g19337 (.A(n_23450),
    .Y(n_10558));
 OAI22xp5_ASAP7_75t_SL g19340 (.A1(n_10563),
    .A2(n_7724),
    .B1(n_10564),
    .B2(n_7721),
    .Y(n_9917));
 XNOR2xp5_ASAP7_75t_SL g19341 (.A(n_7502),
    .B(n_7495),
    .Y(n_10563));
 INVx1_ASAP7_75t_SL g19342 (.A(n_10563),
    .Y(n_10564));
 OAI21x1_ASAP7_75t_SL g19344 (.A1(n_7724),
    .A2(n_10567),
    .B(n_10568),
    .Y(n_10569));
 OAI21xp5_ASAP7_75t_SL g19347 (.A1(n_7721),
    .A2(n_3461),
    .B(n_10563),
    .Y(n_10568));
 NAND2xp5_ASAP7_75t_SL g19360 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_296),
    .B(n_17063),
    .Y(n_10585));
 NOR2xp33_ASAP7_75t_SL g19366 (.A(n_9259),
    .B(n_8016),
    .Y(n_10588));
 AOI21x1_ASAP7_75t_SL g19368 (.A1(n_10591),
    .A2(n_10592),
    .B(n_10594),
    .Y(n_10595));
 OR2x2_ASAP7_75t_SL g19369 (.A(n_21656),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_301),
    .Y(n_10591));
 NAND2xp5_ASAP7_75t_SL g19370 (.A(n_10593),
    .B(n_2163),
    .Y(n_10594));
 INVxp67_ASAP7_75t_SL g19371 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_213),
    .Y(n_10593));
 MAJIxp5_ASAP7_75t_SL g19384 (.A(n_4856),
    .B(n_8943),
    .C(n_21941),
    .Y(n_10608));
 MAJIxp5_ASAP7_75t_SL g19386 (.A(n_26242),
    .B(n_10611),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_30),
    .Y(n_10612));
 INVxp67_ASAP7_75t_SL g19387 (.A(n_10608),
    .Y(n_10611));
 INVx1_ASAP7_75t_SL g19391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_51),
    .Y(n_10613));
 XOR2xp5_ASAP7_75t_SL g19395 (.A(n_19053),
    .B(n_10622),
    .Y(n_10623));
 XNOR2xp5_ASAP7_75t_SL g19397 (.A(n_10621),
    .B(n_14653),
    .Y(n_10622));
 INVxp67_ASAP7_75t_SL g19398 (.A(n_9373),
    .Y(n_10621));
 AND2x2_ASAP7_75t_SL g194 (.A(n_22799),
    .B(n_22800),
    .Y(n_22808));
 NAND2xp5_ASAP7_75t_SL g19403 (.A(n_21247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_375),
    .Y(n_10628));
 XOR2xp5_ASAP7_75t_SL g19405 (.A(n_9441),
    .B(n_15551),
    .Y(n_10629));
 OR2x2_ASAP7_75t_SL g19411 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_100),
    .Y(n_10635));
 OAI22xp5_ASAP7_75t_SL g19415 (.A1(n_10640),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_30),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_158),
    .B2(n_10641),
    .Y(n_10642));
 MAJIxp5_ASAP7_75t_SL g19416 (.A(n_13844),
    .B(n_13845),
    .C(n_13843),
    .Y(n_10640));
 MAJIxp5_ASAP7_75t_SL g19419 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_103),
    .B(n_10645),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_78),
    .Y(n_10646));
 NAND2xp5_ASAP7_75t_SL g19420 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .Y(n_10645));
 XNOR2x1_ASAP7_75t_SL g19421 (.B(n_10647),
    .Y(n_10648),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_123));
 XNOR2xp5_ASAP7_75t_SL g19423 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_210),
    .B(n_21287),
    .Y(n_10650));
 NAND2xp33_ASAP7_75t_SL g19430 (.A(n_21849),
    .B(n_21848),
    .Y(n_10657));
 MAJIxp5_ASAP7_75t_SL g19439 (.A(n_25980),
    .B(n_19572),
    .C(n_10665),
    .Y(n_10666));
 INVxp67_ASAP7_75t_SL g19440 (.A(n_11070),
    .Y(n_10665));
 NAND2xp5_ASAP7_75t_SL g19451 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_11),
    .Y(n_10676));
 OR2x2_ASAP7_75t_SL g19452 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_11),
    .Y(n_10677));
 MAJx2_ASAP7_75t_SL g19458 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_12),
    .B(n_10684),
    .C(n_5660),
    .Y(n_10685));
 INVxp67_ASAP7_75t_SL g19459 (.A(n_19898),
    .Y(n_10684));
 MAJIxp5_ASAP7_75t_SL g19461 (.A(n_22604),
    .B(n_8107),
    .C(n_8109),
    .Y(n_10686));
 MAJIxp5_ASAP7_75t_SL g19464 (.A(n_22724),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(n_10693));
 XOR2xp5_ASAP7_75t_SL g19468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_238),
    .B(n_22724),
    .Y(n_10696));
 NAND2xp5_ASAP7_75t_SL g19471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_207),
    .B(n_8657),
    .Y(n_10697));
 NAND2xp5_ASAP7_75t_SL g19483 (.A(n_23776),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_296),
    .Y(n_10711));
 INVx1_ASAP7_75t_SL g19490 (.A(n_10718),
    .Y(n_10719));
 MAJx2_ASAP7_75t_SL g19491 (.A(n_7497),
    .B(n_7496),
    .C(n_7494),
    .Y(n_10718));
 INVxp67_ASAP7_75t_SL g19493 (.A(n_22151),
    .Y(n_10723));
 NAND2xp5_ASAP7_75t_SL g19495 (.A(n_21789),
    .B(n_10720),
    .Y(n_10721));
 INVxp67_ASAP7_75t_SL g19496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_213),
    .Y(n_10720));
 NOR2xp33_ASAP7_75t_SL g19499 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_211),
    .B(n_10721),
    .Y(n_10725));
 HB1xp67_ASAP7_75t_SL g195 (.A(n_11829),
    .Y(n_6099));
 NOR2xp33_ASAP7_75t_SL g19501 (.A(n_10728),
    .B(n_10730),
    .Y(n_10731));
 INVx1_ASAP7_75t_SL g19502 (.A(n_18703),
    .Y(n_10728));
 XNOR2xp5_ASAP7_75t_SL g19503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_126),
    .Y(n_10730));
 INVx1_ASAP7_75t_SL g19504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_108));
 NAND2xp5_ASAP7_75t_SL g19505 (.A(n_10728),
    .B(n_10730),
    .Y(n_10732));
 OAI21xp5_ASAP7_75t_SL g19506 (.A1(n_18703),
    .A2(n_10730),
    .B(n_10738),
    .Y(n_10739));
 AOI22xp5_ASAP7_75t_SL g19507 (.A1(n_10734),
    .A2(n_18703),
    .B1(n_10737),
    .B2(n_18703),
    .Y(n_10738));
 NOR2xp33_ASAP7_75t_SL g19508 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_126),
    .Y(n_10734));
 NOR2xp33_ASAP7_75t_SL g19510 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_107),
    .B(n_10736),
    .Y(n_10737));
 INVxp67_ASAP7_75t_SL g19511 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_126),
    .Y(n_10736));
 NAND2xp5_ASAP7_75t_SL g19512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_252),
    .B(n_10740),
    .Y(n_10741));
 XNOR2x1_ASAP7_75t_SL g19513 (.B(n_23375),
    .Y(n_10740),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_236));
 INVxp67_ASAP7_75t_SRAM g19515 (.A(n_10740),
    .Y(n_10742));
 NOR2x1_ASAP7_75t_SL g19516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_252),
    .B(n_10740),
    .Y(n_10744));
 XNOR2xp5_ASAP7_75t_SL g19523 (.A(n_10753),
    .B(n_19323),
    .Y(n_10754));
 XNOR2xp5_ASAP7_75t_SL g19524 (.A(n_10752),
    .B(n_19326),
    .Y(n_10753));
 INVx1_ASAP7_75t_SL g19525 (.A(n_19324),
    .Y(n_10752));
 OAI21x1_ASAP7_75t_SL g19527 (.A1(n_11835),
    .A2(n_10755),
    .B(n_10756),
    .Y(n_10757));
 AND2x2_ASAP7_75t_SL g19528 (.A(n_12111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109),
    .Y(n_10755));
 OR2x2_ASAP7_75t_SL g19529 (.A(n_12111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109),
    .Y(n_10756));
 OAI22xp5_ASAP7_75t_SL g19530 (.A1(n_18863),
    .A2(n_10757),
    .B1(n_10759),
    .B2(n_6463),
    .Y(n_10760));
 NOR2xp67_ASAP7_75t_SL g19533 (.A(n_18769),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_314),
    .Y(n_10762));
 INVx1_ASAP7_75t_SL g19539 (.A(n_8322),
    .Y(n_10765));
 INVx2_ASAP7_75t_SL g19543 (.A(n_20311),
    .Y(n_10771));
 MAJIxp5_ASAP7_75t_SL g19544 (.A(n_19905),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_216),
    .C(n_10773),
    .Y(n_10774));
 INVxp67_ASAP7_75t_SL g19545 (.A(n_20311),
    .Y(n_10773));
 XNOR2x1_ASAP7_75t_SL g19546 (.B(n_10776),
    .Y(n_10777),
    .A(n_10775));
 AOI22xp5_ASAP7_75t_SL g19547 (.A1(n_15240),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_91),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_93),
    .Y(n_10775));
 INVxp67_ASAP7_75t_SL g19548 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_126),
    .Y(n_10776));
 NAND2x1_ASAP7_75t_L g19550 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(n_10778));
 MAJIxp5_ASAP7_75t_SL g19559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_196),
    .B(n_10788),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_132),
    .Y(n_10789));
 NAND2xp5_ASAP7_75t_SL g19561 (.A(n_13951),
    .B(n_10790),
    .Y(n_10791));
 XNOR2xp5_ASAP7_75t_SL g19562 (.A(n_6474),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_246),
    .Y(n_10790));
 XNOR2xp5_ASAP7_75t_SL g19563 (.A(n_10792),
    .B(n_13951),
    .Y(n_10793));
 INVxp67_ASAP7_75t_SRAM g19564 (.A(n_10790),
    .Y(n_10792));
 OAI21xp5_ASAP7_75t_SL g19566 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_199),
    .A2(n_10795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_201),
    .Y(n_10796));
 NOR2xp67_ASAP7_75t_SL g19567 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_167),
    .Y(n_10795));
 XNOR2xp5_ASAP7_75t_SL g19569 (.A(n_10798),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_210),
    .Y(n_10799));
 INVxp67_ASAP7_75t_SL g19570 (.A(n_10795),
    .Y(n_10798));
 OAI21x1_ASAP7_75t_SL g19571 (.A1(n_10801),
    .A2(n_10802),
    .B(n_2168),
    .Y(n_10803));
 NOR2xp67_ASAP7_75t_SL g19572 (.A(n_18770),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_314),
    .Y(n_10801));
 AND2x2_ASAP7_75t_SL g19574 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_314),
    .B(n_18770),
    .Y(n_10802));
 NAND2xp5_ASAP7_75t_SL g19584 (.A(n_25132),
    .B(n_8369),
    .Y(n_10814));
 OAI21xp5_ASAP7_75t_SL g19586 (.A1(n_25131),
    .A2(n_14802),
    .B(n_8369),
    .Y(n_10816));
 XNOR2xp5_ASAP7_75t_SL g196 (.A(n_7615),
    .B(n_19910),
    .Y(n_19911));
 MAJx2_ASAP7_75t_SL g19607 (.A(n_6062),
    .B(n_10838),
    .C(n_10840),
    .Y(n_10841));
 HB1xp67_ASAP7_75t_SL g19608 (.A(n_6063),
    .Y(n_10838));
 HB1xp67_ASAP7_75t_SL g19609 (.A(n_10839),
    .Y(n_10840));
 XNOR2x1_ASAP7_75t_SL g19610 (.B(n_5991),
    .Y(n_10839),
    .A(n_5990));
 XNOR2xp5_ASAP7_75t_SL g19611 (.A(n_6063),
    .B(n_10839),
    .Y(n_10842));
 INVxp67_ASAP7_75t_SL g19617 (.A(n_9808),
    .Y(n_10847));
 INVx1_ASAP7_75t_SL g19618 (.A(n_2176),
    .Y(n_10848));
 XOR2xp5_ASAP7_75t_SL g19624 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_99),
    .B(n_12803),
    .Y(n_10856));
 NAND2xp5_ASAP7_75t_SL g19628 (.A(n_13389),
    .B(n_10859),
    .Y(n_10860));
 INVxp67_ASAP7_75t_SL g19629 (.A(n_13390),
    .Y(n_10859));
 MAJIxp5_ASAP7_75t_SL g19630 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_172),
    .B(n_10862),
    .C(n_10864),
    .Y(n_10865));
 INVxp67_ASAP7_75t_SL g19631 (.A(n_18775),
    .Y(n_10862));
 HB1xp67_ASAP7_75t_SL g19633 (.A(n_10863),
    .Y(n_10864));
 XNOR2x1_ASAP7_75t_SL g19634 (.B(n_4969),
    .Y(n_10863),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_27));
 XNOR2x1_ASAP7_75t_SL g19635 (.B(n_10863),
    .Y(n_10866),
    .A(n_18775));
 NAND2x1_ASAP7_75t_SL g19648 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(n_2927),
    .Y(n_10878));
 MAJIxp5_ASAP7_75t_SL g19651 (.A(n_18778),
    .B(n_10878),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_20),
    .Y(n_10882));
 XNOR2xp5_ASAP7_75t_SL g19652 (.A(n_10883),
    .B(n_10885),
    .Y(n_10886));
 INVx1_ASAP7_75t_SL g19653 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_153),
    .Y(n_10883));
 XNOR2xp5_ASAP7_75t_SL g19654 (.A(n_9514),
    .B(n_9516),
    .Y(n_10885));
 MAJIxp5_ASAP7_75t_SL g19656 (.A(n_6916),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_153),
    .C(n_10887),
    .Y(n_10888));
 HB1xp67_ASAP7_75t_SL g19657 (.A(n_10885),
    .Y(n_10887));
 OAI22xp5_ASAP7_75t_SL g19660 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_69),
    .A2(n_13725),
    .B1(n_4038),
    .B2(n_10891),
    .Y(n_10892));
 INVx1_ASAP7_75t_SL g19661 (.A(n_13725),
    .Y(n_10891));
 NAND2xp5_ASAP7_75t_SL g19664 (.A(n_24102),
    .B(n_10894),
    .Y(n_10895));
 INVx1_ASAP7_75t_SL g19665 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_225),
    .Y(n_10894));
 AOI21x1_ASAP7_75t_SL g19670 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_250),
    .A2(n_19543),
    .B(n_10901),
    .Y(n_10902));
 NOR2xp67_ASAP7_75t_SL g19671 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_239),
    .Y(n_10901));
 NAND2xp5_ASAP7_75t_SL g19672 (.A(n_10903),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_250),
    .Y(n_10904));
 INVxp67_ASAP7_75t_SRAM g19673 (.A(n_10901),
    .Y(n_10903));
 NAND2xp5_ASAP7_75t_SL g19676 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .Y(n_10905));
 MAJIxp5_ASAP7_75t_SL g19677 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_74),
    .B(n_10905),
    .C(n_22875),
    .Y(n_10908));
 XOR2xp5_ASAP7_75t_SL g19681 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_465),
    .B(n_22439),
    .Y(n_10912));
 MAJIxp5_ASAP7_75t_SL g19682 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_32),
    .B(n_13178),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_90),
    .Y(n_10915));
 NAND2x1_ASAP7_75t_SL g19684 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(n_14674),
    .Y(n_10913));
 OAI22xp5_ASAP7_75t_SL g19685 (.A1(n_10913),
    .A2(n_13779),
    .B1(n_13178),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_32),
    .Y(n_10916));
 MAJIxp5_ASAP7_75t_SL g19686 (.A(n_10917),
    .B(n_10918),
    .C(n_12114),
    .Y(n_10922));
 INVx1_ASAP7_75t_SL g19687 (.A(n_6421),
    .Y(n_10917));
 INVx1_ASAP7_75t_SL g19688 (.A(n_6420),
    .Y(n_10918));
 INVx1_ASAP7_75t_SL g197 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_108),
    .Y(n_6094));
 XOR2x2_ASAP7_75t_SL g19703 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_22),
    .B(n_12658),
    .Y(n_10933));
 AOI22xp5_ASAP7_75t_SL g19719 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_47),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_67),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_48),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_66),
    .Y(n_10947));
 NOR2xp33_ASAP7_75t_SL g19721 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_269),
    .B(n_10953),
    .Y(n_10954));
 MAJIxp5_ASAP7_75t_SL g19722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_238),
    .B(n_13449),
    .C(n_18737),
    .Y(n_10953));
 OAI21xp5_ASAP7_75t_SL g19727 (.A1(n_19857),
    .A2(n_19860),
    .B(n_10963),
    .Y(n_10964));
 OAI21xp5_ASAP7_75t_SL g19734 (.A1(n_19858),
    .A2(n_19856),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_142),
    .Y(n_10963));
 XNOR2x1_ASAP7_75t_SL g19737 (.B(n_10971),
    .Y(n_10972),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_27));
 OAI22xp5_ASAP7_75t_SL g19738 (.A1(n_10968),
    .A2(n_8781),
    .B1(n_10969),
    .B2(n_10970),
    .Y(n_10971));
 NAND2xp5_ASAP7_75t_R g19739 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .Y(n_10968));
 INVx1_ASAP7_75t_SL g19740 (.A(n_10968),
    .Y(n_10969));
 INVx1_ASAP7_75t_SL g19741 (.A(n_8781),
    .Y(n_10970));
 MAJIxp5_ASAP7_75t_SL g19742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_27),
    .B(n_10969),
    .C(n_8781),
    .Y(n_10973));
 MAJIxp5_ASAP7_75t_SL g19750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_19),
    .C(n_10981),
    .Y(n_10982));
 NAND2xp5_ASAP7_75t_SL g19751 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .Y(n_10981));
 XNOR2xp5_ASAP7_75t_SL g19752 (.A(n_10981),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_19),
    .Y(n_10983));
 XOR2xp5_ASAP7_75t_SL g19759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_187),
    .B(n_10995),
    .Y(n_7620));
 XNOR2xp5_ASAP7_75t_SL g19760 (.A(n_10990),
    .B(n_10994),
    .Y(n_10995));
 INVx1_ASAP7_75t_SL g19761 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_135),
    .Y(n_10990));
 AOI22xp5_ASAP7_75t_SL g19762 (.A1(n_10992),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_150),
    .B1(n_10993),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78),
    .Y(n_10994));
 INVx1_ASAP7_75t_L g19763 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78),
    .Y(n_10992));
 INVx1_ASAP7_75t_SL g19765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_150),
    .Y(n_10993));
 MAJIxp5_ASAP7_75t_SL g19766 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_187),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_150),
    .C(n_10998),
    .Y(n_10999));
 OAI22xp5_ASAP7_75t_SL g19768 (.A1(n_10992),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_135),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78),
    .B2(n_10990),
    .Y(n_10998));
 NAND2xp5_ASAP7_75t_SL g19771 (.A(n_11871),
    .B(n_9498),
    .Y(n_11000));
 MAJx2_ASAP7_75t_SL g19789 (.A(n_19398),
    .B(n_19400),
    .C(n_21469),
    .Y(n_11021));
 XNOR2xp5_ASAP7_75t_SL g19792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_647),
    .B(n_11022),
    .Y(n_11023));
 AND2x2_ASAP7_75t_SL g19793 (.A(n_2179),
    .B(n_13524),
    .Y(n_11022));
 NAND2xp5_ASAP7_75t_SL g19795 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_647),
    .B(n_11022),
    .Y(n_11026));
 OAI21xp5_ASAP7_75t_SL g19796 (.A1(n_11028),
    .A2(n_11029),
    .B(n_11031),
    .Y(n_11032));
 NAND2xp5_ASAP7_75t_SL g19797 (.A(n_11027),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_308),
    .Y(n_11028));
 INVxp67_ASAP7_75t_SL g19798 (.A(n_14382),
    .Y(n_11027));
 INVxp67_ASAP7_75t_SL g19799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_310),
    .Y(n_11029));
 NOR2xp33_ASAP7_75t_SL g198 (.A(n_20036),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_301),
    .Y(n_20037));
 AOI21xp33_ASAP7_75t_SL g19800 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_311),
    .A2(n_11027),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_274),
    .Y(n_11031));
 NAND3xp33_ASAP7_75t_SL g19805 (.A(n_11920),
    .B(n_20099),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278),
    .Y(n_11039));
 AOI21x1_ASAP7_75t_SL g19808 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_303),
    .A2(n_11040),
    .B(n_11042),
    .Y(n_11043));
 HB1xp67_ASAP7_75t_SL g19809 (.A(n_11920),
    .Y(n_11040));
 HB1xp67_ASAP7_75t_SL g19810 (.A(n_11041),
    .Y(n_11042));
 OAI21xp5_ASAP7_75t_SL g19811 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_285),
    .A2(n_11919),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_282),
    .Y(n_11041));
 AOI21xp5_ASAP7_75t_SL g19812 (.A1(n_11044),
    .A2(n_10685),
    .B(n_11919),
    .Y(n_11045));
 HB1xp67_ASAP7_75t_SL g19813 (.A(n_11918),
    .Y(n_11044));
 NAND2xp5_ASAP7_75t_SL g19820 (.A(n_11054),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_155),
    .Y(n_11056));
 XNOR2xp5_ASAP7_75t_SL g19821 (.A(n_18778),
    .B(n_18960),
    .Y(n_11054));
 NOR2xp33_ASAP7_75t_SL g19825 (.A(n_11054),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_155),
    .Y(n_11058));
 AND2x2_ASAP7_75t_SL g19830 (.A(n_7011),
    .B(n_11063),
    .Y(n_11064));
 XNOR2xp5_ASAP7_75t_SL g19831 (.A(n_11062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_238),
    .Y(n_11063));
 XNOR2xp5_ASAP7_75t_SL g19832 (.A(n_8092),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_26),
    .Y(n_11062));
 NOR2xp67_ASAP7_75t_SL g19833 (.A(n_7011),
    .B(n_11063),
    .Y(n_11065));
 XNOR2x1_ASAP7_75t_SL g19834 (.B(n_11069),
    .Y(n_11070),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_192));
 XNOR2x1_ASAP7_75t_SL g19835 (.B(n_20093),
    .Y(n_11069),
    .A(n_11066));
 INVx1_ASAP7_75t_SL g19838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_108),
    .Y(n_11067));
 MAJIxp5_ASAP7_75t_SL g19839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_192),
    .B(n_11071),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_28),
    .Y(n_11072));
 OAI21xp5_ASAP7_75t_SL g19846 (.A1(n_9036),
    .A2(n_5617),
    .B(n_6204),
    .Y(n_11077));
 OAI22xp5_ASAP7_75t_SL g19852 (.A1(n_11084),
    .A2(n_11085),
    .B1(n_15464),
    .B2(n_15223),
    .Y(n_11088));
 NAND2xp5_ASAP7_75t_SL g19853 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .Y(n_11084));
 NAND2x1_ASAP7_75t_SL g19854 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(n_14523),
    .Y(n_11085));
 MAJIxp5_ASAP7_75t_SL g19857 (.A(n_7885),
    .B(n_15223),
    .C(n_15464),
    .Y(n_11090));
 MAJIxp5_ASAP7_75t_SL g19858 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_77),
    .C(n_11094),
    .Y(n_11095));
 HB1xp67_ASAP7_75t_SL g19859 (.A(n_11093),
    .Y(n_11094));
 MAJIxp5_ASAP7_75t_SL g19860 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_99),
    .C(n_11092),
    .Y(n_11093));
 INVx1_ASAP7_75t_SL g19861 (.A(n_11091),
    .Y(n_11092));
 NAND2xp5_ASAP7_75t_SL g19862 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(n_12800),
    .Y(n_11091));
 OAI22xp5_ASAP7_75t_SL g19863 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_76),
    .A2(n_11093),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_77),
    .B2(n_11096),
    .Y(n_11097));
 INVx1_ASAP7_75t_SL g19864 (.A(n_11093),
    .Y(n_11096));
 OAI22xp5_ASAP7_75t_SL g19865 (.A1(n_11091),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_78),
    .B1(n_11092),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_79),
    .Y(n_11098));
 NOR2xp33_ASAP7_75t_SL g19872 (.A(n_11830),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .Y(n_11105));
 AND2x2_ASAP7_75t_SL g19879 (.A(n_13235),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_79),
    .Y(n_11112));
 XNOR2x1_ASAP7_75t_SL g19881 (.B(n_11112),
    .Y(n_11116),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_6));
 XOR2x2_ASAP7_75t_SL g19882 (.A(n_22261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_12),
    .Y(n_11120));
 AND2x2_ASAP7_75t_SL g19887 (.A(n_22078),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_243),
    .Y(n_11124));
 NAND2xp5_ASAP7_75t_SL g19890 (.A(n_11125),
    .B(n_11389),
    .Y(n_11126));
 INVxp67_ASAP7_75t_SL g19891 (.A(n_22078),
    .Y(n_11125));
 MAJIxp5_ASAP7_75t_SL g19892 (.A(n_22077),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_216),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_207),
    .Y(n_11127));
 XNOR2xp5_ASAP7_75t_SL g19893 (.A(n_11129),
    .B(n_11132),
    .Y(n_11133));
 INVx1_ASAP7_75t_SL g19894 (.A(n_11128),
    .Y(n_11129));
 XNOR2xp5_ASAP7_75t_SL g19895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_118),
    .B(n_5896),
    .Y(n_11128));
 AOI22xp5_ASAP7_75t_SL g19896 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_195),
    .A2(n_11130),
    .B1(n_11131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_190),
    .Y(n_11132));
 INVx1_ASAP7_75t_SL g19897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_190),
    .Y(n_11130));
 INVx1_ASAP7_75t_SL g19898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_195),
    .Y(n_11131));
 MAJIxp5_ASAP7_75t_SL g19899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_224),
    .B(n_11134),
    .C(n_11136),
    .Y(n_11137));
 XOR2xp5_ASAP7_75t_SL g199 (.A(n_20121),
    .B(n_23451),
    .Y(n_11517));
 HB1xp67_ASAP7_75t_SL g19900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_190),
    .Y(n_11134));
 XNOR2xp5_ASAP7_75t_SL g19901 (.A(n_11129),
    .B(n_11135),
    .Y(n_11136));
 HB1xp67_ASAP7_75t_SL g19902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_195),
    .Y(n_11135));
 MAJIxp5_ASAP7_75t_SL g19903 (.A(n_11128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_165),
    .Y(n_11138));
 HB1xp67_ASAP7_75t_SL g19909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_21),
    .Y(n_11142));
 XOR2xp5_ASAP7_75t_SL g19910 (.A(n_23682),
    .B(n_23684),
    .Y(n_11145));
 OAI21xp5_ASAP7_75t_SL g19917 (.A1(n_8902),
    .A2(n_11151),
    .B(n_6788),
    .Y(n_11152));
 AOI21x1_ASAP7_75t_SL g19918 (.A1(n_8696),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_297),
    .Y(n_11151));
 OAI21xp33_ASAP7_75t_SL g19928 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_496),
    .A2(n_5331),
    .B(n_11164),
    .Y(n_11165));
 AOI21xp5_ASAP7_75t_SL g19929 (.A1(n_5334),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_496),
    .B(n_18779),
    .Y(n_11164));
 XNOR2x2_ASAP7_75t_SL g19931 (.A(n_11168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_13),
    .Y(n_11169));
 MAJIxp5_ASAP7_75t_SL g19932 (.A(n_15999),
    .B(n_24107),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_717),
    .Y(n_11168));
 MAJIxp5_ASAP7_75t_SL g19939 (.A(n_22230),
    .B(n_10249),
    .C(n_6304),
    .Y(n_11175));
 A2O1A1Ixp33_ASAP7_75t_SL g19940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_31),
    .B(n_22229),
    .C(n_11176),
    .Y(n_11177));
 OR2x2_ASAP7_75t_SL g19941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_31),
    .Y(n_11176));
 OAI21xp5_ASAP7_75t_SL g19943 (.A1(n_9455),
    .A2(n_6102),
    .B(n_7705),
    .Y(n_11178));
 OAI22xp33_ASAP7_75t_SL g19952 (.A1(n_8531),
    .A2(n_18907),
    .B1(n_8532),
    .B2(n_11192),
    .Y(n_11193));
 NAND2xp5_ASAP7_75t_SL g19954 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .Y(n_11189));
 INVxp67_ASAP7_75t_SL g19956 (.A(n_18907),
    .Y(n_11192));
 MAJx2_ASAP7_75t_SL g19957 (.A(n_8530),
    .B(n_18907),
    .C(n_8532),
    .Y(n_11194));
 AND2x2_ASAP7_75t_SL g19958 (.A(n_11189),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_46),
    .Y(n_11195));
 MAJIxp5_ASAP7_75t_SL g19959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_42),
    .C(n_11198),
    .Y(n_3461));
 INVx1_ASAP7_75t_SL g19960 (.A(n_11197),
    .Y(n_11198));
 OR2x2_ASAP7_75t_SL g19961 (.A(n_11196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_92),
    .Y(n_11197));
 NAND2xp5_ASAP7_75t_SL g19962 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .Y(n_11196));
 XNOR2xp5_ASAP7_75t_SL g19963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_117),
    .B(n_11198),
    .Y(n_11200));
 NAND2xp5_ASAP7_75t_SL g19965 (.A(n_11196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_92),
    .Y(n_11201));
 XNOR2xp5_ASAP7_75t_SL g19968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_27),
    .B(n_8032),
    .Y(n_11204));
 MAJIxp5_ASAP7_75t_SL g19971 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_172),
    .B(n_11208),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_136),
    .Y(n_11209));
 INVxp67_ASAP7_75t_SL g19972 (.A(n_11204),
    .Y(n_11208));
 AOI21xp5_ASAP7_75t_SL g19973 (.A1(n_11212),
    .A2(n_9992),
    .B(n_9991),
    .Y(n_11213));
 NOR2xp33_ASAP7_75t_SL g19974 (.A(n_11867),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_260),
    .Y(n_11212));
 NAND2xp33_ASAP7_75t_R g19977 (.A(n_11868),
    .B(n_11215),
    .Y(n_11216));
 OR2x2_ASAP7_75t_SL g19979 (.A(n_11867),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_260),
    .Y(n_11215));
 XNOR2x1_ASAP7_75t_SL g19982 (.B(n_11219),
    .Y(n_11220),
    .A(n_11218));
 XNOR2x1_ASAP7_75t_SL g19983 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_224),
    .Y(n_11218),
    .A(n_19200));
 INVxp67_ASAP7_75t_SL g19984 (.A(n_14868),
    .Y(n_11219));
 OAI22xp5_ASAP7_75t_SL g19995 (.A1(n_11235),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_293),
    .B1(n_13934),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_294),
    .Y(n_11236));
 INVx2_ASAP7_75t_SL g19996 (.A(n_13934),
    .Y(n_11235));
 OR2x2_ASAP7_75t_SL g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_160),
    .Y(n_18695));
 NAND2x1p5_ASAP7_75t_SL g20 (.A(n_9570),
    .B(n_9571),
    .Y(n_3206));
 MAJx2_ASAP7_75t_SL g200 (.A(n_22419),
    .B(n_11519),
    .C(n_11520),
    .Y(n_11521));
 INVxp67_ASAP7_75t_SL g20002 (.A(n_13930),
    .Y(n_11238));
 OAI21xp5_ASAP7_75t_SL g20004 (.A1(n_13930),
    .A2(n_13932),
    .B(n_11151),
    .Y(n_11241));
 OAI21xp33_ASAP7_75t_SL g20005 (.A1(n_8691),
    .A2(n_13930),
    .B(n_8697),
    .Y(n_11242));
 MAJIxp5_ASAP7_75t_SL g20008 (.A(n_9659),
    .B(n_9658),
    .C(n_9657),
    .Y(n_11243));
 MAJIxp5_ASAP7_75t_SL g20009 (.A(n_17754),
    .B(n_11248),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_72),
    .Y(n_11249));
 MAJIxp5_ASAP7_75t_SL g20024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_251),
    .B(n_18780),
    .C(n_11266),
    .Y(n_11267));
 XNOR2xp5_ASAP7_75t_SL g20026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_212),
    .Y(n_11266));
 XNOR2xp5_ASAP7_75t_SL g20027 (.A(n_18780),
    .B(n_11266),
    .Y(n_11268));
 MAJIxp5_ASAP7_75t_SL g20029 (.A(n_11269),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_71),
    .C(n_21184),
    .Y(n_11270));
 NAND2xp5_ASAP7_75t_SL g20030 (.A(n_6965),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .Y(n_11269));
 XNOR2xp5_ASAP7_75t_SL g20036 (.A(n_11269),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_2),
    .Y(n_11277));
 XNOR2x2_ASAP7_75t_SL g20046 (.A(n_11725),
    .B(n_26150),
    .Y(n_11295));
 NAND2x1_ASAP7_75t_SL g20049 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_684),
    .Y(n_11289));
 NOR3xp33_ASAP7_75t_SL g20056 (.A(n_11299),
    .B(n_15088),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_308),
    .Y(n_11300));
 INVx1_ASAP7_75t_SL g20057 (.A(n_11298),
    .Y(n_11299));
 NAND2xp5_ASAP7_75t_SL g20058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_288),
    .B(n_11419),
    .Y(n_11298));
 HB1xp67_ASAP7_75t_SL g20060 (.A(n_11298),
    .Y(n_11302));
 INVxp67_ASAP7_75t_SL g20062 (.A(n_11302),
    .Y(n_11304));
 NAND2xp5_ASAP7_75t_SL g20064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_208),
    .B(n_11308),
    .Y(n_11309));
 XNOR2xp5_ASAP7_75t_SL g20065 (.A(n_7963),
    .B(n_11307),
    .Y(n_11308));
 AOI22xp5_ASAP7_75t_SL g20066 (.A1(n_24754),
    .A2(n_7965),
    .B1(n_7964),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154),
    .Y(n_11307));
 NOR2xp67_ASAP7_75t_SL g20067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_208),
    .B(n_11308),
    .Y(n_11310));
 NAND2xp5_ASAP7_75t_SL g20068 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .B(n_11316),
    .Y(n_11317));
 NOR2xp33_ASAP7_75t_SL g20069 (.A(n_5996),
    .B(n_11315),
    .Y(n_11316));
 INVxp67_ASAP7_75t_SL g20071 (.A(n_23738),
    .Y(n_11315));
 AOI21xp5_ASAP7_75t_L g20075 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .A2(n_23738),
    .B(n_5996),
    .Y(n_11318));
 OAI21xp5_ASAP7_75t_SL g20076 (.A1(n_21266),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_446),
    .B(n_23738),
    .Y(n_11320));
 MAJIxp5_ASAP7_75t_SL g20078 (.A(n_23018),
    .B(n_8027),
    .C(n_11323),
    .Y(n_11324));
 HB1xp67_ASAP7_75t_SL g20079 (.A(n_11322),
    .Y(n_11323));
 MAJIxp5_ASAP7_75t_SL g20080 (.A(n_11321),
    .B(n_8864),
    .C(n_8866),
    .Y(n_11322));
 XNOR2xp5_ASAP7_75t_SL g20081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_89),
    .B(n_10629),
    .Y(n_11321));
 XOR2xp5_ASAP7_75t_SL g20082 (.A(n_8862),
    .B(n_11322),
    .Y(n_11325));
 XOR2xp5_ASAP7_75t_SL g20083 (.A(n_11326),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_186),
    .Y(n_11327));
 INVx1_ASAP7_75t_SL g20084 (.A(n_11321),
    .Y(n_11326));
 AOI22xp5_ASAP7_75t_SL g20087 (.A1(n_14675),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_83),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_84),
    .B2(n_13681),
    .Y(n_11328));
 MAJIxp5_ASAP7_75t_SL g20089 (.A(n_11333),
    .B(n_2437),
    .C(n_8882),
    .Y(n_11334));
 XNOR2x1_ASAP7_75t_SL g20090 (.B(n_11332),
    .Y(n_11333),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41));
 OAI21x1_ASAP7_75t_SL g20091 (.A1(n_2580),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .B(n_8888),
    .Y(n_11332));
 XOR2xp5_ASAP7_75t_SL g20095 (.A(n_11340),
    .B(n_23122),
    .Y(n_11341));
 NOR2xp33_ASAP7_75t_R g20096 (.A(n_5630),
    .B(n_11339),
    .Y(n_11340));
 INVxp33_ASAP7_75t_SL g20097 (.A(n_11338),
    .Y(n_11339));
 NAND2xp5_ASAP7_75t_SL g20098 (.A(n_26222),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_271),
    .Y(n_11338));
 INVxp67_ASAP7_75t_SL g201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_213),
    .Y(n_20035));
 NAND2xp5_ASAP7_75t_SL g20100 (.A(n_11338),
    .B(n_7947),
    .Y(n_11343));
 OAI22xp5_ASAP7_75t_SL g20103 (.A1(n_11346),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_158),
    .B1(n_9138),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30),
    .Y(n_11348));
 AND2x2_ASAP7_75t_SL g20104 (.A(n_11346),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30),
    .Y(n_11350));
 MAJx2_ASAP7_75t_SL g20113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_68),
    .C(n_22876),
    .Y(n_11361));
 OAI22xp5_ASAP7_75t_SL g20121 (.A1(n_10174),
    .A2(n_10169),
    .B1(n_10173),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .Y(n_11374));
 XNOR2x1_ASAP7_75t_SL g20127 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_723),
    .Y(n_11377),
    .A(n_11376));
 XNOR2x1_ASAP7_75t_SL g20128 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_563),
    .Y(n_11376),
    .A(n_11375));
 NAND2xp5_ASAP7_75t_SL g20129 (.A(n_2158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_786),
    .Y(n_11375));
 INVxp67_ASAP7_75t_SL g20132 (.A(n_11375),
    .Y(n_11379));
 OAI21xp5_ASAP7_75t_SL g20133 (.A1(n_11382),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .B(n_11383),
    .Y(n_11384));
 NOR2xp33_ASAP7_75t_SL g20134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_363),
    .B(n_11381),
    .Y(n_11382));
 XNOR2x1_ASAP7_75t_SL g20135 (.B(n_19050),
    .Y(n_11381),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_34));
 NAND2xp5_ASAP7_75t_SL g20136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_363),
    .B(n_11381),
    .Y(n_11383));
 OAI21xp33_ASAP7_75t_SRAM g20137 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_363),
    .A2(n_11381),
    .B(n_11383),
    .Y(n_11385));
 XNOR2xp5_ASAP7_75t_SL g20138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_10),
    .B(n_11387),
    .Y(n_11388));
 XNOR2xp5_ASAP7_75t_SL g20139 (.A(n_5553),
    .B(n_11386),
    .Y(n_11387));
 AOI22xp5_ASAP7_75t_SL g20140 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_126),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_145),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_127),
    .B2(n_15210),
    .Y(n_11386));
 MAJIxp5_ASAP7_75t_SL g20141 (.A(n_11387),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_7),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_165),
    .Y(n_11389));
 NAND2x1_ASAP7_75t_SL g20156 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B(n_19391),
    .Y(n_11401));
 XNOR2xp5_ASAP7_75t_SL g20157 (.A(n_11403),
    .B(n_11404),
    .Y(n_11405));
 INVx2_ASAP7_75t_SL g20158 (.A(n_13782),
    .Y(n_11403));
 NAND2xp5_ASAP7_75t_SL g20160 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_2985),
    .Y(n_11404));
 MAJIxp5_ASAP7_75t_SL g20161 (.A(n_11409),
    .B(n_11401),
    .C(n_11403),
    .Y(n_11411));
 INVxp67_ASAP7_75t_SL g20162 (.A(n_11404),
    .Y(n_11409));
 XNOR2xp5_ASAP7_75t_SL g20164 (.A(n_5129),
    .B(n_11417),
    .Y(n_11418));
 XNOR2x1_ASAP7_75t_SL g20165 (.B(n_11412),
    .Y(n_11417),
    .A(n_14244));
 MAJIxp5_ASAP7_75t_SL g20168 (.A(n_11417),
    .B(n_3243),
    .C(n_13188),
    .Y(n_11419));
 OAI21xp5_ASAP7_75t_SL g20169 (.A1(n_14243),
    .A2(n_11421),
    .B(n_14242),
    .Y(n_11423));
 INVx1_ASAP7_75t_SL g20171 (.A(n_11412),
    .Y(n_11421));
 AO21x1_ASAP7_75t_SL g20174 (.A1(n_11425),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_293),
    .B(n_11430),
    .Y(n_11431));
 AND2x2_ASAP7_75t_SL g20175 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254),
    .B(n_11424),
    .Y(n_11425));
 AND2x2_ASAP7_75t_SL g20176 (.A(n_2151),
    .B(n_5751),
    .Y(n_11424));
 OAI31xp33_ASAP7_75t_SL g20178 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_293),
    .A2(n_11427),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253),
    .B(n_11429),
    .Y(n_11430));
 NAND2xp5_ASAP7_75t_SL g20179 (.A(n_2151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_251),
    .Y(n_11427));
 AOI31xp33_ASAP7_75t_SL g20180 (.A1(n_11424),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254),
    .B(n_11428),
    .Y(n_11429));
 NOR2xp33_ASAP7_75t_SL g20181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254),
    .B(n_11427),
    .Y(n_11428));
 XNOR2xp5_ASAP7_75t_SL g20182 (.A(n_11431),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_14),
    .Y(n_11433));
 NAND2xp5_ASAP7_75t_SL g20188 (.A(n_2307),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .Y(n_11438));
 MAJIxp5_ASAP7_75t_SL g20192 (.A(n_11445),
    .B(n_19679),
    .C(n_19680),
    .Y(n_11446));
 INVx1_ASAP7_75t_SL g20193 (.A(n_11438),
    .Y(n_11445));
 XNOR2xp5_ASAP7_75t_SL g20194 (.A(n_18782),
    .B(n_11451),
    .Y(n_11452));
 XOR2xp5_ASAP7_75t_SL g20197 (.A(n_11449),
    .B(n_11450),
    .Y(n_11451));
 MAJIxp5_ASAP7_75t_SL g20198 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_753),
    .B(n_17732),
    .C(n_17735),
    .Y(n_11449));
 XOR2xp5_ASAP7_75t_SL g20199 (.A(n_8646),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_7),
    .Y(n_11450));
 XNOR2xp5_ASAP7_75t_SL g202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_230),
    .B(n_6365),
    .Y(n_6366));
 NAND2xp5_ASAP7_75t_SL g20200 (.A(n_11453),
    .B(n_6724),
    .Y(n_11454));
 INVx1_ASAP7_75t_SL g20201 (.A(n_11452),
    .Y(n_11453));
 MAJIxp5_ASAP7_75t_SL g20202 (.A(n_18782),
    .B(n_11449),
    .C(n_11455),
    .Y(n_11456));
 INVxp67_ASAP7_75t_SL g20203 (.A(n_11450),
    .Y(n_11455));
 MAJx2_ASAP7_75t_SL g20209 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_75),
    .B(n_7463),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_67),
    .Y(n_11458));
 INVx1_ASAP7_75t_SL g20210 (.A(n_18972),
    .Y(n_11462));
 INVx2_ASAP7_75t_SL g20214 (.A(n_11458),
    .Y(n_11463));
 MAJx2_ASAP7_75t_SL g20216 (.A(n_11463),
    .B(n_11462),
    .C(n_17976),
    .Y(n_11469));
 INVx2_ASAP7_75t_SL g20222 (.A(n_11501),
    .Y(n_11502));
 XNOR2x1_ASAP7_75t_SL g20223 (.B(n_14819),
    .Y(n_11501),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_115));
 MAJIxp5_ASAP7_75t_SL g20228 (.A(n_11502),
    .B(n_11509),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_147),
    .Y(n_11510));
 INVxp67_ASAP7_75t_SRAM g20235 (.A(n_20121),
    .Y(n_11519));
 INVxp67_ASAP7_75t_SL g20236 (.A(n_23451),
    .Y(n_11520));
 XNOR2x1_ASAP7_75t_SL g20241 (.B(n_11528),
    .Y(n_11529),
    .A(n_11525));
 XOR2xp5_ASAP7_75t_SL g20242 (.A(n_11526),
    .B(n_11527),
    .Y(n_11528));
 NAND2xp5_ASAP7_75t_SL g20243 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .Y(n_11526));
 AND2x2_ASAP7_75t_SL g20244 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .Y(n_11527));
 MAJx2_ASAP7_75t_SL g20246 (.A(n_8962),
    .B(n_11529),
    .C(n_13100),
    .Y(n_11533));
 MAJIxp5_ASAP7_75t_SL g20247 (.A(n_11525),
    .B(n_11527),
    .C(n_11526),
    .Y(n_11534));
 NOR2xp67_ASAP7_75t_SL g20248 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .B(n_11539),
    .Y(n_11540));
 XNOR2xp5_ASAP7_75t_SL g20249 (.A(n_11535),
    .B(n_11536),
    .Y(n_11537));
 MAJIxp5_ASAP7_75t_SL g20250 (.A(n_19012),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_211),
    .C(n_13406),
    .Y(n_11535));
 XOR2xp5_ASAP7_75t_SL g20251 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(n_21168),
    .Y(n_11536));
 XOR2xp5_ASAP7_75t_SL g20252 (.A(n_13617),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_276),
    .Y(n_11538));
 NAND2xp5_ASAP7_75t_SL g20253 (.A(n_11539),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .Y(n_11541));
 MAJx2_ASAP7_75t_SL g20254 (.A(n_11538),
    .B(n_11542),
    .C(n_11543),
    .Y(n_11544));
 INVxp67_ASAP7_75t_SL g20255 (.A(n_11535),
    .Y(n_11542));
 HB1xp67_ASAP7_75t_SL g20256 (.A(n_11536),
    .Y(n_11543));
 XNOR2x1_ASAP7_75t_SL g20257 (.B(n_22958),
    .Y(n_11550),
    .A(n_11547));
 XNOR2xp5_ASAP7_75t_SL g20258 (.A(n_11545),
    .B(n_11546),
    .Y(n_11547));
 MAJx2_ASAP7_75t_SL g20259 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_751),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_687),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_591),
    .Y(n_11545));
 XNOR2x1_ASAP7_75t_SL g20260 (.B(n_8235),
    .Y(n_11546),
    .A(n_8245));
 MAJIxp5_ASAP7_75t_SL g20276 (.A(n_11610),
    .B(n_20519),
    .C(n_7727),
    .Y(n_11611));
 XNOR2x1_ASAP7_75t_SL g20287 (.B(n_20128),
    .Y(n_11612),
    .A(n_20520));
 XNOR2x2_ASAP7_75t_SL g20291 (.A(n_18124),
    .B(n_11621),
    .Y(n_11622));
 XNOR2x1_ASAP7_75t_SL g20295 (.B(n_11620),
    .Y(n_11621),
    .A(n_11618));
 AND2x2_ASAP7_75t_SL g20296 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_52),
    .Y(n_11618));
 XNOR2xp5_ASAP7_75t_SL g20297 (.A(n_18718),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_129),
    .Y(n_11620));
 MAJIxp5_ASAP7_75t_SL g20300 (.A(n_11625),
    .B(n_22074),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_147),
    .Y(n_11627));
 INVxp67_ASAP7_75t_SL g20301 (.A(n_11621),
    .Y(n_11625));
 MAJIxp5_ASAP7_75t_SL g20303 (.A(n_3366),
    .B(n_11618),
    .C(n_18718),
    .Y(n_3615));
 NOR2xp33_ASAP7_75t_SL g20363 (.A(n_18783),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_330),
    .Y(n_11722));
 AND2x2_ASAP7_75t_SL g20365 (.A(n_18783),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_330),
    .Y(n_11723));
 OAI21x1_ASAP7_75t_SL g20366 (.A1(n_11725),
    .A2(n_22169),
    .B(n_22170),
    .Y(n_11726));
 AND2x2_ASAP7_75t_SL g20367 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_748),
    .B(n_2151),
    .Y(n_11725));
 NAND2x1_ASAP7_75t_SL g20371 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .B(n_3868),
    .Y(n_11729));
 AOI21x1_ASAP7_75t_SL g20378 (.A1(n_9801),
    .A2(n_11300),
    .B(n_14427),
    .Y(n_11739));
 XNOR2x1_ASAP7_75t_SL g20380 (.B(n_11742),
    .Y(n_11743),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_148));
 OAI22xp5_ASAP7_75t_SL g20381 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_165),
    .A2(n_13056),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_166),
    .B2(n_14204),
    .Y(n_11742));
 OAI22xp5_ASAP7_75t_SL g20389 (.A1(n_11751),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_39),
    .B1(n_11752),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_38),
    .Y(n_11753));
 NAND2x1_ASAP7_75t_SL g20390 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(n_22156),
    .Y(n_11751));
 INVx2_ASAP7_75t_SL g20391 (.A(n_11751),
    .Y(n_11752));
 XNOR2x1_ASAP7_75t_SL g20397 (.B(n_11761),
    .Y(n_11762),
    .A(n_21230));
 XNOR2x2_ASAP7_75t_SL g20398 (.A(n_11760),
    .B(n_19177),
    .Y(n_11761));
 MAJx2_ASAP7_75t_SL g20399 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_166),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_148),
    .Y(n_11760));
 NAND2x1_ASAP7_75t_SL g204 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .B(n_4275),
    .Y(n_20696));
 XNOR2xp5_ASAP7_75t_SL g20402 (.A(n_10765),
    .B(n_17488),
    .Y(n_11763));
 OAI21xp5_ASAP7_75t_SL g20405 (.A1(n_11767),
    .A2(n_19515),
    .B(n_8368),
    .Y(n_11768));
 AOI21xp5_ASAP7_75t_SL g20406 (.A1(n_7342),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_290),
    .B(n_5487),
    .Y(n_11767));
 NAND2xp5_ASAP7_75t_SL g20408 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(n_11770),
    .Y(n_11771));
 AND2x2_ASAP7_75t_SL g20418 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_243),
    .B(n_23019),
    .Y(n_11781));
 OAI33xp33_ASAP7_75t_SL g20420 (.A1(n_11324),
    .A2(n_10558),
    .A3(n_11789),
    .B1(n_11324),
    .B2(n_11788),
    .B3(n_23450),
    .Y(n_11790));
 AOI22x1_ASAP7_75t_SL g20422 (.A1(n_22519),
    .A2(n_7255),
    .B1(n_14213),
    .B2(n_11787),
    .Y(n_11788));
 INVx1_ASAP7_75t_SL g20424 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_149),
    .Y(n_11783));
 XOR2xp5_ASAP7_75t_SL g20427 (.A(n_11800),
    .B(n_20372),
    .Y(n_11793));
 AND2x2_ASAP7_75t_SL g20436 (.A(n_2182),
    .B(n_13405),
    .Y(n_11800));
 NAND2xp5_ASAP7_75t_SL g20437 (.A(n_20988),
    .B(n_18764),
    .Y(n_11808));
 INVx1_ASAP7_75t_SL g20448 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_275),
    .Y(n_11812));
 MAJx2_ASAP7_75t_SL g20453 (.A(n_11818),
    .B(n_12747),
    .C(n_21925),
    .Y(n_11819));
 AND2x2_ASAP7_75t_SL g20454 (.A(n_2165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_674),
    .Y(n_11818));
 OAI22xp5_ASAP7_75t_SL g20456 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_3),
    .A2(n_11821),
    .B1(n_11822),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_140),
    .Y(n_11823));
 MAJIxp5_ASAP7_75t_SL g20457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_60),
    .B(n_23825),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_78),
    .Y(n_11821));
 INVx1_ASAP7_75t_SL g20458 (.A(n_11821),
    .Y(n_11822));
 XNOR2x1_ASAP7_75t_SL g20459 (.B(n_11828),
    .Y(n_11829),
    .A(n_9092));
 NAND2x1p5_ASAP7_75t_SL g20461 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .B(n_2825),
    .Y(n_11826));
 INVx2_ASAP7_75t_SL g20462 (.A(n_11826),
    .Y(n_11827));
 XNOR2xp5_ASAP7_75t_SL g20463 (.A(n_22893),
    .B(n_21673),
    .Y(n_11832));
 OAI22x1_ASAP7_75t_SL g20465 (.A1(n_6669),
    .A2(n_6082),
    .B1(n_18964),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_n_737),
    .Y(n_11830));
 XNOR2x1_ASAP7_75t_SL g20468 (.B(n_7558),
    .Y(n_11835),
    .A(n_26039));
 XOR2xp5_ASAP7_75t_SL g20475 (.A(n_11845),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_140),
    .Y(n_11846));
 NAND2xp5_ASAP7_75t_SL g20476 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(n_2293),
    .Y(n_11845));
 XNOR2xp5_ASAP7_75t_SL g20479 (.A(n_26200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_183),
    .Y(n_11852));
 OAI21x1_ASAP7_75t_SL g20483 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_287),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_289),
    .B(n_11856),
    .Y(n_11857));
 OA21x2_ASAP7_75t_SL g20484 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_280),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_283),
    .B(n_11855),
    .Y(n_11856));
 AOI21xp5_ASAP7_75t_SL g20485 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_276),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_259),
    .B(n_11854),
    .Y(n_11855));
 INVx1_ASAP7_75t_SL g20486 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_8),
    .Y(n_11854));
 NAND2xp5_ASAP7_75t_SL g20489 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_258),
    .B(n_9841),
    .Y(n_11858));
 NOR2xp67_ASAP7_75t_SL g20493 (.A(n_9536),
    .B(n_11865),
    .Y(n_3681));
 XNOR2xp5_ASAP7_75t_SL g20494 (.A(n_10483),
    .B(n_20110),
    .Y(n_11865));
 INVx1_ASAP7_75t_SL g20497 (.A(n_11868),
    .Y(n_11869));
 NAND2xp5_ASAP7_75t_SL g20498 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_260),
    .B(n_11867),
    .Y(n_11868));
 XNOR2x1_ASAP7_75t_SL g20499 (.B(n_11612),
    .Y(n_11867),
    .A(n_7727));
 AOI21xp5_ASAP7_75t_SL g205 (.A1(n_8406),
    .A2(n_22323),
    .B(n_20737),
    .Y(n_20738));
 NAND2xp5_ASAP7_75t_SL g20501 (.A(n_11871),
    .B(n_9501),
    .Y(n_11872));
 NAND2xp5_ASAP7_75t_SL g20502 (.A(n_22022),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_241),
    .Y(n_11871));
 INVx2_ASAP7_75t_SL g20510 (.A(n_11891),
    .Y(n_11892));
 XNOR2x1_ASAP7_75t_SL g20511 (.B(n_26078),
    .Y(n_11891),
    .A(n_11887));
 XOR2xp5_ASAP7_75t_SL g20517 (.A(n_19432),
    .B(n_23551),
    .Y(n_11896));
 AND2x2_ASAP7_75t_SL g20528 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_688),
    .Y(n_11904));
 AOI22x1_ASAP7_75t_SL g20535 (.A1(n_11914),
    .A2(n_11915),
    .B1(n_11913),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_126),
    .Y(n_11916));
 XOR2x2_ASAP7_75t_SL g20537 (.A(n_21137),
    .B(n_11912),
    .Y(n_11913));
 INVx1_ASAP7_75t_SL g20538 (.A(n_6409),
    .Y(n_11912));
 INVx1_ASAP7_75t_SL g20539 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_126),
    .Y(n_11915));
 NOR2xp33_ASAP7_75t_SL g20540 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_277),
    .B(n_11919),
    .Y(n_11920));
 NOR2x1_ASAP7_75t_SL g20541 (.A(n_10685),
    .B(n_11918),
    .Y(n_11919));
 XNOR2x1_ASAP7_75t_SL g20542 (.B(n_19490),
    .Y(n_11918),
    .A(n_21678));
 MAJIxp5_ASAP7_75t_L g20543_dup (.A(n_21046),
    .B(n_21048),
    .C(n_21049),
    .Y(n_14300));
 NAND2xp33_ASAP7_75t_SL g20547 (.A(n_7029),
    .B(n_7027),
    .Y(n_11924));
 INVx1_ASAP7_75t_SL g20548 (.A(n_20825),
    .Y(n_11925));
 OAI21x1_ASAP7_75t_SL g20549 (.A1(n_11928),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_272),
    .B(n_11931),
    .Y(n_11932));
 OA21x2_ASAP7_75t_SL g20550 (.A1(n_18004),
    .A2(n_18003),
    .B(n_8295),
    .Y(n_11928));
 AOI31xp67_ASAP7_75t_SL g20551 (.A1(n_18002),
    .A2(n_8295),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_272),
    .B(n_11930),
    .Y(n_11931));
 INVx1_ASAP7_75t_SL g20553 (.A(n_7595),
    .Y(n_11930));
 XNOR2xp5_ASAP7_75t_SL g20554 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_118),
    .B(n_20118),
    .Y(n_11936));
 XNOR2xp5_ASAP7_75t_SL g20558 (.A(n_11937),
    .B(n_19614),
    .Y(n_11941));
 INVx1_ASAP7_75t_SL g20559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_80),
    .Y(n_11937));
 MAJIxp5_ASAP7_75t_SL g20563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_62),
    .B(n_11942),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_26),
    .Y(n_11943));
 NAND2x1p5_ASAP7_75t_L g20564 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .Y(n_11942));
 XNOR2xp5_ASAP7_75t_SL g20566 (.A(n_12258),
    .B(n_11944),
    .Y(n_11945));
 OAI22xp5_ASAP7_75t_SL g20567 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_222),
    .A2(n_3511),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_226),
    .B2(n_3918),
    .Y(n_11944));
 XNOR2xp5_ASAP7_75t_SL g20577 (.A(n_24769),
    .B(n_11960),
    .Y(n_11961));
 XNOR2xp5_ASAP7_75t_SL g20579 (.A(n_12549),
    .B(n_21974),
    .Y(n_11960));
 XNOR2xp5_ASAP7_75t_SL g20583 (.A(n_11963),
    .B(n_21507),
    .Y(n_11970));
 XOR2xp5_ASAP7_75t_SL g20584 (.A(n_11962),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_252),
    .Y(n_11963));
 HB1xp67_ASAP7_75t_SL g20585 (.A(n_7071),
    .Y(n_11962));
 INVxp67_ASAP7_75t_SL g20587 (.A(n_11965),
    .Y(n_11966));
 NOR2x1_ASAP7_75t_SL g20588 (.A(n_11964),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_264),
    .Y(n_11965));
 BUFx2_ASAP7_75t_SL g20589 (.A(n_21986),
    .Y(n_11964));
 INVx1_ASAP7_75t_SL g20590 (.A(n_11967),
    .Y(n_11968));
 NAND2x1p5_ASAP7_75t_SL g20591 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_264),
    .B(n_11964),
    .Y(n_11967));
 MAJx2_ASAP7_75t_SL g20593 (.A(n_13708),
    .B(n_26003),
    .C(n_11972),
    .Y(n_9138));
 NAND2x1p5_ASAP7_75t_SL g20594 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .B(n_2820),
    .Y(n_11972));
 MAJIxp5_ASAP7_75t_SL g206 (.A(n_19143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_140),
    .Y(n_11515));
 XNOR2xp5_ASAP7_75t_SL g20615 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_711),
    .B(n_11997),
    .Y(n_11998));
 XOR2xp5_ASAP7_75t_SL g20616 (.A(n_11995),
    .B(n_11996),
    .Y(n_11997));
 NAND2xp5_ASAP7_75t_SL g20617 (.A(n_21789),
    .B(n_26238),
    .Y(n_11995));
 NAND2xp5_ASAP7_75t_SL g20619 (.A(n_14141),
    .B(n_2181),
    .Y(n_11996));
 MAJIxp5_ASAP7_75t_SL g20620 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_711),
    .B(n_11999),
    .C(n_12000),
    .Y(n_12001));
 INVxp67_ASAP7_75t_SL g20621 (.A(n_11995),
    .Y(n_11999));
 INVxp67_ASAP7_75t_SL g20622 (.A(n_11996),
    .Y(n_12000));
 NAND2xp5_ASAP7_75t_SL g20637 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .Y(n_12039));
 XOR2x2_ASAP7_75t_SL g20646 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_12),
    .B(n_12062),
    .Y(n_12063));
 XOR2xp5_ASAP7_75t_SL g20647 (.A(n_19677),
    .B(n_12061),
    .Y(n_12062));
 MAJx2_ASAP7_75t_SL g20654 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_12),
    .B(n_12064),
    .C(n_12065),
    .Y(n_12066));
 HB1xp67_ASAP7_75t_SL g20655 (.A(n_19677),
    .Y(n_12064));
 HB1xp67_ASAP7_75t_SL g20656 (.A(n_12061),
    .Y(n_12065));
 XNOR2xp5_ASAP7_75t_SL g20657 (.A(n_12067),
    .B(n_12068),
    .Y(n_12069));
 INVx1_ASAP7_75t_SL g20658 (.A(n_19674),
    .Y(n_12067));
 OAI22xp33_ASAP7_75t_SL g20659 (.A1(n_19676),
    .A2(n_19669),
    .B1(n_19675),
    .B2(n_19670),
    .Y(n_12068));
 INVx1_ASAP7_75t_SL g20667 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .Y(n_12073));
 XNOR2x1_ASAP7_75t_SL g20670 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_27),
    .Y(n_12077),
    .A(n_7435));
 HB1xp67_ASAP7_75t_SL g20672 (.A(n_12079),
    .Y(n_12080));
 XOR2xp5_ASAP7_75t_SL g20673 (.A(n_10456),
    .B(n_21142),
    .Y(n_12079));
 MAJIxp5_ASAP7_75t_SL g20676 (.A(n_4089),
    .B(n_8612),
    .C(n_12087),
    .Y(n_12088));
 INVx1_ASAP7_75t_SL g20677 (.A(n_12631),
    .Y(n_12087));
 MAJIxp5_ASAP7_75t_SL g207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_152),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_166),
    .C(n_11194),
    .Y(n_5781));
 MAJIxp5_ASAP7_75t_SL g20732 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_267),
    .B(n_6324),
    .C(n_10411),
    .Y(n_12186));
 XNOR2xp5_ASAP7_75t_SL g20735 (.A(n_12187),
    .B(n_12186),
    .Y(n_12188));
 INVx1_ASAP7_75t_SL g20736 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_51),
    .Y(n_12187));
 MAJIxp5_ASAP7_75t_SL g20762 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_178),
    .B(n_12217),
    .C(n_11534),
    .Y(n_12218));
 OAI22xp5_ASAP7_75t_SL g20786 (.A1(n_25599),
    .A2(n_12245),
    .B1(n_21793),
    .B2(n_19530),
    .Y(n_12246));
 INVx1_ASAP7_75t_SL g20793 (.A(n_19530),
    .Y(n_12250));
 OAI22xp5_ASAP7_75t_SL g20794 (.A1(n_18842),
    .A2(n_19530),
    .B1(n_12250),
    .B2(n_8766),
    .Y(n_12251));
 MAJIxp5_ASAP7_75t_SL g20796 (.A(n_12252),
    .B(n_26175),
    .C(n_12254),
    .Y(n_12255));
 INVxp67_ASAP7_75t_SL g20799 (.A(n_9120),
    .Y(n_12254));
 XOR2xp5_ASAP7_75t_SL g20803 (.A(n_12259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_332),
    .Y(n_12260));
 AOI21xp5_ASAP7_75t_SL g20804 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_250),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_263),
    .Y(n_12259));
 AND2x2_ASAP7_75t_L g20806 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_6965),
    .Y(n_12262));
 XOR2xp5_ASAP7_75t_SL g20808 (.A(n_12264),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_5),
    .Y(n_12265));
 OR2x2_ASAP7_75t_SL g20809 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_59),
    .Y(n_12264));
 OAI21x1_ASAP7_75t_SL g20815 (.A1(n_7007),
    .A2(n_12271),
    .B(n_7008),
    .Y(n_12272));
 OA21x2_ASAP7_75t_SL g20816 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_260),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_27),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_259),
    .Y(n_12271));
 XNOR2x1_ASAP7_75t_SL g20823 (.B(n_7250),
    .Y(n_12279),
    .A(n_7249));
 XNOR2xp5_ASAP7_75t_SL g20827 (.A(n_11891),
    .B(n_9238),
    .Y(n_12283));
 NAND2xp5_ASAP7_75t_SL g20828 (.A(n_11891),
    .B(n_9238),
    .Y(n_12284));
 XOR2xp5_ASAP7_75t_SL g20829 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_96),
    .B(n_12039),
    .Y(n_12285));
 NOR2xp33_ASAP7_75t_SL g20831 (.A(n_15084),
    .B(n_15085),
    .Y(n_12287));
 XOR2xp5_ASAP7_75t_SL g20832 (.A(n_13061),
    .B(n_6593),
    .Y(n_12288));
 XOR2xp5_ASAP7_75t_SL g20833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_36),
    .Y(n_12289));
 XNOR2xp5_ASAP7_75t_SL g20836 (.A(n_18699),
    .B(n_12303),
    .Y(n_12304));
 MAJIxp5_ASAP7_75t_SL g20841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_41),
    .Y(n_12293));
 XNOR2xp5_ASAP7_75t_SL g20843 (.A(n_12301),
    .B(n_19773),
    .Y(n_12303));
 INVxp67_ASAP7_75t_SL g20844 (.A(n_19183),
    .Y(n_12301));
 XNOR2xp5_ASAP7_75t_SL g20850 (.A(n_12306),
    .B(n_12307),
    .Y(n_12308));
 INVxp67_ASAP7_75t_SL g20851 (.A(n_14741),
    .Y(n_12306));
 AOI22xp5_ASAP7_75t_SL g20853 (.A1(n_7297),
    .A2(n_14746),
    .B1(n_7296),
    .B2(n_14749),
    .Y(n_12307));
 NAND2xp5_ASAP7_75t_SL g20887 (.A(n_12375),
    .B(n_21364),
    .Y(n_12376));
 INVxp67_ASAP7_75t_SL g20888 (.A(n_12374),
    .Y(n_12375));
 NAND2xp5_ASAP7_75t_SL g20889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_23),
    .Y(n_12374));
 OA21x2_ASAP7_75t_SL g20890 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_232),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_240),
    .Y(n_12379));
 INVx1_ASAP7_75t_SL g20891 (.A(n_12377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_240));
 NOR2xp67_ASAP7_75t_SL g20892 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_174),
    .Y(n_12377));
 OAI21xp5_ASAP7_75t_SL g20893 (.A1(n_12377),
    .A2(n_12382),
    .B(n_12383),
    .Y(n_12384));
 NAND2xp5_ASAP7_75t_SL g20894 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_3150),
    .Y(n_12387));
 MAJIxp5_ASAP7_75t_SL g20895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_43),
    .Y(n_12388));
 AOI21x1_ASAP7_75t_SL g20897 (.A1(n_9384),
    .A2(n_18753),
    .B(n_9385),
    .Y(n_12393));
 NOR2xp67_ASAP7_75t_SL g20898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_224),
    .Y(n_12395));
 XOR2x2_ASAP7_75t_SL g209 (.A(n_12219),
    .B(n_6360),
    .Y(n_6361));
 MAJx2_ASAP7_75t_SL g20902 (.A(n_12397),
    .B(n_12398),
    .C(n_12400),
    .Y(n_12402));
 NAND2xp5_ASAP7_75t_SL g20904 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_99),
    .Y(n_12398));
 MAJIxp5_ASAP7_75t_SL g20906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_55),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_74),
    .Y(n_12400));
 MAJIxp5_ASAP7_75t_SL g20915 (.A(n_13880),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_134),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_126),
    .Y(n_12414));
 MAJIxp5_ASAP7_75t_SL g20917 (.A(n_12419),
    .B(n_12420),
    .C(n_12422),
    .Y(n_12424));
 XOR2x2_ASAP7_75t_SL g20918 (.A(n_18978),
    .B(n_12418),
    .Y(n_12419));
 MAJIxp5_ASAP7_75t_SL g20919 (.A(n_13495),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_49),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_40),
    .Y(n_12418));
 MAJIxp5_ASAP7_75t_SL g20921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_45),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_95),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_76),
    .Y(n_12420));
 XNOR2xp5_ASAP7_75t_SL g20923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_98),
    .B(n_11753),
    .Y(n_12422));
 MAJIxp5_ASAP7_75t_SL g20925 (.A(n_12418),
    .B(n_12425),
    .C(n_12427),
    .Y(n_12428));
 NAND2x1_ASAP7_75t_SL g20927 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .B(n_2544),
    .Y(n_12425));
 AND2x2_ASAP7_75t_SL g20928 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(n_2831),
    .Y(n_12427));
 AOI21xp5_ASAP7_75t_SL g20938 (.A1(n_12500),
    .A2(n_19496),
    .B(n_19504),
    .Y(n_12510));
 OAI21xp33_ASAP7_75t_SL g20939 (.A1(n_21577),
    .A2(n_16397),
    .B(n_12499),
    .Y(n_12500));
 INVx1_ASAP7_75t_SL g20945 (.A(n_22497),
    .Y(n_12503));
 MAJIxp5_ASAP7_75t_SL g20947 (.A(n_11761),
    .B(n_10617),
    .C(n_21229),
    .Y(n_12504));
 INVx1_ASAP7_75t_SL g20949 (.A(n_12504),
    .Y(n_12508));
 INVxp67_ASAP7_75t_SL g20950 (.A(n_19496),
    .Y(n_12512));
 AOI21xp5_ASAP7_75t_SL g20951 (.A1(n_12494),
    .A2(n_12513),
    .B(n_12498),
    .Y(n_12514));
 NOR2x1_ASAP7_75t_SL g20953 (.A(n_21534),
    .B(n_12531),
    .Y(n_12532));
 INVxp67_ASAP7_75t_SL g20957 (.A(n_5815),
    .Y(n_12516));
 MAJIxp5_ASAP7_75t_SL g20959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_69),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_106),
    .Y(n_12518));
 XOR2xp5_ASAP7_75t_SL g20961 (.A(n_8416),
    .B(n_8414),
    .Y(n_12520));
 XNOR2x2_ASAP7_75t_SL g20962 (.A(n_12527),
    .B(n_12530),
    .Y(n_12531));
 XNOR2xp5_ASAP7_75t_SL g20963 (.A(n_5817),
    .B(n_12526),
    .Y(n_12527));
 MAJIxp5_ASAP7_75t_SL g20964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_135),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_129),
    .C(n_5815),
    .Y(n_5817));
 XNOR2xp5_ASAP7_75t_SL g20965 (.A(n_12525),
    .B(n_12265),
    .Y(n_12526));
 INVxp67_ASAP7_75t_SL g20966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_141),
    .Y(n_12525));
 XNOR2xp5_ASAP7_75t_SL g20967 (.A(n_12528),
    .B(n_18952),
    .Y(n_12530));
 OAI21x1_ASAP7_75t_SL g20968 (.A1(n_8421),
    .A2(n_8415),
    .B(n_8422),
    .Y(n_12528));
 AND2x2_ASAP7_75t_SL g20979 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_678),
    .Y(n_12540));
 NOR2xp33_ASAP7_75t_SL g20982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_297),
    .B(n_12546),
    .Y(n_12547));
 INVxp33_ASAP7_75t_SRAM g20983 (.A(n_12888),
    .Y(n_12546));
 XOR2xp5_ASAP7_75t_SL g20985 (.A(n_12548),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_170),
    .Y(n_12549));
 XNOR2x1_ASAP7_75t_SL g20986 (.B(n_21056),
    .Y(n_12548),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_140));
 AND2x2_ASAP7_75t_SL g20989 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_576),
    .B(n_2159),
    .Y(n_12550));
 AOI21x1_ASAP7_75t_SL g20994 (.A1(n_18785),
    .A2(n_12559),
    .B(n_12560),
    .Y(n_12561));
 HB1xp67_ASAP7_75t_SL g20996 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_296),
    .Y(n_12559));
 HB1xp67_ASAP7_75t_SL g20997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_299),
    .Y(n_12560));
 AOI21xp5_ASAP7_75t_SL g20998 (.A1(n_4771),
    .A2(n_4772),
    .B(n_4773),
    .Y(n_12562));
 OAI21x1_ASAP7_75t_SL g20999 (.A1(n_12563),
    .A2(n_12564),
    .B(n_2176),
    .Y(n_12565));
 NAND2xp5_ASAP7_75t_SL g21 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(n_9349),
    .Y(n_9571));
 INVx1_ASAP7_75t_SL g210 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_178),
    .Y(n_6360));
 AND2x2_ASAP7_75t_SL g21000 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_309),
    .B(n_5589),
    .Y(n_12563));
 NOR2xp33_ASAP7_75t_SL g21001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_309),
    .B(n_5589),
    .Y(n_12564));
 OAI21xp5_ASAP7_75t_SL g21002 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_283),
    .A2(n_13934),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_281),
    .Y(n_12567));
 XNOR2x1_ASAP7_75t_SL g21006 (.B(n_12570),
    .Y(n_12571),
    .A(n_9813));
 XNOR2x1_ASAP7_75t_SL g21007 (.B(n_9811),
    .Y(n_12570),
    .A(n_23422));
 XNOR2x1_ASAP7_75t_SL g21008 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_132),
    .Y(n_12575),
    .A(n_18986));
 XNOR2xp5_ASAP7_75t_SL g21013 (.A(n_21295),
    .B(n_19688),
    .Y(n_12576));
 XNOR2x1_ASAP7_75t_SL g21014 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_145),
    .Y(n_12580),
    .A(n_12579));
 INVx1_ASAP7_75t_SL g21015 (.A(n_12578),
    .Y(n_12579));
 NAND2xp5_ASAP7_75t_SL g21016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_106),
    .B(n_13240),
    .Y(n_12578));
 NAND2xp5_ASAP7_75t_SL g21017 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .Y(n_12581));
 XOR2xp5_ASAP7_75t_SL g21019 (.A(n_12583),
    .B(n_12593),
    .Y(n_12594));
 XOR2x2_ASAP7_75t_SL g21020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_188),
    .Y(n_12583));
 AO21x1_ASAP7_75t_SL g21021 (.A1(n_12589),
    .A2(n_12591),
    .B(n_12592),
    .Y(n_12593));
 NAND2xp5_ASAP7_75t_SL g21022 (.A(n_23002),
    .B(n_18987),
    .Y(n_12589));
 INVx1_ASAP7_75t_SL g21024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_98),
    .Y(n_12584));
 INVxp67_ASAP7_75t_SL g21027 (.A(n_21976),
    .Y(n_12591));
 NOR2x1_ASAP7_75t_SL g21029 (.A(n_18987),
    .B(n_23002),
    .Y(n_12592));
 XNOR2xp5_ASAP7_75t_SL g21030 (.A(n_12598),
    .B(n_12605),
    .Y(n_12606));
 INVx1_ASAP7_75t_SL g21031 (.A(n_12597),
    .Y(n_12598));
 XNOR2xp5_ASAP7_75t_SL g21032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_6),
    .Y(n_12597));
 AOI22xp5_ASAP7_75t_SL g21033 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_199),
    .A2(n_12604),
    .B1(n_19185),
    .B2(n_12603),
    .Y(n_12605));
 XOR2x2_ASAP7_75t_SL g21038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_149),
    .B(n_23432),
    .Y(n_12603));
 XNOR2xp5_ASAP7_75t_SL g21047 (.A(n_12618),
    .B(n_14723),
    .Y(n_12620));
 XOR2xp5_ASAP7_75t_SL g21048 (.A(n_12616),
    .B(n_15097),
    .Y(n_12618));
 XNOR2xp5_ASAP7_75t_SL g21051 (.A(n_12623),
    .B(n_12624),
    .Y(n_12625));
 NAND2x1_ASAP7_75t_SL g21052 (.A(n_12621),
    .B(n_12622),
    .Y(n_12623));
 NAND2xp5_ASAP7_75t_SL g21053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_0),
    .Y(n_12621));
 OR2x2_ASAP7_75t_SL g21054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_0),
    .Y(n_12622));
 MAJIxp5_ASAP7_75t_SL g21055 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_30),
    .C(n_21797),
    .Y(n_12624));
 MAJIxp5_ASAP7_75t_SL g21059 (.A(n_11431),
    .B(n_22312),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_581),
    .Y(n_9966));
 XNOR2xp5_ASAP7_75t_SL g21062 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_23),
    .B(n_12073),
    .Y(n_12631));
 MAJx2_ASAP7_75t_SL g21065 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_262),
    .B(n_6411),
    .C(n_23670),
    .Y(n_12632));
 XOR2xp5_ASAP7_75t_SL g21066 (.A(n_13072),
    .B(n_8605),
    .Y(n_12634));
 XNOR2xp5_ASAP7_75t_SL g21067 (.A(n_12637),
    .B(n_12641),
    .Y(n_12642));
 NAND2xp5_ASAP7_75t_SL g21068 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_265),
    .Y(n_12637));
 OAI21xp5_ASAP7_75t_SL g21069 (.A1(n_21961),
    .A2(n_12639),
    .B(n_12640),
    .Y(n_12641));
 NOR2x2_ASAP7_75t_SRAM g21071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_249),
    .Y(n_12639));
 NAND2xp5_ASAP7_75t_SL g21072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_249),
    .Y(n_12640));
 MAJx2_ASAP7_75t_SL g21078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_172),
    .Y(n_12648));
 INVx1_ASAP7_75t_SL g21079 (.A(n_12648),
    .Y(n_12649));
 XNOR2xp5_ASAP7_75t_SL g21080 (.A(n_12652),
    .B(n_20101),
    .Y(n_12658));
 MAJIxp5_ASAP7_75t_SL g21082 (.A(n_5393),
    .B(n_17552),
    .C(n_8674),
    .Y(n_12653));
 INVx1_ASAP7_75t_SL g21085 (.A(n_12652),
    .Y(n_12659));
 XNOR2xp5_ASAP7_75t_SL g21087 (.A(n_12665),
    .B(n_12664),
    .Y(n_12666));
 XOR2xp5_ASAP7_75t_SL g21088 (.A(n_12661),
    .B(n_12663),
    .Y(n_12664));
 MAJx2_ASAP7_75t_SL g21089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_187),
    .B(n_3204),
    .C(n_2801),
    .Y(n_12661));
 XNOR2xp5_ASAP7_75t_SL g21090 (.A(n_12662),
    .B(n_10069),
    .Y(n_12663));
 INVx1_ASAP7_75t_SL g21091 (.A(n_19964),
    .Y(n_12662));
 MAJIxp5_ASAP7_75t_SL g21092 (.A(n_20306),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_29),
    .C(n_3360),
    .Y(n_12665));
 INVx1_ASAP7_75t_SL g211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_191),
    .Y(n_7338));
 AOI31xp67_ASAP7_75t_SL g21102 (.A1(n_12696),
    .A2(n_12697),
    .A3(n_12701),
    .B(n_12704),
    .Y(n_12705));
 AOI221xp5_ASAP7_75t_SL g21104 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .B1(n_12702),
    .B2(n_12703),
    .C(n_12700),
    .Y(n_12704));
 INVx1_ASAP7_75t_SL g21105 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .Y(n_12703));
 HB1xp67_ASAP7_75t_SL g21106 (.A(n_12705),
    .Y(n_12706));
 XNOR2xp5_ASAP7_75t_SL g21107 (.A(n_12709),
    .B(n_18992),
    .Y(n_12715));
 INVxp67_ASAP7_75t_SL g21108 (.A(n_12708),
    .Y(n_12709));
 AOI21x1_ASAP7_75t_SL g21109 (.A1(n_11112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_128),
    .Y(n_12708));
 XNOR2x2_ASAP7_75t_SL g21113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_0),
    .Y(n_12712));
 AO21x1_ASAP7_75t_SL g21117 (.A1(n_12717),
    .A2(n_21624),
    .B(n_12719),
    .Y(n_12720));
 NAND2xp5_ASAP7_75t_SL g21118 (.A(n_21334),
    .B(n_7116),
    .Y(n_12717));
 NOR2xp67_ASAP7_75t_SL g21120 (.A(n_21334),
    .B(n_7116),
    .Y(n_12719));
 NOR2xp67_ASAP7_75t_SL g21124 (.A(n_12738),
    .B(n_12744),
    .Y(n_12745));
 MAJIxp5_ASAP7_75t_SL g21125 (.A(n_7480),
    .B(n_7481),
    .C(n_7482),
    .Y(n_12738));
 XNOR2x1_ASAP7_75t_SL g21126 (.B(n_18993),
    .Y(n_12744),
    .A(n_12740));
 XNOR2xp5_ASAP7_75t_SL g21127 (.A(n_12739),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_168),
    .Y(n_12740));
 INVx1_ASAP7_75t_SL g21128 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_1),
    .Y(n_12739));
 INVx1_ASAP7_75t_SL g21132 (.A(n_12740),
    .Y(n_12746));
 XNOR2x1_ASAP7_75t_SL g21133 (.B(n_21925),
    .Y(n_12754),
    .A(n_12747));
 AND2x2_ASAP7_75t_SL g21134 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_546),
    .Y(n_12747));
 NAND2xp5_ASAP7_75t_SL g21136 (.A(n_12748),
    .B(n_12749),
    .Y(n_12750));
 AND3x4_ASAP7_75t_SL g21137 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[6]),
    .Y(n_12748));
 INVx1_ASAP7_75t_SL g21138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_226),
    .Y(n_12749));
 NAND2xp5_ASAP7_75t_SL g21140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_226),
    .B(n_12748),
    .Y(n_12752));
 XNOR2x1_ASAP7_75t_SL g21160 (.B(n_12786),
    .Y(n_12787),
    .A(n_12785));
 NOR2x1p5_ASAP7_75t_SL g21161 (.A(n_12782),
    .B(n_14736),
    .Y(n_12785));
 INVxp67_ASAP7_75t_SL g21162 (.A(n_12781),
    .Y(n_12782));
 AND3x1_ASAP7_75t_SL g21163 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[2]),
    .Y(n_12781));
 OAI21x1_ASAP7_75t_SL g21166 (.A1(n_11723),
    .A2(n_11722),
    .B(n_2158),
    .Y(n_12786));
 XNOR2xp5_ASAP7_75t_SL g21175 (.A(n_12801),
    .B(n_12802),
    .Y(n_12803));
 NAND2xp5_ASAP7_75t_SL g21176 (.A(n_12800),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .Y(n_12801));
 NAND2x1_ASAP7_75t_SL g21177 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(n_14985),
    .Y(n_12802));
 NOR2xp33_ASAP7_75t_SL g21178 (.A(n_146),
    .B(n_3433),
    .Y(n_12806));
 XNOR2xp5_ASAP7_75t_SL g21181 (.A(n_19186),
    .B(n_19187),
    .Y(n_12817));
 XNOR2xp5_ASAP7_75t_SL g21186 (.A(n_12833),
    .B(n_21802),
    .Y(n_12839));
 INVx1_ASAP7_75t_SL g21187 (.A(n_15719),
    .Y(n_12833));
 INVxp67_ASAP7_75t_SL g21189 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_755),
    .Y(n_12831));
 XOR2x2_ASAP7_75t_SL g21192 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_6),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_723),
    .Y(n_12834));
 XNOR2xp5_ASAP7_75t_SL g212 (.A(n_7404),
    .B(n_7405),
    .Y(n_7406));
 MAJIxp5_ASAP7_75t_SL g21223 (.A(n_12882),
    .B(n_12884),
    .C(n_10173),
    .Y(n_12887));
 XOR2xp5_ASAP7_75t_SL g21224 (.A(n_12878),
    .B(n_18996),
    .Y(n_12882));
 AND2x2_ASAP7_75t_SL g21225 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_720),
    .Y(n_12878));
 MAJIxp5_ASAP7_75t_SL g21230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_755),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_691),
    .Y(n_12884));
 XNOR2x1_ASAP7_75t_SL g21232 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_753),
    .Y(n_10173),
    .A(n_17734));
 NAND2xp5_ASAP7_75t_SL g21233 (.A(n_12888),
    .B(n_14090),
    .Y(n_12892));
 NAND2xp5_ASAP7_75t_SL g21234 (.A(n_11945),
    .B(n_14091),
    .Y(n_12888));
 MAJIxp5_ASAP7_75t_SL g21238 (.A(n_12893),
    .B(n_12894),
    .C(n_12899),
    .Y(n_12900));
 XNOR2xp5_ASAP7_75t_SL g21239 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_113),
    .Y(n_12893));
 XNOR2xp5_ASAP7_75t_SL g21240 (.A(n_15798),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_6),
    .Y(n_12894));
 MAJIxp5_ASAP7_75t_SL g21241 (.A(n_12895),
    .B(n_12896),
    .C(n_12897),
    .Y(n_12899));
 NAND2xp5_ASAP7_75t_SL g21242 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_61),
    .Y(n_12895));
 NAND2x1_ASAP7_75t_SL g21243 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .B(n_2831),
    .Y(n_12896));
 NAND2xp5_ASAP7_75t_SL g21245 (.A(n_23016),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .Y(n_12897));
 MAJIxp5_ASAP7_75t_SL g21247 (.A(n_12902),
    .B(n_12903),
    .C(n_12904),
    .Y(n_12905));
 INVx2_ASAP7_75t_SL g21248 (.A(n_12901),
    .Y(n_12902));
 NAND2x1_ASAP7_75t_SL g21249 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(n_3479),
    .Y(n_12901));
 NAND2x1_ASAP7_75t_SL g21250 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .Y(n_12903));
 AND2x2_ASAP7_75t_SL g21251 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(n_2927),
    .Y(n_12904));
 MAJx2_ASAP7_75t_SL g21252 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_21),
    .C(n_22870),
    .Y(n_12906));
 NOR2x1_ASAP7_75t_SL g21256 (.A(n_19189),
    .B(n_12922),
    .Y(n_12923));
 XNOR2xp5_ASAP7_75t_SL g21262 (.A(n_12918),
    .B(n_18999),
    .Y(n_12922));
 INVxp67_ASAP7_75t_SL g21263 (.A(n_12917),
    .Y(n_12918));
 MAJIxp5_ASAP7_75t_SL g21264 (.A(n_21497),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_86),
    .C(n_21546),
    .Y(n_12917));
 XNOR2x1_ASAP7_75t_SL g21269 (.B(n_12928),
    .Y(n_12929),
    .A(n_12924));
 NAND2xp5_ASAP7_75t_SL g21271 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .B(n_2855),
    .Y(n_12924));
 XOR2xp5_ASAP7_75t_SL g21272 (.A(n_12926),
    .B(n_12927),
    .Y(n_12928));
 NAND2x1_ASAP7_75t_SL g21273 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(n_2325),
    .Y(n_12926));
 NAND2x1_ASAP7_75t_L g21274 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .B(n_6965),
    .Y(n_12927));
 XNOR2xp5_ASAP7_75t_SL g21275 (.A(n_12930),
    .B(n_12933),
    .Y(n_12934));
 NAND2x1_ASAP7_75t_SL g21276 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .Y(n_12930));
 XOR2xp5_ASAP7_75t_SL g21277 (.A(n_12931),
    .B(n_12932),
    .Y(n_12933));
 NAND2xp5_ASAP7_75t_SL g21278 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(n_4831),
    .Y(n_12931));
 AND2x2_ASAP7_75t_SL g21279 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_18039),
    .Y(n_12932));
 INVx1_ASAP7_75t_SL g21280 (.A(n_12931),
    .Y(n_12935));
 OAI22xp5_ASAP7_75t_SL g21284 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_81),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_19),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_82),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_132),
    .Y(n_12938));
 XNOR2xp5_ASAP7_75t_SL g21287 (.A(n_12940),
    .B(n_19001),
    .Y(n_12945));
 INVx1_ASAP7_75t_SL g21288 (.A(n_12939),
    .Y(n_12940));
 NAND2xp5_ASAP7_75t_SL g21289 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .B(n_2544),
    .Y(n_12939));
 INVx1_ASAP7_75t_SL g213 (.A(n_7403),
    .Y(n_7404));
 XNOR2x2_ASAP7_75t_SL g21303 (.A(n_11401),
    .B(n_11405),
    .Y(n_12956));
 XNOR2x1_ASAP7_75t_SL g21305 (.B(n_23541),
    .Y(n_12962),
    .A(n_12959));
 MAJIxp5_ASAP7_75t_SL g21306 (.A(n_11729),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_52),
    .C(n_3950),
    .Y(n_12959));
 INVxp33_ASAP7_75t_SL g21312 (.A(n_23541),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_176));
 AND2x2_ASAP7_75t_SL g21317 (.A(n_2168),
    .B(n_2160),
    .Y(n_12979));
 AND2x2_ASAP7_75t_SL g21319 (.A(n_12511),
    .B(n_2168),
    .Y(n_12986));
 XNOR2x1_ASAP7_75t_SL g21320 (.B(n_12995),
    .Y(n_12996),
    .A(n_14812));
 OR2x2_ASAP7_75t_SL g21322 (.A(n_12990),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_279),
    .Y(n_12991));
 NAND2xp5_ASAP7_75t_SL g21326 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_279),
    .Y(n_12993));
 NAND2xp5_ASAP7_75t_SL g21327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_562),
    .B(n_2182),
    .Y(n_12995));
 INVxp67_ASAP7_75t_SRAM g21328 (.A(n_12995),
    .Y(n_12997));
 OAI21xp5_ASAP7_75t_SL g21338 (.A1(n_13013),
    .A2(n_13011),
    .B(n_13015),
    .Y(n_13016));
 AOI21x1_ASAP7_75t_SL g21339 (.A1(n_13007),
    .A2(n_13008),
    .B(n_13010),
    .Y(n_13011));
 NOR2x1_ASAP7_75t_SL g21340 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_290),
    .B(n_14135),
    .Y(n_13007));
 NAND2x2_ASAP7_75t_SL g21341 (.A(n_6025),
    .B(n_13458),
    .Y(n_13008));
 INVxp67_ASAP7_75t_SL g21342 (.A(n_13009),
    .Y(n_13010));
 OAI21xp5_ASAP7_75t_SL g21343 (.A1(n_14136),
    .A2(n_23103),
    .B(n_23102),
    .Y(n_13009));
 NOR2xp67_ASAP7_75t_SL g21345 (.A(n_23105),
    .B(n_22967),
    .Y(n_13012));
 NAND2xp5_ASAP7_75t_SL g21346 (.A(n_22967),
    .B(n_23105),
    .Y(n_13014));
 XNOR2xp5_ASAP7_75t_SL g21347 (.A(n_13017),
    .B(n_21613),
    .Y(n_13025));
 XOR2xp5_ASAP7_75t_SL g21348 (.A(n_18846),
    .B(n_15231),
    .Y(n_13017));
 XNOR2x2_ASAP7_75t_SL g21352 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_15),
    .Y(n_13021));
 INVxp67_ASAP7_75t_SL g21354 (.A(n_13022),
    .Y(n_13023));
 MAJIxp5_ASAP7_75t_SL g21355 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_103),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_78),
    .Y(n_13022));
 INVxp67_ASAP7_75t_SL g21356 (.A(n_13017),
    .Y(n_5719));
 OAI21x1_ASAP7_75t_SL g21359 (.A1(n_13028),
    .A2(n_19525),
    .B(n_13030),
    .Y(n_13031));
 AND2x2_ASAP7_75t_SL g21360 (.A(n_19523),
    .B(n_20239),
    .Y(n_13028));
 AND3x2_ASAP7_75t_SL g21362 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[2]),
    .Y(n_13030));
 XNOR2xp5_ASAP7_75t_SL g21363 (.A(n_13034),
    .B(n_21634),
    .Y(n_13040));
 XNOR2x2_ASAP7_75t_SL g21364 (.A(n_13033),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_199),
    .Y(n_13034));
 INVxp67_ASAP7_75t_SL g21365 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_189),
    .Y(n_13033));
 XNOR2x1_ASAP7_75t_SL g21368 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_194),
    .Y(n_13036),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_149));
 INVx2_ASAP7_75t_SL g21370 (.A(n_13036),
    .Y(n_13038));
 OAI22xp5_ASAP7_75t_SL g21383 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_109),
    .A2(n_13052),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_110),
    .B2(n_13053),
    .Y(n_13054));
 NAND2x1_ASAP7_75t_SL g21384 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(n_3479),
    .Y(n_13052));
 INVx2_ASAP7_75t_SL g21385 (.A(n_13052),
    .Y(n_13053));
 MAJIxp5_ASAP7_75t_SL g21386 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_109),
    .C(n_13053),
    .Y(n_13056));
 INVx1_ASAP7_75t_SL g21388 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_705),
    .Y(n_13057));
 XNOR2xp5_ASAP7_75t_SL g21389 (.A(n_18157),
    .B(n_13060),
    .Y(n_13061));
 OAI22xp5_ASAP7_75t_SL g21390 (.A1(n_19868),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_135),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .B2(n_13059),
    .Y(n_13060));
 INVx2_ASAP7_75t_SL g21391 (.A(n_19868),
    .Y(n_13059));
 OAI22xp5_ASAP7_75t_SL g21392 (.A1(n_23389),
    .A2(n_19868),
    .B1(n_23393),
    .B2(n_13059),
    .Y(n_6045));
 MAJx2_ASAP7_75t_SL g21396 (.A(n_8605),
    .B(n_3657),
    .C(n_13065),
    .Y(n_13067));
 XOR2x2_ASAP7_75t_SL g21398 (.A(n_26076),
    .B(n_22180),
    .Y(n_13065));
 MAJIxp5_ASAP7_75t_SL g214 (.A(n_13667),
    .B(n_7402),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_298),
    .Y(n_7403));
 INVxp67_ASAP7_75t_SL g21400 (.A(n_13067),
    .Y(n_13069));
 OAI22xp5_ASAP7_75t_SL g21401 (.A1(n_13071),
    .A2(n_3657),
    .B1(n_8606),
    .B2(n_13065),
    .Y(n_13072));
 INVx1_ASAP7_75t_SL g21402 (.A(n_13065),
    .Y(n_13071));
 NAND2xp5_ASAP7_75t_SL g21409 (.A(n_13080),
    .B(n_10922),
    .Y(n_13081));
 XOR2xp5_ASAP7_75t_SL g21410 (.A(n_22188),
    .B(n_13079),
    .Y(n_13080));
 XNOR2xp5_ASAP7_75t_SL g21411 (.A(n_26101),
    .B(n_10760),
    .Y(n_13079));
 NOR2x1_ASAP7_75t_SL g21412 (.A(n_10922),
    .B(n_13080),
    .Y(n_13082));
 OAI21xp5_ASAP7_75t_SL g21417 (.A1(n_13088),
    .A2(n_11790),
    .B(n_13089),
    .Y(n_13090));
 NOR2xp33_ASAP7_75t_SL g21418 (.A(n_13087),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_269),
    .Y(n_13088));
 XNOR2xp5_ASAP7_75t_SL g21419 (.A(n_22419),
    .B(n_11517),
    .Y(n_13087));
 NAND2xp5_ASAP7_75t_SL g21420 (.A(n_13087),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_269),
    .Y(n_13089));
 NOR2xp33_ASAP7_75t_SRAM g21421 (.A(n_13088),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_290),
    .Y(n_13091));
 OAI21x1_ASAP7_75t_SL g21427 (.A1(n_9053),
    .A2(n_24766),
    .B(n_9054),
    .Y(n_13097));
 XNOR2xp5_ASAP7_75t_SL g21430 (.A(n_13098),
    .B(n_18935),
    .Y(n_13100));
 INVx1_ASAP7_75t_SL g21431 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_74),
    .Y(n_13098));
 MAJIxp5_ASAP7_75t_SL g21433 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_224),
    .B(n_13103),
    .C(n_13106),
    .Y(n_13107));
 HB1xp67_ASAP7_75t_SL g21434 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_190),
    .Y(n_13103));
 XNOR2xp5_ASAP7_75t_SL g21435 (.A(n_13104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_195),
    .Y(n_13106));
 XOR2x2_ASAP7_75t_SL g21436 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_56),
    .Y(n_13104));
 XNOR2xp5_ASAP7_75t_SL g21438 (.A(n_13104),
    .B(n_19006),
    .Y(n_13111));
 MAJIxp5_ASAP7_75t_SL g21441 (.A(n_21588),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_77),
    .C(n_13104),
    .Y(n_13112));
 MAJIxp5_ASAP7_75t_SL g21448 (.A(n_13124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_135),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_121),
    .Y(n_13125));
 XNOR2x1_ASAP7_75t_SL g21449 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_91),
    .Y(n_13123),
    .A(n_19449));
 XNOR2xp5_ASAP7_75t_SL g21454 (.A(n_8261),
    .B(n_13123),
    .Y(n_13126));
 NOR2x1_ASAP7_75t_SL g21455 (.A(n_22295),
    .B(n_13129),
    .Y(n_13130));
 XNOR2x2_ASAP7_75t_SL g21456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_232),
    .B(n_13128),
    .Y(n_13129));
 XNOR2xp5_ASAP7_75t_SL g21457 (.A(n_13127),
    .B(n_10294),
    .Y(n_13128));
 INVx1_ASAP7_75t_SL g21458 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_219),
    .Y(n_13127));
 INVxp67_ASAP7_75t_SL g21466 (.A(n_19007),
    .Y(n_13138));
 A2O1A1Ixp33_ASAP7_75t_SL g21467 (.A1(n_22422),
    .A2(n_19007),
    .B(n_13141),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_119),
    .Y(n_13142));
 NOR2xp33_ASAP7_75t_SL g21469 (.A(n_22422),
    .B(n_19007),
    .Y(n_13141));
 XNOR2xp5_ASAP7_75t_SL g21470 (.A(n_13143),
    .B(n_19008),
    .Y(n_13148));
 INVx1_ASAP7_75t_SL g21471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_112),
    .Y(n_13143));
 NAND2x1_ASAP7_75t_SL g21473 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(n_2820),
    .Y(n_13144));
 MAJIxp5_ASAP7_75t_SL g21476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_112),
    .C(n_13144),
    .Y(n_13149));
 MAJIxp5_ASAP7_75t_SL g215 (.A(n_26152),
    .B(n_22235),
    .C(n_22234),
    .Y(n_21976));
 NAND3x2_ASAP7_75t_L g21534 (.B(n_22250),
    .C(n_2657),
    .Y(n_13233),
    .A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]));
 XNOR2xp5_ASAP7_75t_SL g21595 (.A(n_13293),
    .B(n_11823),
    .Y(n_13294));
 XNOR2xp5_ASAP7_75t_SL g21596 (.A(n_15589),
    .B(n_13292),
    .Y(n_13293));
 MAJIxp5_ASAP7_75t_SL g21598 (.A(n_13293),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_157),
    .Y(n_13295));
 MAJIxp5_ASAP7_75t_SL g216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_46),
    .B(n_22874),
    .C(n_12154),
    .Y(n_19252));
 MAJx2_ASAP7_75t_SL g21622 (.A(n_18665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_132),
    .C(n_25992),
    .Y(n_13321));
 XOR2xp5_ASAP7_75t_SL g21626 (.A(n_9810),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_54),
    .Y(n_13324));
 XOR2xp5_ASAP7_75t_SL g21629 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_40),
    .Y(n_13327));
 XNOR2xp5_ASAP7_75t_SL g21632 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_8),
    .B(n_10299),
    .Y(n_13330));
 XOR2x2_ASAP7_75t_SL g21634 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_177),
    .B(n_12293),
    .Y(n_13332));
 XOR2xp5_ASAP7_75t_SL g21635 (.A(n_8594),
    .B(n_8596),
    .Y(n_13333));
 XNOR2xp5_ASAP7_75t_SL g21654 (.A(n_9713),
    .B(n_13358),
    .Y(n_13359));
 MAJIxp5_ASAP7_75t_SL g21655 (.A(n_10643),
    .B(n_9714),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_152),
    .Y(n_13358));
 XOR2x2_ASAP7_75t_SL g21656 (.A(n_6824),
    .B(n_13360),
    .Y(n_13361));
 AOI22xp5_ASAP7_75t_SL g21657 (.A1(n_13295),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_204),
    .B1(n_6825),
    .B2(n_15213),
    .Y(n_13360));
 NOR2xp33_ASAP7_75t_SL g21658 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283),
    .B(n_13362),
    .Y(n_13363));
 NOR2x1_ASAP7_75t_SL g21659 (.A(n_7670),
    .B(n_20974),
    .Y(n_13362));
 XOR2x2_ASAP7_75t_SL g21679 (.A(n_22174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_105),
    .Y(n_13387));
 NAND2xp5_ASAP7_75t_SL g21685 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_209),
    .B(n_23415),
    .Y(n_13389));
 NOR2xp67_ASAP7_75t_SL g21686 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_209),
    .B(n_23415),
    .Y(n_13390));
 XNOR2xp5_ASAP7_75t_SL g21687 (.A(n_5494),
    .B(n_13589),
    .Y(n_13397));
 INVx1_ASAP7_75t_SL g21689 (.A(n_21977),
    .Y(n_13393));
 XOR2xp5_ASAP7_75t_SL g21692 (.A(n_4041),
    .B(n_18988),
    .Y(n_13401));
 XNOR2xp5_ASAP7_75t_SL g21696 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_225),
    .B(n_13404),
    .Y(n_13405));
 AOI21xp5_ASAP7_75t_SL g21697 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_298),
    .A2(n_22596),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_301),
    .Y(n_13404));
 XNOR2xp5_ASAP7_75t_SL g217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_189),
    .Y(n_12061));
 XOR2x2_ASAP7_75t_SL g21701 (.A(n_19011),
    .B(n_19012),
    .Y(n_13412));
 INVx1_ASAP7_75t_SL g21707 (.A(n_22017),
    .Y(n_13413));
 OAI21x1_ASAP7_75t_SL g21709 (.A1(n_9080),
    .A2(n_13419),
    .B(n_13420),
    .Y(n_11359));
 AND2x2_ASAP7_75t_SL g21710 (.A(n_13418),
    .B(n_9077),
    .Y(n_13419));
 AND2x2_ASAP7_75t_SL g21711 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .Y(n_13418));
 OR2x2_ASAP7_75t_SL g21712 (.A(n_13418),
    .B(n_9077),
    .Y(n_13420));
 XNOR2xp5_ASAP7_75t_SL g21722 (.A(n_21601),
    .B(n_13435),
    .Y(n_13437));
 XNOR2xp5_ASAP7_75t_SL g21725 (.A(n_18969),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_172),
    .Y(n_13435));
 OAI22xp5_ASAP7_75t_SL g21730 (.A1(n_9763),
    .A2(n_13439),
    .B1(n_9762),
    .B2(n_13440),
    .Y(n_13441));
 INVx2_ASAP7_75t_SL g21731 (.A(n_9762),
    .Y(n_13439));
 XNOR2xp5_ASAP7_75t_SL g21733 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_238),
    .B(n_13447),
    .Y(n_13448));
 XNOR2xp5_ASAP7_75t_SL g21734 (.A(n_18737),
    .B(n_14368),
    .Y(n_13447));
 XOR2x2_ASAP7_75t_SL g21739 (.A(n_13450),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_56),
    .Y(n_13451));
 XNOR2xp5_ASAP7_75t_SL g21740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_81),
    .B(n_7269),
    .Y(n_13450));
 AND2x2_ASAP7_75t_SL g21745 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .Y(n_13456));
 NAND2xp5_ASAP7_75t_SL g21747 (.A(n_6025),
    .B(n_13458),
    .Y(n_13459));
 OA21x2_ASAP7_75t_SL g21748 (.A1(n_20758),
    .A2(n_6019),
    .B(n_20759),
    .Y(n_13458));
 XNOR2x1_ASAP7_75t_SL g21751 (.B(n_13465),
    .Y(n_2445),
    .A(n_18790));
 XOR2xp5_ASAP7_75t_SL g21753 (.A(n_13464),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_655),
    .Y(n_13465));
 NAND2xp5_ASAP7_75t_SL g21754 (.A(n_2179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_622),
    .Y(n_13464));
 MAJIxp5_ASAP7_75t_SL g21760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_141),
    .C(n_13475),
    .Y(n_13476));
 XNOR2x1_ASAP7_75t_SL g21761 (.B(n_5930),
    .Y(n_13475),
    .A(n_13474));
 AND2x2_ASAP7_75t_SL g21762 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_742),
    .B(n_2151),
    .Y(n_13474));
 OR2x2_ASAP7_75t_SL g21765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_117),
    .Y(n_13477));
 NOR2xp33_ASAP7_75t_SL g21766 (.A(n_13481),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_258),
    .Y(n_13482));
 NOR2xp33_ASAP7_75t_SL g21767 (.A(n_13480),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_230),
    .Y(n_13481));
 INVxp67_ASAP7_75t_SL g21768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_221),
    .Y(n_13483));
 XNOR2xp5_ASAP7_75t_SL g21777 (.A(n_13495),
    .B(n_13499),
    .Y(n_12411));
 INVx1_ASAP7_75t_SL g21778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_40),
    .Y(n_13498));
 MAJx2_ASAP7_75t_SL g21780 (.A(n_9379),
    .B(n_9375),
    .C(n_14653),
    .Y(n_13502));
 AOI22xp5_ASAP7_75t_SL g21784 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_45),
    .A2(n_13504),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_44),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_76),
    .Y(n_13505));
 AOI22xp5_ASAP7_75t_SL g21788 (.A1(n_13697),
    .A2(n_13784),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_95),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_32),
    .Y(n_13508));
 HB1xp67_ASAP7_75t_SL g21793 (.A(n_14117),
    .Y(n_13519));
 XNOR2xp5_ASAP7_75t_SL g21799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_287),
    .B(n_13523),
    .Y(n_13524));
 NAND2xp5_ASAP7_75t_SL g218 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_96),
    .B(n_20494),
    .Y(n_19913));
 AOI31xp33_ASAP7_75t_SL g21801 (.A1(n_13007),
    .A2(n_13459),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_310),
    .B(n_13521),
    .Y(n_13522));
 XNOR2xp5_ASAP7_75t_SL g21802 (.A(n_20850),
    .B(n_21067),
    .Y(n_13530));
 INVx1_ASAP7_75t_SL g21804 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_10),
    .Y(n_13525));
 XNOR2xp5_ASAP7_75t_SL g21814 (.A(n_13537),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_79),
    .Y(n_13538));
 AND2x2_ASAP7_75t_SL g21815 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .Y(n_13537));
 OAI22x1_ASAP7_75t_SL g21818 (.A1(n_13542),
    .A2(n_13541),
    .B1(n_13543),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_315),
    .Y(n_13544));
 NAND2xp5_ASAP7_75t_SL g21819 (.A(n_22164),
    .B(n_13540),
    .Y(n_13541));
 INVx1_ASAP7_75t_SL g21820 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_226),
    .Y(n_13540));
 INVx2_ASAP7_75t_SL g21821 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_315),
    .Y(n_13542));
 NAND2xp5_ASAP7_75t_SL g21822 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_226),
    .B(n_22164),
    .Y(n_13543));
 HB1xp67_ASAP7_75t_SL g21823 (.A(n_12428),
    .Y(n_13546));
 XNOR2xp5_ASAP7_75t_SL g21824 (.A(n_12424),
    .B(n_16142),
    .Y(n_13551));
 XNOR2xp5_ASAP7_75t_SL g21829 (.A(n_15922),
    .B(n_16140),
    .Y(n_13552));
 OAI21xp5_ASAP7_75t_SL g21842 (.A1(n_13566),
    .A2(n_8196),
    .B(n_8197),
    .Y(n_13567));
 NOR2xp67_ASAP7_75t_SL g21843 (.A(n_20023),
    .B(n_9972),
    .Y(n_13566));
 NAND2xp5_ASAP7_75t_SL g21844 (.A(n_3645),
    .B(n_23290),
    .Y(n_13570));
 OAI21xp5_ASAP7_75t_SL g21846 (.A1(n_20738),
    .A2(n_3644),
    .B(n_23289),
    .Y(n_13571));
 MAJIxp5_ASAP7_75t_SL g21847 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_115),
    .C(n_13574),
    .Y(n_13575));
 HB1xp67_ASAP7_75t_SL g21848 (.A(n_13573),
    .Y(n_13574));
 MAJIxp5_ASAP7_75t_SL g21849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_42),
    .B(n_13572),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_68),
    .Y(n_13573));
 NAND2xp5_ASAP7_75t_SL g21850 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(n_19645),
    .Y(n_13572));
 XOR2xp5_ASAP7_75t_SL g21851 (.A(n_13573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_115),
    .Y(n_13576));
 XOR2x2_ASAP7_75t_SL g21852 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_146),
    .B(n_13572),
    .Y(n_13577));
 INVx1_ASAP7_75t_SL g21856 (.A(n_6968),
    .Y(n_13578));
 MAJIxp5_ASAP7_75t_SL g21858 (.A(n_22232),
    .B(n_6242),
    .C(n_14838),
    .Y(n_13586));
 XNOR2xp5_ASAP7_75t_SL g21861 (.A(n_13393),
    .B(n_13588),
    .Y(n_13589));
 XNOR2x1_ASAP7_75t_SL g21862 (.B(n_26017),
    .Y(n_13588),
    .A(n_19376));
 INVx1_ASAP7_75t_SL g21865 (.A(n_19376),
    .Y(n_13590));
 XNOR2x1_ASAP7_75t_SL g21866 (.B(n_8135),
    .Y(n_13596),
    .A(n_22016));
 INVx1_ASAP7_75t_SL g21870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_99),
    .Y(n_13593));
 MAJIxp5_ASAP7_75t_SL g21871 (.A(n_21971),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_153),
    .C(n_13597),
    .Y(n_13598));
 AO21x2_ASAP7_75t_SL g21874 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_32),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_258),
    .Y(n_13599));
 OAI311xp33_ASAP7_75t_SL g21875 (.A1(n_13600),
    .A2(n_25606),
    .A3(n_19381),
    .B1(n_13608),
    .C1(n_4250),
    .Y(n_13609));
 NAND2xp5_ASAP7_75t_SL g21876 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273),
    .B(n_13606),
    .Y(n_13608));
 XOR2xp5_ASAP7_75t_SL g21878 (.A(n_25607),
    .B(n_13600),
    .Y(n_13612));
 MAJIxp5_ASAP7_75t_SL g21879 (.A(n_13616),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(n_13617));
 XNOR2x2_ASAP7_75t_SL g21880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .B(n_19018),
    .Y(n_13616));
 OAI21xp33_ASAP7_75t_SL g21885 (.A1(n_13621),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_285),
    .B(n_23233),
    .Y(n_13622));
 AOI21x1_ASAP7_75t_SL g21886 (.A1(n_12720),
    .A2(n_21560),
    .B(n_21559),
    .Y(n_13621));
 INVx2_ASAP7_75t_SL g21889 (.A(n_13621),
    .Y(n_13623));
 XOR2xp5_ASAP7_75t_SL g21890 (.A(n_13623),
    .B(n_23232),
    .Y(n_13625));
 NAND2xp5_ASAP7_75t_SL g21892 (.A(n_21560),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_296),
    .Y(n_13627));
 NAND2xp5_ASAP7_75t_SL g21894 (.A(n_13628),
    .B(n_12028),
    .Y(n_13629));
 INVx1_ASAP7_75t_SL g21895 (.A(n_9865),
    .Y(n_13628));
 NAND2x1p5_ASAP7_75t_SL g21897 (.A(n_12018),
    .B(n_12023),
    .Y(n_13631));
 OAI21xp33_ASAP7_75t_L g21898 (.A1(n_15560),
    .A2(n_13631),
    .B(n_12028),
    .Y(n_13634));
 INVx1_ASAP7_75t_L g21900 (.A(n_12028),
    .Y(n_13635));
 NOR2xp67_ASAP7_75t_SL g21901 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_180),
    .B(n_21631),
    .Y(n_13640));
 INVx1_ASAP7_75t_SL g21904 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_106),
    .Y(n_13637));
 NAND2xp5_ASAP7_75t_SL g21905 (.A(n_21631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_180),
    .Y(n_13641));
 MAJIxp5_ASAP7_75t_SL g21908 (.A(n_5890),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_131),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_139),
    .Y(n_13644));
 INVxp33_ASAP7_75t_SRAM g21909 (.A(n_13649),
    .Y(n_13650));
 XNOR2x1_ASAP7_75t_SL g21910 (.B(n_13648),
    .Y(n_13649),
    .A(n_13647));
 XNOR2x1_ASAP7_75t_SL g21911 (.B(n_13646),
    .Y(n_13647),
    .A(n_13645));
 XNOR2xp5_ASAP7_75t_SL g21912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_61),
    .B(n_5804),
    .Y(n_13645));
 MAJIxp5_ASAP7_75t_SL g21913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_107),
    .B(n_6646),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_88),
    .Y(n_13646));
 XNOR2x2_ASAP7_75t_SL g21914 (.A(n_7544),
    .B(n_7548),
    .Y(n_13648));
 OAI21xp5_ASAP7_75t_SL g21915 (.A1(n_13653),
    .A2(n_6658),
    .B(n_13654),
    .Y(n_13655));
 NOR2x1_ASAP7_75t_SL g21916 (.A(n_13649),
    .B(n_13652),
    .Y(n_13653));
 INVxp67_ASAP7_75t_SL g21917 (.A(n_13644),
    .Y(n_13652));
 MAJx2_ASAP7_75t_SL g21918 (.A(n_13648),
    .B(n_13656),
    .C(n_13657),
    .Y(n_13658));
 INVxp67_ASAP7_75t_SL g21919 (.A(n_13646),
    .Y(n_13656));
 HB1xp67_ASAP7_75t_SL g21920 (.A(n_13645),
    .Y(n_13657));
 NOR2xp33_ASAP7_75t_SL g2194 (.A(n_20621),
    .B(n_22012),
    .Y(n_20623));
 AOI21xp33_ASAP7_75t_SL g2195 (.A1(n_23819),
    .A2(n_23818),
    .B(n_17443),
    .Y(n_20637));
 NAND2xp5_ASAP7_75t_SL g21951 (.A(n_13707),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .Y(n_13708));
 NAND2xp5_ASAP7_75t_SL g21953 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .B(n_13707),
    .Y(n_13709));
 NAND2x1_ASAP7_75t_SL g21967 (.A(n_13707),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .Y(n_13723));
 NAND2x1_ASAP7_75t_SL g21968 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .B(n_13707),
    .Y(n_13724));
 NAND2x1_ASAP7_75t_SL g21969 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .B(n_13707),
    .Y(n_13725));
 NAND2x1_ASAP7_75t_SL g21970 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .B(n_3528),
    .Y(n_13726));
 AOI21xp5_ASAP7_75t_SL g2199 (.A1(n_21892),
    .A2(n_22011),
    .B(n_19981),
    .Y(n_20624));
 NAND2xp5_ASAP7_75t_SL g22 (.A(n_21479),
    .B(n_16316),
    .Y(n_21126));
 OAI22xp5_ASAP7_75t_SL g220 (.A1(n_21505),
    .A2(n_20013),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_171),
    .B2(n_20012),
    .Y(n_20248));
 NAND2xp5_ASAP7_75t_SL g2200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .B(n_9974),
    .Y(n_20621));
 NAND2x1p5_ASAP7_75t_SL g22011 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .B(n_16763),
    .Y(n_13767));
 NAND2xp5_ASAP7_75t_SL g22013 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .Y(n_13769));
 NAND2xp5_ASAP7_75t_SL g22014 (.A(n_16763),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .Y(n_13770));
 NAND2x2_ASAP7_75t_SL g22026 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(n_16769),
    .Y(n_13782));
 OR2x2_ASAP7_75t_SL g2205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_373),
    .B(n_17442),
    .Y(n_20633));
 AND2x2_ASAP7_75t_SL g2206 (.A(n_25445),
    .B(n_25981),
    .Y(n_20629));
 AND2x2_ASAP7_75t_SL g2207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_373),
    .B(n_17442),
    .Y(n_20630));
 INVxp67_ASAP7_75t_SL g2208 (.A(n_9974),
    .Y(n_20625));
 MAJx2_ASAP7_75t_SL g22090 (.A(n_14035),
    .B(n_14031),
    .C(n_14033),
    .Y(n_13848));
 INVx1_ASAP7_75t_SL g221 (.A(n_9575),
    .Y(n_12056));
 AOI21x1_ASAP7_75t_SL g22168 (.A1(n_13931),
    .A2(n_13933),
    .B(n_11152),
    .Y(n_13934));
 INVx1_ASAP7_75t_SL g22169 (.A(n_13930),
    .Y(n_13931));
 AOI21x1_ASAP7_75t_SL g22170 (.A1(n_17063),
    .A2(n_13929),
    .B(n_8694),
    .Y(n_13930));
 AO21x1_ASAP7_75t_SL g22171 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_266),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_277),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_264),
    .Y(n_13929));
 NOR2xp67_ASAP7_75t_SL g22172 (.A(n_8902),
    .B(n_13932),
    .Y(n_13933));
 NAND2xp5_ASAP7_75t_SL g22173 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_290),
    .B(n_8690),
    .Y(n_13932));
 NAND2x1p5_ASAP7_75t_SL g22174 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(n_16772),
    .Y(n_13936));
 OAI321xp33_ASAP7_75t_SL g22184 (.A1(n_13082),
    .A2(n_22862),
    .A3(n_13952),
    .B1(n_13952),
    .B2(n_13081),
    .C(n_10791),
    .Y(n_13953));
 NOR2x1_ASAP7_75t_SL g22185 (.A(n_10790),
    .B(n_13951),
    .Y(n_13952));
 OAI21x1_ASAP7_75t_SL g22186 (.A1(n_13945),
    .A2(n_13947),
    .B(n_19019),
    .Y(n_13951));
 NOR2xp33_ASAP7_75t_SL g22187 (.A(n_6463),
    .B(n_6471),
    .Y(n_13945));
 AO21x1_ASAP7_75t_SL g22188 (.A1(n_10758),
    .A2(n_22188),
    .B(n_13946),
    .Y(n_13947));
 NOR2xp33_ASAP7_75t_SL g22189 (.A(n_18863),
    .B(n_26101),
    .Y(n_13946));
 AOI21xp5_ASAP7_75t_SL g22197 (.A1(n_19021),
    .A2(n_13958),
    .B(n_13959),
    .Y(n_13960));
 NAND2xp33_ASAP7_75t_SL g22201 (.A(n_21577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_293),
    .Y(n_13958));
 INVx1_ASAP7_75t_SL g22202 (.A(n_2168),
    .Y(n_13959));
 XNOR2xp5_ASAP7_75t_SL g22205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .B(n_13970),
    .Y(n_13971));
 OAI22xp5_ASAP7_75t_SL g22206 (.A1(n_8505),
    .A2(n_13968),
    .B1(n_13969),
    .B2(n_8507),
    .Y(n_13970));
 XNOR2xp5_ASAP7_75t_SL g22207 (.A(n_26004),
    .B(n_13966),
    .Y(n_13968));
 OAI22xp5_ASAP7_75t_SL g22208 (.A1(n_20833),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_135),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_162),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .Y(n_13966));
 INVx1_ASAP7_75t_SL g22210 (.A(n_13968),
    .Y(n_13969));
 OAI21x1_ASAP7_75t_SL g22211 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_255),
    .A2(n_4151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_254),
    .Y(n_13975));
 NAND2xp5_ASAP7_75t_SL g22212 (.A(n_19890),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_227),
    .Y(n_4151));
 NAND2xp5_ASAP7_75t_SL g22254 (.A(n_13007),
    .B(n_13459),
    .Y(n_14018));
 NAND2xp5_ASAP7_75t_SL g22258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_260),
    .B(n_7543),
    .Y(n_14024));
 NAND2xp5_ASAP7_75t_SL g22259 (.A(n_7539),
    .B(n_5277),
    .Y(n_14025));
 XNOR2xp5_ASAP7_75t_SL g22261 (.A(n_14031),
    .B(n_19022),
    .Y(n_14038));
 AOI21xp5_ASAP7_75t_SL g22263 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_128),
    .Y(n_14031));
 XNOR2x2_ASAP7_75t_SL g22266 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_0),
    .Y(n_14033));
 XNOR2xp5_ASAP7_75t_SL g22267 (.A(n_13843),
    .B(n_13846),
    .Y(n_14035));
 XNOR2x2_ASAP7_75t_SL g22275 (.A(n_14045),
    .B(n_19023),
    .Y(n_14048));
 AND2x2_ASAP7_75t_SL g22276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_0),
    .Y(n_14045));
 XNOR2x2_ASAP7_75t_SL g22280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_3),
    .B(n_14049),
    .Y(n_14050));
 INVxp67_ASAP7_75t_SL g22281 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_73),
    .Y(n_14049));
 INVxp67_ASAP7_75t_SL g22289 (.A(n_22465),
    .Y(n_14061));
 INVxp67_ASAP7_75t_SL g22291 (.A(n_19270),
    .Y(n_14067));
 AO22x2_ASAP7_75t_SL g22293 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_149),
    .A2(n_14062),
    .B1(n_6579),
    .B2(n_14063),
    .Y(n_14064));
 INVx1_ASAP7_75t_SL g22294 (.A(n_6579),
    .Y(n_14062));
 INVx1_ASAP7_75t_SL g22295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_149),
    .Y(n_14063));
 XNOR2xp5_ASAP7_75t_SL g223 (.A(n_20785),
    .B(n_22960),
    .Y(n_20786));
 NOR2xp67_ASAP7_75t_SL g22315 (.A(n_19339),
    .B(n_14088),
    .Y(n_14089));
 XNOR2xp5_ASAP7_75t_SL g22316 (.A(n_21580),
    .B(n_14087),
    .Y(n_14088));
 XNOR2xp5_ASAP7_75t_SL g22317 (.A(n_20496),
    .B(n_5339),
    .Y(n_14087));
 NAND2xp5_ASAP7_75t_SL g22318 (.A(n_14088),
    .B(n_19339),
    .Y(n_14090));
 AOI21xp5_ASAP7_75t_SL g22319 (.A1(n_14087),
    .A2(n_21581),
    .B(n_21582),
    .Y(n_14091));
 NAND2xp5_ASAP7_75t_SL g22322 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .Y(n_14092));
 OAI22xp5_ASAP7_75t_SL g22328 (.A1(n_18915),
    .A2(n_14101),
    .B1(n_14102),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_222),
    .Y(n_14103));
 MAJIxp5_ASAP7_75t_SL g22329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_171),
    .B(n_14100),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_1),
    .Y(n_14101));
 MAJx2_ASAP7_75t_SL g22330 (.A(n_7234),
    .B(n_7233),
    .C(n_7231),
    .Y(n_14100));
 MAJx2_ASAP7_75t_SL g22332 (.A(n_13401),
    .B(n_14102),
    .C(n_8747),
    .Y(n_14105));
 INVx2_ASAP7_75t_SL g22333 (.A(n_14101),
    .Y(n_14102));
 XNOR2xp5_ASAP7_75t_SL g22334 (.A(n_14100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_11),
    .Y(n_14106));
 OAI21xp5_ASAP7_75t_SL g22335 (.A1(n_14108),
    .A2(n_6298),
    .B(n_14109),
    .Y(n_14110));
 NOR2xp33_ASAP7_75t_SL g22336 (.A(n_20327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_14108));
 NAND2xp5_ASAP7_75t_SL g22338 (.A(n_20327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_14109));
 OAI21xp5_ASAP7_75t_SL g22339 (.A1(n_17416),
    .A2(n_14108),
    .B(n_14109),
    .Y(n_14111));
 OAI22xp5_ASAP7_75t_SL g22343 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_293),
    .A2(n_14120),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_294),
    .B2(n_22541),
    .Y(n_14121));
 INVx2_ASAP7_75t_SL g22344 (.A(n_22541),
    .Y(n_14120));
 MAJIxp5_ASAP7_75t_SL g22346 (.A(n_26264),
    .B(n_14123),
    .C(n_14124),
    .Y(n_14125));
 HB1xp67_ASAP7_75t_SL g22347 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_294),
    .Y(n_14123));
 HB1xp67_ASAP7_75t_SL g22348 (.A(n_22541),
    .Y(n_14124));
 AND2x2_ASAP7_75t_SL g22355 (.A(n_25302),
    .B(n_21996),
    .Y(n_14135));
 NOR2xp67_ASAP7_75t_SL g22358 (.A(n_25302),
    .B(n_21996),
    .Y(n_14136));
 MAJIxp5_ASAP7_75t_SL g22359 (.A(n_21621),
    .B(n_5959),
    .C(n_21994),
    .Y(n_14137));
 OAI22xp5_ASAP7_75t_SL g22360 (.A1(n_14140),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_293),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_294),
    .B2(n_23125),
    .Y(n_14141));
 INVx2_ASAP7_75t_SL g22361 (.A(n_23125),
    .Y(n_14140));
 INVx1_ASAP7_75t_SL g22368 (.A(n_20234),
    .Y(n_14143));
 NOR2x1_ASAP7_75t_SL g22369 (.A(n_20863),
    .B(n_20867),
    .Y(n_14147));
 NOR2x1_ASAP7_75t_SL g22370 (.A(n_18791),
    .B(n_24213),
    .Y(n_14151));
 NAND2xp5_ASAP7_75t_SL g22374 (.A(n_18791),
    .B(n_24213),
    .Y(n_14152));
 XNOR2xp5_ASAP7_75t_SL g22375 (.A(n_18798),
    .B(n_19197),
    .Y(n_10012));
 NAND2xp5_ASAP7_75t_SL g22377 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .Y(n_14153));
 MAJIxp5_ASAP7_75t_SL g22380 (.A(n_14153),
    .B(n_15332),
    .C(n_14158),
    .Y(n_14159));
 AOI21xp5_ASAP7_75t_SL g22382 (.A1(n_14708),
    .A2(n_19953),
    .B(n_19952),
    .Y(n_14162));
 NAND2xp33_ASAP7_75t_L g22442 (.A(n_14241),
    .B(n_11413),
    .Y(n_14242));
 XOR2x2_ASAP7_75t_SL g22443 (.A(n_19027),
    .B(n_14238),
    .Y(n_14241));
 NOR2xp33_ASAP7_75t_SL g22446 (.A(n_11413),
    .B(n_14241),
    .Y(n_14243));
 XNOR2x1_ASAP7_75t_SL g22447 (.B(n_14241),
    .Y(n_14244),
    .A(n_11413));
 XNOR2xp5_ASAP7_75t_SL g225 (.A(n_2588),
    .B(n_14121),
    .Y(n_14122));
 MAJIxp5_ASAP7_75t_SL g22501 (.A(n_9009),
    .B(n_14298),
    .C(n_12988),
    .Y(n_14299));
 MAJIxp5_ASAP7_75t_SL g22502 (.A(n_21046),
    .B(n_21048),
    .C(n_21049),
    .Y(n_14298));
 XNOR2xp5_ASAP7_75t_SL g22503 (.A(n_12988),
    .B(n_14300),
    .Y(n_14301));
 NAND2xp5_ASAP7_75t_SL g22529 (.A(n_18577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_280),
    .Y(n_14327));
 NAND2xp5_ASAP7_75t_SL g22530 (.A(n_14329),
    .B(n_12567),
    .Y(n_14330));
 NOR2xp33_ASAP7_75t_SL g22531 (.A(n_5799),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_280),
    .Y(n_14329));
 OAI21xp5_ASAP7_75t_SL g22533 (.A1(n_14333),
    .A2(n_14334),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_270),
    .Y(n_14335));
 NAND2xp5_ASAP7_75t_SL g22534 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_271),
    .B(n_6392),
    .Y(n_14333));
 INVxp67_ASAP7_75t_SL g22536 (.A(n_6397),
    .Y(n_14334));
 NAND2x1_ASAP7_75t_SL g22537 (.A(n_6392),
    .B(n_6397),
    .Y(n_14336));
 MAJx2_ASAP7_75t_SL g22540 (.A(n_7819),
    .B(n_14339),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_709),
    .Y(n_14340));
 AND2x4_ASAP7_75t_SL g22541 (.A(n_2173),
    .B(n_12101),
    .Y(n_14339));
 XNOR2x1_ASAP7_75t_SL g22543 (.B(n_26174),
    .Y(n_14344),
    .A(n_6361));
 NAND2xp5_ASAP7_75t_SL g22552 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .Y(n_14353));
 OAI22xp5_ASAP7_75t_SL g22554 (.A1(n_13596),
    .A2(n_8141),
    .B1(n_8137),
    .B2(n_8140),
    .Y(n_14354));
 XNOR2xp5_ASAP7_75t_SL g22562 (.A(n_14364),
    .B(n_14367),
    .Y(n_14368));
 INVx1_ASAP7_75t_SL g22563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_150),
    .Y(n_14364));
 AOI22xp5_ASAP7_75t_SL g22564 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_145),
    .A2(n_7263),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_146),
    .B2(n_19144),
    .Y(n_14367));
 NOR2x1_ASAP7_75t_SL g22574 (.A(n_14928),
    .B(n_19235),
    .Y(n_14382));
 AOI22x1_ASAP7_75t_SL g22579 (.A1(n_14384),
    .A2(n_23493),
    .B1(n_14383),
    .B2(n_12956),
    .Y(n_14386));
 INVx2_ASAP7_75t_L g22580 (.A(n_14383),
    .Y(n_14384));
 XNOR2x2_ASAP7_75t_SL g22581 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_63),
    .B(n_21930),
    .Y(n_14383));
 XNOR2xp5_ASAP7_75t_SL g22584 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_192),
    .B(n_19029),
    .Y(n_14394));
 NOR2xp33_ASAP7_75t_SL g226 (.A(n_20776),
    .B(n_20777),
    .Y(n_20778));
 MAJx2_ASAP7_75t_SL g22602 (.A(n_14407),
    .B(n_14408),
    .C(n_14414),
    .Y(n_14415));
 INVxp67_ASAP7_75t_SL g22603 (.A(n_8596),
    .Y(n_14407));
 INVx1_ASAP7_75t_SL g22604 (.A(n_8594),
    .Y(n_14408));
 MAJIxp5_ASAP7_75t_SL g22605 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_202),
    .B(n_14411),
    .C(n_14413),
    .Y(n_14414));
 HB1xp67_ASAP7_75t_SL g22609 (.A(n_14412),
    .Y(n_14413));
 XNOR2xp5_ASAP7_75t_SL g22610 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_132),
    .Y(n_14412));
 XNOR2xp5_ASAP7_75t_SL g22611 (.A(n_14416),
    .B(n_13333),
    .Y(n_14417));
 INVxp67_ASAP7_75t_SL g22612 (.A(n_14414),
    .Y(n_14416));
 XNOR2xp5_ASAP7_75t_SL g22613 (.A(n_14411),
    .B(n_14412),
    .Y(n_14418));
 OAI21xp5_ASAP7_75t_SL g22620 (.A1(n_15091),
    .A2(n_8787),
    .B(n_15087),
    .Y(n_14427));
 NOR2xp67_ASAP7_75t_SL g22622 (.A(n_11419),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_288),
    .Y(n_14425));
 OAI21xp5_ASAP7_75t_SL g22623 (.A1(n_11304),
    .A2(n_6265),
    .B(n_14429),
    .Y(n_14430));
 NAND2xp5_ASAP7_75t_SL g22626 (.A(n_11302),
    .B(n_14429),
    .Y(n_14431));
 INVxp67_ASAP7_75t_SRAM g22628 (.A(n_14706),
    .Y(n_14434));
 XNOR2xp5_ASAP7_75t_SL g22631 (.A(n_6774),
    .B(n_14706),
    .Y(n_14436));
 INVx1_ASAP7_75t_SL g22632 (.A(n_14437),
    .Y(n_14438));
 MAJx2_ASAP7_75t_SL g22633 (.A(n_9359),
    .B(n_13477),
    .C(n_10281),
    .Y(n_14437));
 INVx1_ASAP7_75t_SL g22634 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_10),
    .Y(n_14440));
 INVx1_ASAP7_75t_SL g22635 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_171),
    .Y(n_14441));
 XNOR2xp5_ASAP7_75t_SL g22641 (.A(n_14451),
    .B(n_12079),
    .Y(n_14452));
 MAJx2_ASAP7_75t_SL g22642 (.A(n_6452),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .Y(n_14451));
 HB1xp67_ASAP7_75t_SL g22644 (.A(n_14451),
    .Y(n_14454));
 XNOR2xp5_ASAP7_75t_SL g22647 (.A(n_14456),
    .B(n_12631),
    .Y(n_14457));
 XNOR2xp5_ASAP7_75t_SL g22648 (.A(n_8612),
    .B(n_12634),
    .Y(n_14456));
 MAJIxp5_ASAP7_75t_SL g227 (.A(n_12069),
    .B(n_6372),
    .C(n_18700),
    .Y(n_6373));
 AND2x2_ASAP7_75t_SL g22791 (.A(n_12781),
    .B(n_10106),
    .Y(n_14643));
 XNOR2x1_ASAP7_75t_SL g22792 (.B(n_13772),
    .Y(n_14645),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_67));
 NAND2xp5_ASAP7_75t_SL g22793 (.A(n_13772),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_67),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_111));
 MAJIxp5_ASAP7_75t_SL g22799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_81),
    .B(n_14652),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_20),
    .Y(n_14653));
 AND2x2_ASAP7_75t_SL g228 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_193),
    .Y(n_20773));
 NAND2x1_ASAP7_75t_SL g22800 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(n_13707),
    .Y(n_14652));
 XNOR2xp5_ASAP7_75t_SL g22810 (.A(n_18793),
    .B(n_14664),
    .Y(n_2442));
 XNOR2x1_ASAP7_75t_SL g22812 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_655),
    .Y(n_14664),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_623));
 XNOR2x2_ASAP7_75t_SL g22813 (.A(n_19032),
    .B(n_14669),
    .Y(n_11509));
 INVxp67_ASAP7_75t_SL g22817 (.A(n_22620),
    .Y(n_14669));
 NAND2xp67_ASAP7_75t_SL g22820 (.A(n_14674),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .Y(n_14675));
 INVx2_ASAP7_75t_SL g22829 (.A(n_14683),
    .Y(n_14684));
 XNOR2x1_ASAP7_75t_SL g22830 (.B(n_11793),
    .Y(n_14683),
    .A(n_4957));
 NOR2x1_ASAP7_75t_SL g22832 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_250),
    .B(n_14687),
    .Y(n_14688));
 XNOR2xp5_ASAP7_75t_L g22833 (.A(n_18794),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_146),
    .Y(n_14687));
 NOR2x1p5_ASAP7_75t_SL g22836 (.A(n_6218),
    .B(n_22955),
    .Y(n_14689));
 NAND2xp5_ASAP7_75t_SL g22843 (.A(n_10953),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_269),
    .Y(n_14695));
 MAJIxp5_ASAP7_75t_SL g22845 (.A(n_19253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_172),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_186),
    .Y(n_14698));
 XOR2xp5_ASAP7_75t_SL g22847 (.A(n_14701),
    .B(n_9669),
    .Y(n_14702));
 XNOR2x1_ASAP7_75t_SL g22848 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_20),
    .Y(n_14701),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_709));
 XNOR2xp5_ASAP7_75t_SL g22849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_61),
    .B(n_14705),
    .Y(n_14706));
 OAI22xp33_ASAP7_75t_SL g22850 (.A1(n_14703),
    .A2(n_13718),
    .B1(n_14704),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_95),
    .Y(n_14705));
 NAND2x1_ASAP7_75t_SL g22851 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_11770),
    .Y(n_14703));
 INVx1_ASAP7_75t_SL g22852 (.A(n_14703),
    .Y(n_14704));
 XNOR2xp5_ASAP7_75t_SL g22853 (.A(n_19956),
    .B(n_14708),
    .Y(n_14709));
 XNOR2xp5_ASAP7_75t_SL g22854 (.A(n_14437),
    .B(n_18849),
    .Y(n_14708));
 XOR2xp5_ASAP7_75t_SL g22858 (.A(n_18702),
    .B(n_19041),
    .Y(n_14713));
 XNOR2x1_ASAP7_75t_SL g22861 (.B(n_14717),
    .Y(n_14718),
    .A(n_14716));
 XNOR2xp5_ASAP7_75t_SL g22862 (.A(n_15584),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_109),
    .Y(n_14716));
 HB1xp67_ASAP7_75t_SL g22864 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_65),
    .Y(n_14717));
 XOR2xp5_ASAP7_75t_SL g22866 (.A(n_14722),
    .B(n_6186),
    .Y(n_14723));
 XNOR2xp5_ASAP7_75t_SL g22867 (.A(n_14721),
    .B(n_21513),
    .Y(n_14722));
 MAJx2_ASAP7_75t_SL g22868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_5),
    .B(n_14720),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_32),
    .Y(n_14721));
 NOR2xp33_ASAP7_75t_SL g22869 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_80),
    .Y(n_14720));
 NOR2xp33_ASAP7_75t_SL g22870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_80),
    .Y(n_14724));
 AND2x2_ASAP7_75t_SL g22874 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .Y(n_14725));
 XNOR2xp5_ASAP7_75t_SL g22875 (.A(n_14729),
    .B(n_14735),
    .Y(n_14736));
 OA21x2_ASAP7_75t_SL g22876 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_167),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_189),
    .Y(n_14729));
 OAI21xp5_ASAP7_75t_SL g22877 (.A1(n_14731),
    .A2(n_14732),
    .B(n_14734),
    .Y(n_14735));
 INVxp67_ASAP7_75t_SL g22878 (.A(n_14730),
    .Y(n_14731));
 NOR2xp33_ASAP7_75t_SL g22879 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_246),
    .Y(n_14730));
 OA21x2_ASAP7_75t_SL g22880 (.A1(n_16663),
    .A2(n_8290),
    .B(n_15188),
    .Y(n_14732));
 OAI21xp5_ASAP7_75t_SL g22881 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_244),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_236),
    .Y(n_14733));
 OAI21xp5_ASAP7_75t_SL g22884 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_128),
    .A2(n_14739),
    .B(n_14740),
    .Y(n_14741));
 OAI21xp5_ASAP7_75t_SL g22885 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_141),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_5),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_103),
    .Y(n_14740));
 INVx1_ASAP7_75t_SL g22886 (.A(n_14746),
    .Y(n_7296));
 XNOR2x1_ASAP7_75t_SL g22895 (.B(n_14762),
    .Y(n_14763),
    .A(n_14760));
 XNOR2x1_ASAP7_75t_SL g22896 (.B(n_14759),
    .Y(n_14760),
    .A(n_14758));
 AND2x2_ASAP7_75t_SL g22897 (.A(n_20825),
    .B(n_20983),
    .Y(n_14758));
 AND2x4_ASAP7_75t_SL g22898 (.A(n_2161),
    .B(n_19584),
    .Y(n_14759));
 INVx2_ASAP7_75t_L g22899 (.A(n_14761),
    .Y(n_14762));
 MAJIxp5_ASAP7_75t_SL g229 (.A(n_26249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .C(n_6253),
    .Y(n_6254));
 AND2x2_ASAP7_75t_SL g22900 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_770),
    .Y(n_14761));
 AOI31xp33_ASAP7_75t_SL g22901 (.A1(n_14764),
    .A2(n_14769),
    .A3(n_14770),
    .B(n_14771),
    .Y(n_14772));
 NAND2xp5_ASAP7_75t_SL g22902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .Y(n_14764));
 NAND2xp5_ASAP7_75t_SL g22903 (.A(n_19034),
    .B(n_14768),
    .Y(n_14769));
 MAJIxp5_ASAP7_75t_SL g22907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_325),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .Y(n_14768));
 NAND2xp5_ASAP7_75t_SL g22908 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(n_14770));
 NOR2xp67_ASAP7_75t_SL g22909 (.A(n_14768),
    .B(n_19034),
    .Y(n_14771));
 HB1xp67_ASAP7_75t_SL g22910 (.A(n_14772),
    .Y(n_14773));
 OAI21xp5_ASAP7_75t_SL g22911 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(n_14774));
 MAJIxp5_ASAP7_75t_SL g22918 (.A(n_14781),
    .B(n_14783),
    .C(n_14784),
    .Y(n_14785));
 AND2x2_ASAP7_75t_SL g22919 (.A(n_14987),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .Y(n_14781));
 AND2x2_ASAP7_75t_SL g22920 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(n_19645),
    .Y(n_14783));
 NAND2x2_ASAP7_75t_SL g22922 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .Y(n_14784));
 NAND2xp5_ASAP7_75t_SL g22923 (.A(n_19645),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .Y(n_14786));
 XNOR2x2_ASAP7_75t_SL g22926 (.A(n_14788),
    .B(n_3235),
    .Y(n_14791));
 NOR2x1_ASAP7_75t_SL g22927 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_57),
    .Y(n_14788));
 OAI22xp5_ASAP7_75t_SL g22928 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_51),
    .Y(n_3235));
 OAI21xp5_ASAP7_75t_SL g22934 (.A1(n_14798),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_285),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_292),
    .Y(n_14799));
 AOI21x1_ASAP7_75t_SL g22935 (.A1(n_14809),
    .A2(n_23776),
    .B(n_8826),
    .Y(n_14798));
 OAI22xp33_ASAP7_75t_SL g22939 (.A1(n_14800),
    .A2(n_14803),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_304),
    .B2(n_14798),
    .Y(n_14804));
 INVxp67_ASAP7_75t_SL g22940 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_304),
    .Y(n_14803));
 XNOR2xp5_ASAP7_75t_SL g22941 (.A(n_10711),
    .B(n_14805),
    .Y(n_14806));
 HB1xp67_ASAP7_75t_SL g22942 (.A(n_14809),
    .Y(n_14805));
 AO21x1_ASAP7_75t_SL g22943 (.A1(n_8821),
    .A2(n_14808),
    .B(n_8823),
    .Y(n_14809));
 OAI21xp5_ASAP7_75t_SL g22944 (.A1(n_14807),
    .A2(n_8666),
    .B(n_10697),
    .Y(n_14808));
 NOR2xp67_ASAP7_75t_SL g22945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_207),
    .B(n_8657),
    .Y(n_14807));
 OAI22x1_ASAP7_75t_SL g22946 (.A1(n_14810),
    .A2(n_12991),
    .B1(n_14811),
    .B2(n_12993),
    .Y(n_14812));
 NAND2xp5_ASAP7_75t_SL g22948 (.A(n_10697),
    .B(n_14813),
    .Y(n_14814));
 INVxp67_ASAP7_75t_SRAM g22949 (.A(n_14807),
    .Y(n_14813));
 XOR2xp5_ASAP7_75t_SL g22950 (.A(n_7162),
    .B(n_19199),
    .Y(n_14819));
 NAND2xp5_ASAP7_75t_SL g22952 (.A(n_3706),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .Y(n_14815));
 INVxp67_ASAP7_75t_SRAM g22954 (.A(n_14815),
    .Y(n_14820));
 OAI22xp5_ASAP7_75t_SL g22956 (.A1(n_14822),
    .A2(n_14823),
    .B1(n_14824),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_43),
    .Y(n_14825));
 NAND2xp5_ASAP7_75t_SL g22957 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .Y(n_14822));
 INVx1_ASAP7_75t_SL g22958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_43),
    .Y(n_14823));
 INVx1_ASAP7_75t_SL g22959 (.A(n_14822),
    .Y(n_14824));
 MAJIxp5_ASAP7_75t_SL g22960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_152),
    .B(n_14824),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_43),
    .Y(n_14826));
 NAND2xp5_ASAP7_75t_SL g22961 (.A(n_22090),
    .B(n_20335),
    .Y(n_14835));
 XOR2x2_ASAP7_75t_SL g22963 (.A(n_14829),
    .B(n_14831),
    .Y(n_14832));
 OAI22xp5_ASAP7_75t_SL g22964 (.A1(n_14827),
    .A2(n_6156),
    .B1(n_6157),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_13),
    .Y(n_14829));
 INVx1_ASAP7_75t_SL g22965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_13),
    .Y(n_14827));
 MAJIxp5_ASAP7_75t_SL g22967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_133),
    .B(n_6243),
    .C(n_20329),
    .Y(n_14831));
 NOR2xp67_ASAP7_75t_SL g22970 (.A(n_20335),
    .B(n_22090),
    .Y(n_14836));
 MAJIxp5_ASAP7_75t_SL g22971 (.A(n_14832),
    .B(n_23431),
    .C(n_6128),
    .Y(n_14837));
 MAJIxp5_ASAP7_75t_SL g22972 (.A(n_6157),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_13),
    .C(n_14831),
    .Y(n_14838));
 MAJIxp5_ASAP7_75t_SL g22990 (.A(n_18940),
    .B(n_14878),
    .C(n_16352),
    .Y(n_14864));
 MAJIxp5_ASAP7_75t_SL g22995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_49),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_67),
    .Y(n_14857));
 AND2x2_ASAP7_75t_SL g23 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(n_13231),
    .Y(n_19607));
 HB1xp67_ASAP7_75t_SL g230 (.A(n_15626),
    .Y(n_6253));
 MAJIxp5_ASAP7_75t_SL g23000 (.A(n_20478),
    .B(n_9419),
    .C(n_14867),
    .Y(n_14868));
 INVx1_ASAP7_75t_SL g23001 (.A(n_16347),
    .Y(n_14867));
 OAI22xp5_ASAP7_75t_SL g23003 (.A1(n_17998),
    .A2(n_9279),
    .B1(n_17997),
    .B2(n_26137),
    .Y(n_14877));
 NAND2xp5_ASAP7_75t_SL g23005 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_15192),
    .Y(n_14871));
 XOR2xp5_ASAP7_75t_SL g23006 (.A(n_14872),
    .B(n_14873),
    .Y(n_14874));
 NAND2xp5_ASAP7_75t_SL g23007 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(n_18031),
    .Y(n_14872));
 AND2x2_ASAP7_75t_SL g23008 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .B(n_3218),
    .Y(n_14873));
 AO21x1_ASAP7_75t_SL g23010 (.A1(n_17998),
    .A2(n_21459),
    .B(n_21458),
    .Y(n_14878));
 MAJIxp5_ASAP7_75t_SL g23011 (.A(n_14871),
    .B(n_14873),
    .C(n_14872),
    .Y(n_9419));
 XNOR2xp5_ASAP7_75t_SL g23014 (.A(n_14881),
    .B(n_15453),
    .Y(n_14883));
 INVxp67_ASAP7_75t_SL g23017 (.A(n_15453),
    .Y(n_14887));
 NOR2xp33_ASAP7_75t_SL g23018 (.A(n_17870),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_425),
    .Y(n_14891));
 AND2x2_ASAP7_75t_SL g23022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_462),
    .B(n_3942),
    .Y(n_14894));
 INVxp67_ASAP7_75t_SL g23023 (.A(n_2850),
    .Y(n_14896));
 MAJIxp5_ASAP7_75t_SL g23024 (.A(n_14906),
    .B(n_6774),
    .C(n_14434),
    .Y(n_14907));
 XNOR2x1_ASAP7_75t_SL g23025 (.B(n_14905),
    .Y(n_14906),
    .A(n_18836));
 XNOR2xp5_ASAP7_75t_SL g23027 (.A(n_14902),
    .B(n_14904),
    .Y(n_14905));
 NAND2xp5_ASAP7_75t_SL g23028 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_3374),
    .Y(n_14902));
 INVx2_ASAP7_75t_SL g23029 (.A(n_14903),
    .Y(n_14904));
 NAND2xp5_ASAP7_75t_SL g23030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_121),
    .Y(n_14903));
 XOR2xp5_ASAP7_75t_SL g23031 (.A(n_14436),
    .B(n_14906),
    .Y(n_14908));
 OAI21x1_ASAP7_75t_SL g23032 (.A1(n_14909),
    .A2(n_18836),
    .B(n_14911),
    .Y(n_14912));
 AND2x2_ASAP7_75t_SL g23033 (.A(n_14903),
    .B(n_14902),
    .Y(n_14909));
 NAND2xp5_ASAP7_75t_SL g23034 (.A(n_14910),
    .B(n_14904),
    .Y(n_14911));
 NAND2xp5_ASAP7_75t_SL g23036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_270),
    .B(n_14920),
    .Y(n_14921));
 XNOR2xp5_ASAP7_75t_SL g23037 (.A(n_14914),
    .B(n_19037),
    .Y(n_14920));
 MAJx2_ASAP7_75t_SL g23038 (.A(n_18942),
    .B(n_3088),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_182),
    .Y(n_14914));
 MAJIxp5_ASAP7_75t_SL g23041 (.A(n_7863),
    .B(n_7862),
    .C(n_10100),
    .Y(n_14915));
 NOR2x1_ASAP7_75t_SL g23046 (.A(n_14920),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_270),
    .Y(n_14925));
 MAJIxp5_ASAP7_75t_SL g23047 (.A(n_14926),
    .B(n_14915),
    .C(n_14927),
    .Y(n_14928));
 INVx1_ASAP7_75t_SL g23048 (.A(n_14914),
    .Y(n_14926));
 HB1xp67_ASAP7_75t_SL g23049 (.A(n_19038),
    .Y(n_14927));
 NAND2xp5_ASAP7_75t_SL g23050 (.A(n_14940),
    .B(n_9950),
    .Y(n_14941));
 OAI21xp5_ASAP7_75t_SL g23051 (.A1(n_14929),
    .A2(n_14937),
    .B(n_14939),
    .Y(n_14940));
 AOI21xp5_ASAP7_75t_SL g23052 (.A1(n_14932),
    .A2(n_14934),
    .B(n_14936),
    .Y(n_14937));
 NAND2xp5_ASAP7_75t_SL g23053 (.A(n_18795),
    .B(n_14931),
    .Y(n_14932));
 NAND2xp5_ASAP7_75t_SL g23054 (.A(n_14933),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_201),
    .Y(n_14934));
 INVx1_ASAP7_75t_SL g23055 (.A(n_14935),
    .Y(n_14936));
 MAJIxp5_ASAP7_75t_SL g23056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_117),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_128),
    .Y(n_14935));
 NAND2xp5_ASAP7_75t_SL g23057 (.A(n_14936),
    .B(n_14938),
    .Y(n_14939));
 AOI22xp5_ASAP7_75t_SL g23058 (.A1(n_18795),
    .A2(n_14931),
    .B1(n_14933),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_201),
    .Y(n_14938));
 AND2x2_ASAP7_75t_SL g23059 (.A(n_14943),
    .B(n_10446),
    .Y(n_14944));
 NAND2xp5_ASAP7_75t_SL g23060 (.A(n_9950),
    .B(n_14940),
    .Y(n_14943));
 XNOR2xp5_ASAP7_75t_SL g23062 (.A(n_10443),
    .B(n_14945),
    .Y(n_14946));
 INVxp67_ASAP7_75t_SRAM g23063 (.A(n_14940),
    .Y(n_14945));
 XNOR2xp5_ASAP7_75t_SL g23064 (.A(n_14948),
    .B(n_14949),
    .Y(n_14950));
 XNOR2xp5_ASAP7_75t_SL g23065 (.A(n_14935),
    .B(n_14947),
    .Y(n_14948));
 INVxp67_ASAP7_75t_SL g23067 (.A(n_14929),
    .Y(n_14949));
 OAI21xp5_ASAP7_75t_SL g231 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_133),
    .A2(n_9405),
    .B(n_9406),
    .Y(n_9407));
 MAJIxp5_ASAP7_75t_SL g23141 (.A(n_11423),
    .B(n_4107),
    .C(n_5649),
    .Y(n_15084));
 AOI21xp5_ASAP7_75t_SL g23143 (.A1(n_14425),
    .A2(n_15086),
    .B(n_12287),
    .Y(n_15087));
 NAND2xp5_ASAP7_75t_SL g23144 (.A(n_15084),
    .B(n_15085),
    .Y(n_15086));
 AND2x2_ASAP7_75t_SL g23146 (.A(n_15086),
    .B(n_6266),
    .Y(n_15090));
 NAND2xp5_ASAP7_75t_SL g23148 (.A(n_15086),
    .B(n_11298),
    .Y(n_15091));
 MAJx2_ASAP7_75t_SL g23152 (.A(n_14718),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_33),
    .C(n_15096),
    .Y(n_15097));
 XNOR2x1_ASAP7_75t_SL g232 (.B(n_9074),
    .Y(n_9408),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_13));
 NAND2xp5_ASAP7_75t_SL g23206 (.A(n_6833),
    .B(n_10513),
    .Y(n_15153));
 AND2x2_ASAP7_75t_SL g23212 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .Y(n_15156));
 OR2x2_ASAP7_75t_SL g23214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_58),
    .Y(n_15158));
 NAND2xp5_ASAP7_75t_SL g23218 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .Y(n_15163));
 XOR2xp5_ASAP7_75t_SL g23293 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_96),
    .Y(n_15289));
 MAJIxp5_ASAP7_75t_SL g233 (.A(n_6853),
    .B(n_19314),
    .C(n_26008),
    .Y(n_19316));
 INVx1_ASAP7_75t_SL g234 (.A(n_18858),
    .Y(n_6128));
 AND2x2_ASAP7_75t_SL g23420 (.A(n_10778),
    .B(n_13456),
    .Y(n_15449));
 MAJx2_ASAP7_75t_SL g23423 (.A(n_15567),
    .B(n_18664),
    .C(n_4793),
    .Y(n_15453));
 XOR2xp5_ASAP7_75t_SL g23426 (.A(n_12962),
    .B(n_19002),
    .Y(n_15456));
 XNOR2x1_ASAP7_75t_SL g23427 (.B(n_19002),
    .Y(n_15457),
    .A(n_12962));
 OA21x2_ASAP7_75t_SL g235 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_298),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_301),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_211),
    .Y(n_10592));
 NAND2xp33_ASAP7_75t_SL g23517 (.A(n_24102),
    .B(n_19970),
    .Y(n_15549));
 AND2x2_ASAP7_75t_SL g23519 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(n_16769),
    .Y(n_15551));
 NAND2xp5_ASAP7_75t_SL g23520 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(n_16772),
    .Y(n_15552));
 XNOR2xp5_ASAP7_75t_SL g23521 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_42),
    .B(n_22994),
    .Y(n_15553));
 NOR2x1p5_ASAP7_75t_SL g23528 (.A(n_15560),
    .B(n_13631),
    .Y(n_15561));
 AND2x2_ASAP7_75t_SL g23529 (.A(n_12013),
    .B(n_15559),
    .Y(n_15560));
 NOR2x1_ASAP7_75t_SL g23530 (.A(n_17560),
    .B(n_10348),
    .Y(n_15559));
 XNOR2x2_ASAP7_75t_SL g23532 (.A(n_15568),
    .B(n_15569),
    .Y(n_15570));
 XNOR2xp5_ASAP7_75t_SL g23533 (.A(n_18664),
    .B(n_15567),
    .Y(n_15568));
 XOR2xp5_ASAP7_75t_SL g23534 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_48),
    .B(n_18953),
    .Y(n_15567));
 INVxp67_ASAP7_75t_SL g23538 (.A(n_4793),
    .Y(n_15569));
 XOR2xp5_ASAP7_75t_SL g23540 (.A(n_15579),
    .B(n_22802),
    .Y(n_15581));
 OAI21xp5_ASAP7_75t_SL g23542 (.A1(n_15575),
    .A2(n_7638),
    .B(n_15578),
    .Y(n_15579));
 NAND2xp5_ASAP7_75t_SL g23543 (.A(n_15573),
    .B(n_15574),
    .Y(n_15575));
 INVxp67_ASAP7_75t_SL g23544 (.A(n_15572),
    .Y(n_15573));
 NAND2xp5_ASAP7_75t_SL g23545 (.A(n_12748),
    .B(n_15571),
    .Y(n_15572));
 INVxp67_ASAP7_75t_SL g23546 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_217),
    .Y(n_15571));
 INVx1_ASAP7_75t_SL g23547 (.A(n_7644),
    .Y(n_15574));
 AOI31xp33_ASAP7_75t_SL g23548 (.A1(n_15574),
    .A2(n_15576),
    .A3(n_15573),
    .B(n_15577),
    .Y(n_15578));
 INVxp67_ASAP7_75t_SL g23549 (.A(n_7637),
    .Y(n_15576));
 NOR2xp33_ASAP7_75t_SL g23550 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_213),
    .B(n_15572),
    .Y(n_15577));
 NAND2x1p5_ASAP7_75t_SL g23551 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .B(n_24402),
    .Y(n_15584));
 NAND2x1_ASAP7_75t_SL g23561 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .Y(n_6932));
 XOR2x1_ASAP7_75t_SL g23594 (.A(n_8770),
    .Y(n_15626),
    .B(n_24202));
 INVxp67_ASAP7_75t_SL g236 (.A(n_9313),
    .Y(n_19314));
 XNOR2xp5_ASAP7_75t_SL g23608 (.A(n_15641),
    .B(n_19036),
    .Y(n_15645));
 INVx1_ASAP7_75t_SL g23609 (.A(n_18940),
    .Y(n_15641));
 XNOR2x1_ASAP7_75t_SL g23614 (.B(n_18800),
    .Y(n_15651),
    .A(n_19043));
 XNOR2xp5_ASAP7_75t_SL g23683 (.A(n_12831),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_89),
    .Y(n_15719));
 MAJx2_ASAP7_75t_SL g23684 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_693),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_757),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_597),
    .Y(n_15720));
 OAI21xp5_ASAP7_75t_SL g23770 (.A1(n_15813),
    .A2(n_19382),
    .B(n_15815),
    .Y(n_15816));
 NAND2x1p5_ASAP7_75t_SL g23771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_264),
    .B(n_10533),
    .Y(n_15813));
 NAND2xp5_ASAP7_75t_SL g23773 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263),
    .Y(n_15815));
 OAI22xp5_ASAP7_75t_SL g238 (.A1(n_10908),
    .A2(n_11359),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_166),
    .B2(n_11356),
    .Y(n_11357));
 NAND2xp5_ASAP7_75t_SL g23834 (.A(n_12088),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_400),
    .Y(n_15886));
 XNOR2x1_ASAP7_75t_SL g23866 (.B(n_15921),
    .Y(n_15922),
    .A(n_15920));
 MAJx2_ASAP7_75t_SL g23867 (.A(n_11752),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_39),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_98),
    .Y(n_15920));
 NAND2x1_ASAP7_75t_SL g23868 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(n_15014),
    .Y(n_15921));
 MAJx2_ASAP7_75t_SL g23885 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_284),
    .B(n_17489),
    .C(n_3782),
    .Y(n_15939));
 XNOR2xp5_ASAP7_75t_SL g239 (.A(n_19341),
    .B(n_19138),
    .Y(n_6125));
 AO21x1_ASAP7_75t_SL g23903 (.A1(n_21553),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_278),
    .B(n_21554),
    .Y(n_15962));
 INVxp67_ASAP7_75t_SL g23905 (.A(n_21554),
    .Y(n_15960));
 XNOR2xp5_ASAP7_75t_SL g23940 (.A(n_24107),
    .B(n_15999),
    .Y(n_16000));
 AND2x2_ASAP7_75t_SL g23942 (.A(n_2182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_556),
    .Y(n_15999));
 XOR2xp5_ASAP7_75t_SL g23996 (.A(n_16058),
    .B(n_16059),
    .Y(n_16060));
 MAJIxp5_ASAP7_75t_SL g23997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_267),
    .B(n_4070),
    .C(n_22995),
    .Y(n_16058));
 OAI21xp5_ASAP7_75t_SL g23998 (.A1(n_21978),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(n_16059));
 XNOR2xp5_ASAP7_75t_SL g23999 (.A(n_22873),
    .B(n_16062),
    .Y(n_16063));
 OAI21xp5_ASAP7_75t_SL g24 (.A1(n_20162),
    .A2(n_20163),
    .B(n_9661),
    .Y(n_20164));
 INVx1_ASAP7_75t_SL g240 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_37),
    .Y(n_19307));
 NAND2xp5_ASAP7_75t_SL g24001 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(n_3479),
    .Y(n_16062));
 AOI21xp5_ASAP7_75t_SL g24007 (.A1(n_16069),
    .A2(n_16070),
    .B(n_7716),
    .Y(n_16071));
 NAND2x1_ASAP7_75t_SL g24008 (.A(n_10395),
    .B(n_23092),
    .Y(n_16069));
 XNOR2xp5_ASAP7_75t_SL g24076 (.A(n_16140),
    .B(n_19016),
    .Y(n_16142));
 XNOR2xp5_ASAP7_75t_SL g24077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_119),
    .Y(n_16140));
 OAI22xp5_ASAP7_75t_SL g24087 (.A1(n_18009),
    .A2(n_8959),
    .B1(n_18008),
    .B2(n_10527),
    .Y(n_16149));
 AND2x2_ASAP7_75t_SL g24092 (.A(n_8588),
    .B(n_8586),
    .Y(n_16155));
 NOR2xp67_ASAP7_75t_SL g24093 (.A(n_8588),
    .B(n_8586),
    .Y(n_16156));
 NOR3xp33_ASAP7_75t_SL g24097 (.A(n_16155),
    .B(n_16156),
    .C(n_18954),
    .Y(n_16158));
 AOI21xp5_ASAP7_75t_SL g24099 (.A1(n_12774),
    .A2(n_12775),
    .B(n_16158),
    .Y(n_16162));
 INVx1_ASAP7_75t_SL g241 (.A(n_23431),
    .Y(n_6131));
 XNOR2xp5_ASAP7_75t_SL g24164 (.A(n_16226),
    .B(n_16227),
    .Y(n_16228));
 NAND2xp5_ASAP7_75t_SL g24165 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_786),
    .Y(n_16226));
 NAND2xp5_ASAP7_75t_SL g24166 (.A(n_2181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_562),
    .Y(n_16227));
 INVxp67_ASAP7_75t_SL g24167 (.A(n_16226),
    .Y(n_9978));
 INVx1_ASAP7_75t_SL g24168 (.A(n_16227),
    .Y(n_16230));
 AO21x2_ASAP7_75t_SL g24187 (.A1(n_22323),
    .A2(n_21319),
    .B(n_21318),
    .Y(n_16253));
 OAI331xp33_ASAP7_75t_SL g24189 (.A1(n_16255),
    .A2(n_16253),
    .A3(n_5332),
    .B1(n_5332),
    .B2(n_16257),
    .B3(n_16256),
    .C1(n_16258),
    .Y(n_16259));
 INVx1_ASAP7_75t_SL g24192 (.A(n_16255),
    .Y(n_16257));
 OR2x2_ASAP7_75t_SL g24193 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[16]),
    .B(n_17936),
    .Y(n_16258));
 XOR2xp5_ASAP7_75t_SL g242 (.A(n_12419),
    .B(n_18985),
    .Y(n_4487));
 INVxp33_ASAP7_75t_SL g24251 (.A(n_21126),
    .Y(n_16319));
 NAND2xp5_ASAP7_75t_SL g24256 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_205),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_224),
    .Y(n_16324));
 OAI21xp5_ASAP7_75t_SL g24257 (.A1(n_5412),
    .A2(n_8347),
    .B(n_8349),
    .Y(n_16325));
 NOR2xp67_ASAP7_75t_SL g24258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_205),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_224),
    .Y(n_16326));
 XNOR2x2_ASAP7_75t_SL g24278 (.A(n_14857),
    .B(n_19035),
    .Y(n_16347));
 XNOR2xp5_ASAP7_75t_SL g24280 (.A(n_16347),
    .B(n_16348),
    .Y(n_16349));
 XNOR2xp5_ASAP7_75t_SL g24281 (.A(n_9420),
    .B(n_20376),
    .Y(n_16348));
 XNOR2xp5_ASAP7_75t_SL g24296 (.A(n_16365),
    .B(n_20936),
    .Y(n_16367));
 MAJIxp5_ASAP7_75t_SL g24297 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_41),
    .Y(n_16365));
 XNOR2x1_ASAP7_75t_SL g243 (.B(n_20987),
    .Y(n_20988),
    .A(n_20984));
 NOR2xp33_ASAP7_75t_SL g24348 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[13]),
    .B(n_17869),
    .Y(n_16418));
 OR2x2_ASAP7_75t_SL g24384 (.A(n_19205),
    .B(n_17654),
    .Y(n_16456));
 XNOR2xp5_ASAP7_75t_SL g24390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_88),
    .B(n_19045),
    .Y(n_16466));
 OAI21xp5_ASAP7_75t_SL g24399 (.A1(n_16681),
    .A2(n_18802),
    .B(n_16476),
    .Y(n_16477));
 HB1xp67_ASAP7_75t_SL g244 (.A(n_6593),
    .Y(n_6599));
 AOI21xp33_ASAP7_75t_SL g24401 (.A1(n_16681),
    .A2(n_16475),
    .B(n_9305),
    .Y(n_16476));
 NOR2xp33_ASAP7_75t_SL g24402 (.A(n_5332),
    .B(n_24027),
    .Y(n_16475));
 AOI22xp5_ASAP7_75t_SL g24451 (.A1(n_16528),
    .A2(n_17936),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[9]),
    .Y(n_16529));
 INVxp67_ASAP7_75t_SL g24453 (.A(n_16071),
    .Y(n_16530));
 NAND2xp33_ASAP7_75t_SL g24454 (.A(n_17874),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_436),
    .Y(n_16532));
 NAND2xp5_ASAP7_75t_SL g24456 (.A(n_16533),
    .B(n_17874),
    .Y(n_16534));
 INVx1_ASAP7_75t_SL g24457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_436),
    .Y(n_16533));
 OR2x2_ASAP7_75t_SL g24458 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[9]),
    .B(n_17874),
    .Y(n_16535));
 AOI22xp5_ASAP7_75t_SL g24462 (.A1(n_16540),
    .A2(n_17936),
    .B1(n_5332),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[13]),
    .Y(n_16541));
 XNOR2x1_ASAP7_75t_SL g24475 (.B(n_18897),
    .Y(n_16557),
    .A(n_8007));
 MAJx2_ASAP7_75t_SL g24477 (.A(n_20872),
    .B(n_20869),
    .C(n_2764),
    .Y(n_16558));
 XOR2x2_ASAP7_75t_SL g24478 (.A(n_21355),
    .B(n_6453),
    .Y(n_16559));
 AO21x1_ASAP7_75t_SL g24479 (.A1(n_16558),
    .A2(n_16559),
    .B(n_16676),
    .Y(n_16561));
 INVxp67_ASAP7_75t_SL g24484 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_259),
    .Y(n_16563));
 OA21x2_ASAP7_75t_SL g24485 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_274),
    .A2(n_6976),
    .B(n_24917),
    .Y(n_16564));
 INVxp67_ASAP7_75t_SL g24486 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_261),
    .Y(n_16565));
 MAJIxp5_ASAP7_75t_SL g245 (.A(n_14045),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_34),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_15),
    .Y(n_12412));
 AOI21xp5_ASAP7_75t_SL g24500 (.A1(n_25833),
    .A2(n_21881),
    .B(n_21882),
    .Y(n_16579));
 XNOR2xp5_ASAP7_75t_SL g24515 (.A(n_22853),
    .B(n_16596),
    .Y(n_16597));
 AO21x1_ASAP7_75t_SL g24517 (.A1(n_3987),
    .A2(n_3938),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_424),
    .Y(n_16596));
 OAI311xp33_ASAP7_75t_SL g24532 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_451),
    .A2(n_10455),
    .A3(n_17870),
    .B1(n_16615),
    .C1(n_16614),
    .Y(n_16616));
 OR2x2_ASAP7_75t_SL g24535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[14]),
    .B(n_17869),
    .Y(n_16614));
 NAND3xp33_ASAP7_75t_SL g24536 (.A(n_17869),
    .B(n_10455),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_451),
    .Y(n_16615));
 INVx1_ASAP7_75t_SL g24583 (.A(n_16663),
    .Y(n_16664));
 AOI21x1_ASAP7_75t_SL g24584 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_28),
    .A2(n_7858),
    .B(n_7855),
    .Y(n_16663));
 NOR2x1_ASAP7_75t_SL g24594 (.A(n_16558),
    .B(n_16559),
    .Y(n_16676));
 AOI21xp5_ASAP7_75t_SL g24595 (.A1(n_24021),
    .A2(n_23266),
    .B(n_22324),
    .Y(n_16681));
 XNOR2xp5_ASAP7_75t_SL g246 (.A(n_8670),
    .B(n_8673),
    .Y(n_8674));
 XNOR2xp5_ASAP7_75t_SL g24621 (.A(n_16705),
    .B(n_16706),
    .Y(n_16707));
 XOR2x2_ASAP7_75t_SL g24622 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_277),
    .B(n_12887),
    .Y(n_16705));
 NAND2xp5_ASAP7_75t_SL g24623 (.A(n_6727),
    .B(n_11454),
    .Y(n_16706));
 MAJIxp5_ASAP7_75t_SL g24671 (.A(n_16779),
    .B(n_16780),
    .C(n_16781),
    .Y(n_16782));
 INVx1_ASAP7_75t_SL g24672 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_332),
    .Y(n_16779));
 INVxp67_ASAP7_75t_SL g24673 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .Y(n_16780));
 INVxp67_ASAP7_75t_SL g24674 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_291),
    .Y(n_16781));
 XOR2xp5_ASAP7_75t_SL g24675 (.A(n_10171),
    .B(n_16784),
    .Y(n_16785));
 INVx1_ASAP7_75t_SL g24676 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_32),
    .Y(n_16784));
 XOR2xp5_ASAP7_75t_SL g247 (.A(n_8671),
    .B(n_8672),
    .Y(n_8673));
 INVxp67_ASAP7_75t_SRAM g248 (.A(n_8671),
    .Y(n_5400));
 NAND2xp5_ASAP7_75t_SL g249 (.A(n_19182),
    .B(n_2159),
    .Y(n_8671));
 BUFx4f_ASAP7_75t_SL g24905 (.A(n_12981),
    .Y(n_6879));
 XNOR2xp5_ASAP7_75t_SL g24906 (.A(n_17020),
    .B(n_26091),
    .Y(n_17024));
 INVx1_ASAP7_75t_SL g24907 (.A(n_17019),
    .Y(n_17020));
 AND2x2_ASAP7_75t_SL g24908 (.A(n_6879),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_748),
    .Y(n_17019));
 XNOR2xp5_ASAP7_75t_SL g24941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_142),
    .B(n_19861),
    .Y(n_17057));
 OR2x2_ASAP7_75t_SL g24947 (.A(n_18704),
    .B(n_12050),
    .Y(n_17063));
 MAJIxp5_ASAP7_75t_SL g24951 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_565),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_725),
    .Y(n_17064));
 XOR2xp5_ASAP7_75t_SL g24952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_627),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_659),
    .Y(n_17066));
 NOR2xp67_ASAP7_75t_SL g24958 (.A(n_16782),
    .B(n_16785),
    .Y(n_17073));
 AND2x2_ASAP7_75t_SL g25 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_317),
    .B(n_20161),
    .Y(n_20162));
 AND2x2_ASAP7_75t_SL g250 (.A(n_9259),
    .B(n_8016),
    .Y(n_11746));
 XOR2x2_ASAP7_75t_SL g251 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_95),
    .Y(n_12397));
 OR2x2_ASAP7_75t_SL g25123 (.A(n_46),
    .B(n_445),
    .Y(n_17240));
 NAND2xp5_ASAP7_75t_SL g25125 (.A(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .Y(n_17241));
 INVxp67_ASAP7_75t_SL g25126 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .Y(n_17242));
 NOR2xp33_ASAP7_75t_SL g252 (.A(n_9973),
    .B(n_13971),
    .Y(n_8196));
 XNOR2xp5_ASAP7_75t_SL g25275 (.A(n_17066),
    .B(n_17400),
    .Y(n_17401));
 OAI22xp5_ASAP7_75t_SL g25276 (.A1(n_17398),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_154),
    .B1(n_17397),
    .B2(n_17064),
    .Y(n_17400));
 INVx1_ASAP7_75t_SL g25277 (.A(n_17397),
    .Y(n_17398));
 MAJIxp5_ASAP7_75t_SL g25278 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_661),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_629),
    .Y(n_17397));
 INVx2_ASAP7_75t_SL g25279 (.A(n_17064),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_154));
 OAI22xp5_ASAP7_75t_SL g25280 (.A1(n_17064),
    .A2(n_17066),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_154),
    .B2(n_17403),
    .Y(n_17404));
 INVx1_ASAP7_75t_SL g25282 (.A(n_17066),
    .Y(n_17403));
 XNOR2xp5_ASAP7_75t_SL g25289 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .B(n_18842),
    .Y(n_17413));
 MAJx2_ASAP7_75t_SL g25290 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_545),
    .B(n_24712),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117));
 INVx1_ASAP7_75t_SL g25292 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .Y(n_17414));
 NAND2xp5_ASAP7_75t_SL g253 (.A(n_13971),
    .B(n_9973),
    .Y(n_8197));
 XNOR2xp5_ASAP7_75t_SL g25314 (.A(n_17440),
    .B(n_17441),
    .Y(n_17442));
 MAJIxp5_ASAP7_75t_SL g25315 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_298),
    .B(n_14110),
    .C(n_2580),
    .Y(n_17440));
 AOI22xp5_ASAP7_75t_SL g25316 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .A2(n_26077),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .B2(n_3457),
    .Y(n_17441));
 XOR2xp5_ASAP7_75t_SL g25356 (.A(n_17486),
    .B(n_17487),
    .Y(n_17488));
 MAJIxp5_ASAP7_75t_SL g25357 (.A(n_13720),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_65),
    .Y(n_17486));
 AO22x2_ASAP7_75t_SL g25358 (.A1(n_8326),
    .A2(n_8325),
    .B1(n_8324),
    .B2(n_8323),
    .Y(n_17487));
 XNOR2xp5_ASAP7_75t_SL g25359 (.A(n_17490),
    .B(n_17491),
    .Y(n_17492));
 INVx1_ASAP7_75t_SL g25360 (.A(n_17489),
    .Y(n_17490));
 MAJIxp5_ASAP7_75t_SL g25361 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_74),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_72),
    .Y(n_17489));
 XNOR2x1_ASAP7_75t_SL g25362 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_197),
    .Y(n_17491),
    .A(n_11023));
 MAJx2_ASAP7_75t_SL g25418 (.A(n_9653),
    .B(n_17551),
    .C(n_9651),
    .Y(n_17552));
 NAND2xp5_ASAP7_75t_SL g25419 (.A(n_2174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_748),
    .Y(n_17551));
 INVx1_ASAP7_75t_SL g25420 (.A(n_17551),
    .Y(n_17553));
 OA21x2_ASAP7_75t_SL g25425 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_290),
    .A2(n_10954),
    .B(n_14695),
    .Y(n_17559));
 INVx1_ASAP7_75t_SL g25426 (.A(n_14695),
    .Y(n_17560));
 NAND2xp5_ASAP7_75t_SL g25516 (.A(n_19205),
    .B(n_17654),
    .Y(n_17655));
 AND2x2_ASAP7_75t_SL g25518 (.A(n_11550),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .Y(n_17651));
 XNOR2xp5_ASAP7_75t_SL g25520 (.A(n_10046),
    .B(n_18765),
    .Y(n_17654));
 MAJx2_ASAP7_75t_SL g25526 (.A(n_9827),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .C(n_2897),
    .Y(n_17661));
 NOR2x1_ASAP7_75t_SL g25529 (.A(n_17661),
    .B(n_20873),
    .Y(n_17663));
 AOI21x1_ASAP7_75t_SL g25534 (.A1(n_4349),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_249),
    .B(n_17669),
    .Y(n_17670));
 OAI21xp5_ASAP7_75t_SL g25539 (.A1(n_8624),
    .A2(n_17670),
    .B(n_8629),
    .Y(n_17673));
 XNOR2xp5_ASAP7_75t_SL g25579 (.A(n_20688),
    .B(n_9218),
    .Y(n_17712));
 OR2x2_ASAP7_75t_SL g256 (.A(n_10256),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_301),
    .Y(n_10261));
 XNOR2xp5_ASAP7_75t_SL g25601 (.A(n_17732),
    .B(n_17733),
    .Y(n_17734));
 AND2x2_ASAP7_75t_SL g25602 (.A(n_2162),
    .B(n_13612),
    .Y(n_17732));
 NAND2x1_ASAP7_75t_SL g25603 (.A(n_2159),
    .B(n_11496),
    .Y(n_17733));
 INVx1_ASAP7_75t_SL g25604 (.A(n_17733),
    .Y(n_17735));
 NAND3xp33_ASAP7_75t_SL g25638 (.A(n_17772),
    .B(n_17773),
    .C(n_17774),
    .Y(n_17775));
 NAND3xp33_ASAP7_75t_SL g25639 (.A(n_14894),
    .B(n_16685),
    .C(n_14891),
    .Y(n_17772));
 OAI21xp33_ASAP7_75t_SL g25640 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_425),
    .A2(n_16684),
    .B(n_14897),
    .Y(n_17773));
 AOI21xp33_ASAP7_75t_SL g25641 (.A1(n_14894),
    .A2(n_14893),
    .B(n_16418),
    .Y(n_17774));
 MAJIxp5_ASAP7_75t_SL g25676 (.A(n_22958),
    .B(n_11545),
    .C(n_11546),
    .Y(n_17808));
 AO21x1_ASAP7_75t_SL g25694 (.A1(n_17829),
    .A2(n_17830),
    .B(n_17831),
    .Y(n_17832));
 NAND2xp5_ASAP7_75t_SL g25695 (.A(n_20728),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_246),
    .Y(n_17829));
 OAI21xp5_ASAP7_75t_SL g25696 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_247),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_249),
    .Y(n_17830));
 NOR2xp67_ASAP7_75t_SL g25697 (.A(n_20728),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_246),
    .Y(n_17831));
 OAI211xp5_ASAP7_75t_SL g25727 (.A1(n_17863),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_490),
    .B(n_17867),
    .C(n_17866),
    .Y(n_17868));
 NAND2xp5_ASAP7_75t_SL g25728 (.A(n_25130),
    .B(n_23932),
    .Y(n_17863));
 NAND2xp5_ASAP7_75t_SL g25730 (.A(n_17865),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_490),
    .Y(n_17866));
 NOR2xp33_ASAP7_75t_SL g25731 (.A(n_25130),
    .B(n_17882),
    .Y(n_17865));
 OR2x2_ASAP7_75t_SL g25733 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[11]),
    .B(n_23932),
    .Y(n_17867));
 OAI322xp33_ASAP7_75t_SL g25734 (.A1(n_16160),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_436),
    .A3(n_17870),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[9]),
    .B2(n_17869),
    .C1(n_17871),
    .C2(n_17872),
    .Y(n_17873));
 INVx3_ASAP7_75t_SL g25735 (.A(n_17869),
    .Y(n_17870));
 AND2x6_ASAP7_75t_SL g25736 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_pvld[7]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_pvld[7]),
    .Y(n_17869));
 NAND2xp5_ASAP7_75t_SL g25737 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_436),
    .Y(n_17871));
 INVxp67_ASAP7_75t_SL g25738 (.A(n_16160),
    .Y(n_17872));
 OAI21xp33_ASAP7_75t_SL g25739 (.A1(n_17875),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_494),
    .B(n_17879),
    .Y(n_17880));
 NAND2xp5_ASAP7_75t_SL g25740 (.A(n_17874),
    .B(n_20280),
    .Y(n_17875));
 BUFx8_ASAP7_75t_L g25741 (.A(n_2146),
    .Y(n_17874));
 AOI21xp5_ASAP7_75t_SL g25742 (.A1(n_17877),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_494),
    .B(n_17878),
    .Y(n_17879));
 NOR2xp33_ASAP7_75t_SL g25743 (.A(n_17876),
    .B(n_20280),
    .Y(n_17877));
 INVx3_ASAP7_75t_SL g25744 (.A(n_17874),
    .Y(n_17876));
 NOR2xp33_ASAP7_75t_SL g25745 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[13]),
    .B(n_17874),
    .Y(n_17878));
 OAI321xp33_ASAP7_75t_SL g25746 (.A1(n_19983),
    .A2(n_16579),
    .A3(n_17882),
    .B1(n_17884),
    .B2(n_17883),
    .C(n_17885),
    .Y(n_17886));
 INVx6_ASAP7_75t_L g25747 (.A(n_23932),
    .Y(n_17882));
 NAND2xp5_ASAP7_75t_SL g25749 (.A(n_23932),
    .B(n_19983),
    .Y(n_17883));
 INVx1_ASAP7_75t_SL g25750 (.A(n_16579),
    .Y(n_17884));
 OR2x2_ASAP7_75t_SL g25751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[13]),
    .B(n_23932),
    .Y(n_17885));
 AOI22xp5_ASAP7_75t_SL g25772 (.A1(n_17909),
    .A2(n_17874),
    .B1(n_17876),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[10]),
    .Y(n_17910));
 OAI322xp33_ASAP7_75t_SL g25801 (.A1(n_5332),
    .A2(n_13570),
    .A3(n_20738),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[14]),
    .B2(n_17936),
    .C1(n_17939),
    .C2(n_17938),
    .Y(n_17940));
 INVx6_ASAP7_75t_SL g25802 (.A(n_17936),
    .Y(n_5332));
 BUFx8_ASAP7_75t_L g25803 (.A(n_9301),
    .Y(n_17936));
 INVxp67_ASAP7_75t_SL g25804 (.A(n_20738),
    .Y(n_17938));
 NAND2xp5_ASAP7_75t_SL g25805 (.A(n_13570),
    .B(n_17936),
    .Y(n_17939));
 XNOR2x1_ASAP7_75t_SL g25841 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_125),
    .Y(n_17976),
    .A(n_22883));
 MAJIxp5_ASAP7_75t_SL g25842 (.A(n_17978),
    .B(n_7237),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_174),
    .Y(n_17979));
 XNOR2xp5_ASAP7_75t_SL g25843 (.A(n_17976),
    .B(n_17977),
    .Y(n_17978));
 AOI22xp5_ASAP7_75t_SL g25844 (.A1(n_11458),
    .A2(n_11462),
    .B1(n_11463),
    .B2(n_18972),
    .Y(n_17977));
 XNOR2xp5_ASAP7_75t_SL g25861 (.A(n_14871),
    .B(n_14874),
    .Y(n_17997));
 INVx1_ASAP7_75t_SL g25862 (.A(n_17997),
    .Y(n_17998));
 NAND3xp33_ASAP7_75t_SL g25866 (.A(n_8167),
    .B(n_8292),
    .C(n_13363),
    .Y(n_18002));
 INVxp33_ASAP7_75t_SRAM g25867 (.A(n_8292),
    .Y(n_18004));
 INVx1_ASAP7_75t_SL g25871 (.A(n_18008),
    .Y(n_18009));
 XOR2xp5_ASAP7_75t_SL g25872 (.A(n_8674),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_247),
    .Y(n_18008));
 MAJx2_ASAP7_75t_SL g25892 (.A(n_18063),
    .B(n_18065),
    .C(n_18068),
    .Y(n_18069));
 MAJx2_ASAP7_75t_SL g25893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_138),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_164),
    .Y(n_18063));
 INVxp67_ASAP7_75t_SL g25894 (.A(n_18064),
    .Y(n_18065));
 MAJIxp5_ASAP7_75t_SL g25895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_659),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_627),
    .Y(n_18064));
 INVxp67_ASAP7_75t_SL g25896 (.A(n_18067),
    .Y(n_18068));
 XNOR2x1_ASAP7_75t_SL g25897 (.B(n_18803),
    .Y(n_18067),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_100));
 XOR2xp5_ASAP7_75t_SL g259 (.A(n_6872),
    .B(n_6877),
    .Y(n_6878));
 XOR2xp5_ASAP7_75t_SL g25917 (.A(n_18092),
    .B(n_18093),
    .Y(n_18094));
 INVx1_ASAP7_75t_SL g25918 (.A(n_18091),
    .Y(n_18092));
 MAJx2_ASAP7_75t_SL g25919 (.A(n_18899),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_20),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_17),
    .Y(n_18091));
 XNOR2xp5_ASAP7_75t_SL g25920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_171),
    .B(n_8003),
    .Y(n_18093));
 INVxp67_ASAP7_75t_SRAM g25921 (.A(n_18093),
    .Y(n_3729));
 XNOR2xp5_ASAP7_75t_SL g25947 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_147),
    .B(n_22073),
    .Y(n_18124));
 XNOR2xp5_ASAP7_75t_SL g25966 (.A(n_18141),
    .B(n_19206),
    .Y(n_18144));
 XOR2xp5_ASAP7_75t_SL g25968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_125),
    .Y(n_18141));
 AO21x2_ASAP7_75t_SL g25987 (.A1(n_18165),
    .A2(n_18166),
    .B(n_18167),
    .Y(n_18168));
 NAND2xp67_ASAP7_75t_SL g25988 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_209),
    .B(n_11622),
    .Y(n_18165));
 OAI21xp5_ASAP7_75t_SL g25989 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_229),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_228),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_231),
    .Y(n_18166));
 NOR2x1_ASAP7_75t_SL g25990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_209),
    .B(n_11622),
    .Y(n_18167));
 MAJx2_ASAP7_75t_SL g25997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_75),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_35),
    .Y(n_18175));
 NAND2xp5_ASAP7_75t_SL g26 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_266),
    .B(n_26118),
    .Y(n_20082));
 XNOR2x1_ASAP7_75t_SL g262 (.B(n_10601),
    .Y(n_19268),
    .A(n_4967));
 MAJIxp5_ASAP7_75t_SL g263 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_126),
    .B(n_21800),
    .C(n_21801),
    .Y(n_11413));
 MAJIxp5_ASAP7_75t_SL g26371 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_717),
    .B(n_18579),
    .C(n_5681),
    .Y(n_18582));
 NOR2xp33_ASAP7_75t_SL g26447 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_182),
    .Y(n_18666));
 NOR2xp33_ASAP7_75t_SL g26448 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_253),
    .B(n_10220),
    .Y(n_18667));
 MAJIxp5_ASAP7_75t_SL g26451 (.A(n_15149),
    .B(n_15150),
    .C(n_15151),
    .Y(n_6833));
 HB1xp67_ASAP7_75t_SL g26466 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .Y(n_18692));
 OR2x2_ASAP7_75t_SL g26471 (.A(n_15169),
    .B(n_15172),
    .Y(n_18698));
 MAJx2_ASAP7_75t_SL g26472 (.A(n_16466),
    .B(n_12293),
    .C(n_19566),
    .Y(n_18699));
 MAJx2_ASAP7_75t_SL g26473 (.A(n_18141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_132),
    .C(n_18175),
    .Y(n_18700));
 MAJx2_ASAP7_75t_SL g26474 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_19),
    .Y(n_18701));
 AND2x2_ASAP7_75t_SL g26475 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B(n_3709),
    .Y(n_18702));
 MAJx2_ASAP7_75t_SL g26476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_19),
    .Y(n_18703));
 MAJx2_ASAP7_75t_SL g26477 (.A(n_20018),
    .B(n_14174),
    .C(n_14912),
    .Y(n_18704));
 AND2x2_ASAP7_75t_SL g26478 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .Y(n_14158));
 AND2x2_ASAP7_75t_SL g26480 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(n_18707));
 AND2x2_ASAP7_75t_SL g26483 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .B(n_9273),
    .Y(n_18710));
 AND2x2_ASAP7_75t_SL g26484 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(n_14674),
    .Y(n_18711));
 AND2x2_ASAP7_75t_SL g26485 (.A(n_21224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_282),
    .Y(n_18712));
 AND2x2_ASAP7_75t_SL g26489 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_282),
    .Y(n_18716));
 NAND2xp5_ASAP7_75t_SL g26490 (.A(n_11021),
    .B(n_8158),
    .Y(n_18717));
 AND2x2_ASAP7_75t_SL g26491 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B(n_3706),
    .Y(n_18718));
 MAJx2_ASAP7_75t_SL g26492 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_19),
    .Y(n_18719));
 AND2x2_ASAP7_75t_SL g26493 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_18720));
 XOR2xp5_ASAP7_75t_SL g26494 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_379),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_387),
    .Y(n_18721));
 MAJx2_ASAP7_75t_SL g26499 (.A(n_22443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_120),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .Y(n_18726));
 MAJx2_ASAP7_75t_SL g265 (.A(n_4518),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_30),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_152),
    .Y(n_11412));
 MAJIxp5_ASAP7_75t_SL g26502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_753),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_689),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_593),
    .Y(n_18729));
 OR2x2_ASAP7_75t_SL g26503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_277),
    .B(n_10744),
    .Y(n_18730));
 MAJx2_ASAP7_75t_SL g26504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_94),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_85),
    .Y(n_18731));
 XNOR2xp5_ASAP7_75t_SL g26505 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_115),
    .Y(n_18732));
 MAJx2_ASAP7_75t_SL g26510 (.A(n_12934),
    .B(n_7382),
    .C(n_7383),
    .Y(n_18737));
 MAJx2_ASAP7_75t_SL g26511 (.A(n_7612),
    .B(n_7608),
    .C(n_21668),
    .Y(n_18738));
 AND2x2_ASAP7_75t_SL g26512 (.A(n_22865),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .Y(n_18739));
 MAJx2_ASAP7_75t_SL g26513 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_94),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_85),
    .Y(n_18740));
 MAJx2_ASAP7_75t_SL g26521 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_143),
    .C(n_15070),
    .Y(n_18748));
 OR2x2_ASAP7_75t_SL g26522 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_144),
    .Y(n_18749));
 AND2x2_ASAP7_75t_SL g26524 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .Y(n_18751));
 XOR2xp5_ASAP7_75t_SL g26525 (.A(n_13598),
    .B(n_13111),
    .Y(n_18752));
 OA21x2_ASAP7_75t_SL g26526 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_258),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_261),
    .Y(n_18753));
 AND2x2_ASAP7_75t_SL g26527 (.A(n_2930),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .Y(n_18754));
 AND2x2_ASAP7_75t_SL g26529 (.A(n_3528),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .Y(n_18756));
 XNOR2xp5_ASAP7_75t_SL g26530 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_6),
    .Y(n_18757));
 MAJx2_ASAP7_75t_SL g26531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_150),
    .B(n_20882),
    .C(n_20885),
    .Y(n_18758));
 NAND2xp5_ASAP7_75t_SL g26533 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_94),
    .Y(n_18760));
 AO21x1_ASAP7_75t_SL g26534 (.A1(n_13196),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252),
    .B(n_20680),
    .Y(n_18761));
 AND2x2_ASAP7_75t_SL g26536 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_194),
    .Y(n_18763));
 MAJx2_ASAP7_75t_SL g26537 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_691),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_595),
    .Y(n_18764));
 XOR2xp5_ASAP7_75t_SL g26538 (.A(n_17808),
    .B(n_19049),
    .Y(n_18765));
 XNOR2xp5_ASAP7_75t_SL g26539 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_201),
    .Y(n_18766));
 AO21x1_ASAP7_75t_SL g26540 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_213),
    .Y(n_18767));
 OR2x2_ASAP7_75t_SL g26542 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_257),
    .Y(n_18769));
 OR2x2_ASAP7_75t_SL g26543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_257),
    .Y(n_18770));
 NAND2xp5_ASAP7_75t_SL g26544 (.A(n_21873),
    .B(n_22740),
    .Y(n_18771));
 AO21x1_ASAP7_75t_SL g26547 (.A1(n_22969),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_217),
    .B(n_19174),
    .Y(n_18774));
 MAJx2_ASAP7_75t_SL g26548 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_58),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_75),
    .Y(n_18775));
 MAJx2_ASAP7_75t_SL g26549 (.A(n_19310),
    .B(n_19306),
    .C(n_19316),
    .Y(n_18776));
 AND2x2_ASAP7_75t_SL g26551 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(n_2359),
    .Y(n_18778));
 AND2x2_ASAP7_75t_SL g26552 (.A(n_5329),
    .B(n_5332),
    .Y(n_18779));
 MAJIxp5_ASAP7_75t_SL g26553 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_131),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_139),
    .Y(n_18780));
 XOR2x2_ASAP7_75t_SL g26554 (.A(n_19681),
    .B(n_11438),
    .Y(n_18781));
 XOR2xp5_ASAP7_75t_SL g26555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_751),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_12),
    .Y(n_18782));
 AO21x1_ASAP7_75t_SL g26556 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_213),
    .Y(n_18783));
 AO21x1_ASAP7_75t_SL g26558 (.A1(n_4771),
    .A2(n_4772),
    .B(n_4773),
    .Y(n_18785));
 MAJx2_ASAP7_75t_SL g26559 (.A(n_19621),
    .B(n_21163),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_176),
    .Y(n_18786));
 AND2x2_ASAP7_75t_SL g26560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_8),
    .Y(n_18787));
 MAJx2_ASAP7_75t_SL g26563 (.A(n_20990),
    .B(n_20989),
    .C(n_20984),
    .Y(n_18790));
 MAJx2_ASAP7_75t_SL g26564 (.A(n_2429),
    .B(n_25598),
    .C(n_7371),
    .Y(n_18791));
 MAJx2_ASAP7_75t_SL g26565 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_113),
    .B(n_21520),
    .C(n_9155),
    .Y(n_14411));
 MAJx2_ASAP7_75t_SL g26566 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_785),
    .C(n_12878),
    .Y(n_18793));
 MAJx2_ASAP7_75t_SL g26567 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_64),
    .Y(n_18794));
 XNOR2x1_ASAP7_75t_SL g26568 (.B(n_14713),
    .Y(n_18795),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_115));
 MAJx2_ASAP7_75t_SL g26570 (.A(n_18765),
    .B(n_4539),
    .C(n_13519),
    .Y(n_18797));
 AND2x2_ASAP7_75t_SL g26571 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(n_19411),
    .Y(n_18798));
 AND2x2_ASAP7_75t_SL g26572 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(n_18799));
 MAJx2_ASAP7_75t_SL g26573 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_789),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_565),
    .Y(n_18800));
 NAND2xp5_ASAP7_75t_SL g26575 (.A(n_24027),
    .B(n_9301),
    .Y(n_18802));
 MAJx2_ASAP7_75t_SL g26576 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_563),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_723),
    .C(n_11379),
    .Y(n_18803));
 XOR2xp5_ASAP7_75t_SL g26577 (.A(n_16684),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_458),
    .Y(n_18804));
 XNOR2xp5_ASAP7_75t_SL g26579 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_166),
    .Y(n_18806));
 XNOR2xp5_ASAP7_75t_SL g26580 (.A(n_14725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_45),
    .Y(n_18807));
 XNOR2xp5_ASAP7_75t_SL g26582 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_132),
    .B(n_10295),
    .Y(n_18809));
 XNOR2xp5_ASAP7_75t_SL g26584 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_30),
    .B(n_10608),
    .Y(n_18811));
 XNOR2xp5_ASAP7_75t_SL g26585 (.A(n_6932),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_77),
    .Y(n_18812));
 OR2x2_ASAP7_75t_SL g26588 (.A(n_10666),
    .B(n_10117),
    .Y(n_18815));
 OR2x2_ASAP7_75t_SL g26590 (.A(n_21247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_375),
    .Y(n_10627));
 XOR2xp5_ASAP7_75t_SL g26592 (.A(n_14671),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_55),
    .Y(n_18819));
 NOR2xp33_ASAP7_75t_SL g26593 (.A(n_10774),
    .B(n_19605),
    .Y(n_18820));
 XNOR2xp5_ASAP7_75t_SL g26595 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_113),
    .B(n_12581),
    .Y(n_18822));
 XOR2xp5_ASAP7_75t_SL g26596 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .B(n_11550),
    .Y(n_18823));
 XOR2xp5_ASAP7_75t_SL g26598 (.A(n_11593),
    .B(n_18902),
    .Y(n_18825));
 XNOR2xp5_ASAP7_75t_SL g26599 (.A(n_9344),
    .B(n_9342),
    .Y(n_18826));
 OR3x1_ASAP7_75t_SL g266 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_291),
    .B(n_20361),
    .C(n_20362),
    .Y(n_20363));
 XNOR2xp5_ASAP7_75t_SL g26600 (.A(n_22876),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_68),
    .Y(n_18827));
 OR2x2_ASAP7_75t_SL g26601 (.A(n_2564),
    .B(n_10340),
    .Y(n_18828));
 XOR2xp5_ASAP7_75t_SL g26604 (.A(n_9658),
    .B(n_9657),
    .Y(n_18831));
 XNOR2xp5_ASAP7_75t_SL g26605 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_86),
    .Y(n_18832));
 XNOR2xp5_ASAP7_75t_SL g26608 (.A(n_5529),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_87),
    .Y(n_18835));
 XNOR2x2_ASAP7_75t_SL g26609 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_79),
    .B(n_13244),
    .Y(n_18836));
 XOR2xp5_ASAP7_75t_SL g26611 (.A(n_5575),
    .B(n_11763),
    .Y(n_18838));
 XNOR2x1_ASAP7_75t_SL g26612 (.B(n_12540),
    .Y(n_18839),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_583));
 XOR2x2_ASAP7_75t_SL g26615 (.A(n_15581),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_737),
    .Y(n_18842));
 XNOR2x2_ASAP7_75t_SL g26616 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_169),
    .B(n_5645),
    .Y(n_18843));
 XOR2xp5_ASAP7_75t_SL g26619 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_116),
    .Y(n_18846));
 XOR2xp5_ASAP7_75t_SL g26621 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_43),
    .Y(n_18848));
 XOR2xp5_ASAP7_75t_SL g26622 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_10),
    .Y(n_18849));
 XNOR2xp5_ASAP7_75t_SL g26623 (.A(n_5886),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_107),
    .Y(n_18850));
 XNOR2xp5_ASAP7_75t_SL g26624 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_673),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_577),
    .Y(n_18851));
 XNOR2x1_ASAP7_75t_SL g26629 (.B(n_18857),
    .Y(n_18856),
    .A(n_10509));
 XOR2xp5_ASAP7_75t_SL g26630 (.A(n_23391),
    .B(n_8474),
    .Y(n_18857));
 XOR2xp5_ASAP7_75t_SL g26631 (.A(n_6238),
    .B(n_6125),
    .Y(n_18858));
 XOR2xp5_ASAP7_75t_SL g26635 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_751),
    .B(n_19020),
    .Y(n_18862));
 XNOR2x1_ASAP7_75t_SL g26636 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_137),
    .Y(n_18863),
    .A(n_22190));
 XOR2xp5_ASAP7_75t_SL g26638 (.A(n_7869),
    .B(n_6569),
    .Y(n_18865));
 XNOR2xp5_ASAP7_75t_SL g26639 (.A(n_22634),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_71),
    .Y(n_18866));
 XOR2xp5_ASAP7_75t_SL g26640 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_57),
    .Y(n_18867));
 OR2x2_ASAP7_75t_SL g26641 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_180),
    .B(n_7573),
    .Y(n_18868));
 XOR2xp5_ASAP7_75t_SL g26643 (.A(n_13727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_107),
    .Y(n_18870));
 XOR2x2_ASAP7_75t_SL g26644 (.A(n_18870),
    .B(n_6766),
    .Y(n_18871));
 XNOR2xp5_ASAP7_75t_SL g26647 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_78),
    .Y(n_18874));
 XNOR2x1_ASAP7_75t_SL g26648 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_683),
    .Y(n_18875),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_587));
 XOR2xp5_ASAP7_75t_SL g26654 (.A(n_19441),
    .B(n_9634),
    .Y(n_18881));
 XNOR2xp5_ASAP7_75t_SL g26656 (.A(n_15166),
    .B(n_15167),
    .Y(n_18883));
 XOR2xp5_ASAP7_75t_SL g26657 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_174),
    .B(n_7318),
    .Y(n_18884));
 XNOR2x2_ASAP7_75t_SL g26658 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_57),
    .Y(n_18885));
 XOR2xp5_ASAP7_75t_SL g26659 (.A(n_22631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_71),
    .Y(n_18886));
 XOR2xp5_ASAP7_75t_SL g26662 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_50),
    .B(n_7447),
    .Y(n_18889));
 XOR2xp5_ASAP7_75t_SL g26664 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_278),
    .B(n_11832),
    .Y(n_18891));
 XOR2xp5_ASAP7_75t_SL g26669 (.A(n_11238),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_304),
    .Y(n_18896));
 XOR2xp5_ASAP7_75t_SL g26670 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_73),
    .Y(n_18897));
 XOR2x2_ASAP7_75t_SL g26671 (.A(n_18899),
    .B(n_18900),
    .Y(n_15166));
 XOR2xp5_ASAP7_75t_SL g26672 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_95),
    .B(n_18807),
    .Y(n_18899));
 XOR2xp5_ASAP7_75t_SL g26673 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_17),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_20),
    .Y(n_18900));
 XOR2xp5_ASAP7_75t_SL g26674 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_49),
    .Y(n_18901));
 XOR2xp5_ASAP7_75t_SL g26675 (.A(n_11021),
    .B(n_8158),
    .Y(n_18902));
 XOR2xp5_ASAP7_75t_SL g26676 (.A(n_8248),
    .B(n_19404),
    .Y(n_18903));
 OR2x2_ASAP7_75t_SL g26677 (.A(n_13126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_180),
    .Y(n_18904));
 XNOR2xp5_ASAP7_75t_SL g26680 (.A(n_11189),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_46),
    .Y(n_18907));
 XOR2xp5_ASAP7_75t_SL g26687 (.A(n_8719),
    .B(n_8722),
    .Y(n_18914));
 XOR2xp5_ASAP7_75t_SL g26688 (.A(n_8739),
    .B(n_18997),
    .Y(n_18915));
 XNOR2xp5_ASAP7_75t_SL g26689 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_115),
    .Y(n_18916));
 XOR2xp5_ASAP7_75t_SL g26691 (.A(n_8871),
    .B(n_8878),
    .Y(n_8881));
 XNOR2x1_ASAP7_75t_SL g26692 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_89),
    .Y(n_18919),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_33));
 XNOR2x1_ASAP7_75t_SL g26698 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_29),
    .Y(n_18925),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_9));
 XNOR2xp5_ASAP7_75t_SL g26699 (.A(n_6853),
    .B(n_9313),
    .Y(n_18926));
 INVx1_ASAP7_75t_SL g267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_22),
    .Y(n_6062));
 XOR2x2_ASAP7_75t_SL g26700 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_59),
    .Y(n_18927));
 XOR2xp5_ASAP7_75t_SL g26701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_194),
    .Y(n_18928));
 XOR2xp5_ASAP7_75t_SL g26702 (.A(n_11169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_210),
    .Y(n_18929));
 XOR2xp5_ASAP7_75t_SL g26703 (.A(n_6209),
    .B(n_6211),
    .Y(n_18930));
 XOR2x2_ASAP7_75t_SL g26706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .B(n_20327),
    .Y(n_18933));
 XNOR2xp5_ASAP7_75t_SL g26707 (.A(n_3206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_31),
    .Y(n_18934));
 XOR2xp5_ASAP7_75t_SL g26708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_55),
    .B(n_9842),
    .Y(n_18935));
 XOR2xp5_ASAP7_75t_SL g26711 (.A(n_22525),
    .B(n_22252),
    .Y(n_18938));
 XNOR2xp5_ASAP7_75t_SL g26712 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_49),
    .B(n_10947),
    .Y(n_18939));
 MAJx2_ASAP7_75t_SL g26713 (.A(n_19649),
    .B(n_19647),
    .C(n_19648),
    .Y(n_18940));
 XNOR2xp5_ASAP7_75t_SL g26714 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_86),
    .Y(n_18941));
 XOR2x2_ASAP7_75t_SL g26715 (.A(n_10100),
    .B(n_18943),
    .Y(n_18942));
 XOR2xp5_ASAP7_75t_SL g26716 (.A(n_7862),
    .B(n_7863),
    .Y(n_18943));
 XOR2xp5_ASAP7_75t_SL g26718 (.A(n_9740),
    .B(n_9739),
    .Y(n_18945));
 XNOR2xp5_ASAP7_75t_SL g26719 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_148),
    .Y(n_10157));
 XOR2xp5_ASAP7_75t_SL g26720 (.A(n_14092),
    .B(n_10163),
    .Y(n_18947));
 OR2x2_ASAP7_75t_SL g26721 (.A(n_9617),
    .B(n_9618),
    .Y(n_18948));
 XNOR2xp5_ASAP7_75t_SL g26722 (.A(n_22881),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_86),
    .Y(n_18949));
 XOR2xp5_ASAP7_75t_SL g26725 (.A(n_10224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_149),
    .Y(n_18952));
 XNOR2xp5_ASAP7_75t_SL g26726 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_40),
    .B(n_10344),
    .Y(n_18953));
 MAJx2_ASAP7_75t_SL g26727 (.A(n_2903),
    .B(n_22974),
    .C(n_19050),
    .Y(n_18954));
 XOR2x2_ASAP7_75t_SL g26729 (.A(n_14698),
    .B(n_9541),
    .Y(n_18956));
 XOR2xp5_ASAP7_75t_SL g26730 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_132),
    .B(n_10788),
    .Y(n_18957));
 XNOR2xp5_ASAP7_75t_SL g26731 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_25),
    .Y(n_10788));
 XOR2xp5_ASAP7_75t_SL g26733 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_20),
    .B(n_10878),
    .Y(n_18960));
 XNOR2xp5_ASAP7_75t_SL g26734 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_65),
    .Y(n_18961));
 XNOR2x1_ASAP7_75t_L g26737 (.B(n_6668),
    .Y(n_18964),
    .A(n_6667));
 XOR2xp5_ASAP7_75t_SL g26740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_74),
    .B(n_22884),
    .Y(n_18967));
 XOR2xp5_ASAP7_75t_SL g26741 (.A(n_5826),
    .B(n_9069),
    .Y(n_18968));
 XNOR2xp5_ASAP7_75t_SL g26742 (.A(n_11204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_136),
    .Y(n_18969));
 XOR2xp5_ASAP7_75t_SL g26743 (.A(n_11220),
    .B(n_14864),
    .Y(n_18970));
 XNOR2xp5_ASAP7_75t_SL g26745 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_64),
    .Y(n_18972));
 XNOR2xp5_ASAP7_75t_SL g26746 (.A(n_23433),
    .B(n_10188),
    .Y(n_18973));
 XOR2xp5_ASAP7_75t_SL g26747 (.A(n_11529),
    .B(n_13100),
    .Y(n_18974));
 XOR2xp5_ASAP7_75t_SL g26751 (.A(n_12425),
    .B(n_12427),
    .Y(n_18978));
 OR2x2_ASAP7_75t_SL g26756 (.A(n_7029),
    .B(n_7027),
    .Y(n_18983));
 XOR2xp5_ASAP7_75t_SL g26758 (.A(n_12420),
    .B(n_12422),
    .Y(n_18985));
 XNOR2xp5_ASAP7_75t_SL g26759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_99),
    .Y(n_18986));
 XOR2x1_ASAP7_75t_SL g26760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_150),
    .Y(n_18987),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_116));
 XOR2xp5_ASAP7_75t_SL g26761 (.A(n_18987),
    .B(n_23002),
    .Y(n_18988));
 XNOR2xp5_ASAP7_75t_SL g26765 (.A(n_22068),
    .B(n_12712),
    .Y(n_18992));
 XNOR2xp5_ASAP7_75t_SL g26766 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_150),
    .B(n_20235),
    .Y(n_18993));
 XNOR2xp5_ASAP7_75t_SL g26769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_785),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_561),
    .Y(n_18996));
 XNOR2xp5_ASAP7_75t_SL g26770 (.A(n_12905),
    .B(n_12906),
    .Y(n_18997));
 XNOR2xp5_ASAP7_75t_SL g26772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_184),
    .Y(n_18999));
 XOR2xp5_ASAP7_75t_SL g26773 (.A(n_12938),
    .B(n_12945),
    .Y(n_12948));
 XNOR2x1_ASAP7_75t_SL g26774 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_89),
    .Y(n_19001),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_33));
 XOR2x2_ASAP7_75t_SL g26775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_163),
    .Y(n_19002));
 XOR2xp5_ASAP7_75t_SL g26779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_195),
    .Y(n_19006));
 XOR2xp5_ASAP7_75t_SL g26780 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_71),
    .B(n_13133),
    .Y(n_19007));
 XOR2xp5_ASAP7_75t_SL g26781 (.A(n_13144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_54),
    .Y(n_19008));
 XOR2xp5_ASAP7_75t_SL g26784 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_273),
    .Y(n_19011));
 XOR2xp5_ASAP7_75t_SL g26785 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_757),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .Y(n_19012));
 OR2x2_ASAP7_75t_SL g26786 (.A(n_19193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_189),
    .Y(n_19013));
 XNOR2xp5_ASAP7_75t_SL g26787 (.A(n_8241),
    .B(n_13416),
    .Y(n_19014));
 XOR2xp5_ASAP7_75t_SL g26788 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_191),
    .Y(n_19015));
 XNOR2xp5_ASAP7_75t_SL g26789 (.A(n_12428),
    .B(n_15922),
    .Y(n_19016));
 XNOR2xp5_ASAP7_75t_SL g26790 (.A(n_25605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_293),
    .Y(n_19017));
 XNOR2xp5_ASAP7_75t_SL g26791 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_661),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_629),
    .Y(n_19018));
 OR2x2_ASAP7_75t_SL g26792 (.A(n_10758),
    .B(n_22188),
    .Y(n_19019));
 XNOR2xp5_ASAP7_75t_SL g26793 (.A(n_13960),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_687),
    .Y(n_19020));
 OR2x2_ASAP7_75t_SL g26794 (.A(n_21577),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_293),
    .Y(n_19021));
 XOR2xp5_ASAP7_75t_SL g26795 (.A(n_14033),
    .B(n_14035),
    .Y(n_19022));
 XNOR2xp5_ASAP7_75t_SL g26796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_34),
    .Y(n_19023));
 XOR2xp5_ASAP7_75t_SL g26797 (.A(n_14048),
    .B(n_14050),
    .Y(n_19024));
 XNOR2x1_ASAP7_75t_SL g268 (.B(n_6923),
    .Y(n_6924),
    .A(n_10471));
 XNOR2xp5_ASAP7_75t_SL g26800 (.A(n_14237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_112),
    .Y(n_19027));
 XNOR2xp5_ASAP7_75t_SL g26801 (.A(n_9628),
    .B(n_22626),
    .Y(n_19028));
 XOR2xp5_ASAP7_75t_SL g26802 (.A(n_19028),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_80),
    .Y(n_19029));
 XNOR2xp5_ASAP7_75t_SL g26805 (.A(n_13776),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_101),
    .Y(n_19032));
 XOR2xp5_ASAP7_75t_SL g26806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_34),
    .Y(n_19033));
 XNOR2xp5_ASAP7_75t_SL g26807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .Y(n_19034));
 XOR2xp5_ASAP7_75t_SL g26808 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_43),
    .Y(n_19035));
 XOR2xp5_ASAP7_75t_SL g26809 (.A(n_16349),
    .B(n_14878),
    .Y(n_19036));
 XNOR2xp5_ASAP7_75t_SL g26810 (.A(n_14915),
    .B(n_19038),
    .Y(n_19037));
 XOR2xp5_ASAP7_75t_SL g26811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_171),
    .Y(n_19038));
 XOR2xp5_ASAP7_75t_SL g26812 (.A(n_14920),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_270),
    .Y(n_19039));
 XNOR2xp5_ASAP7_75t_SL g26814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_58),
    .Y(n_19041));
 XNOR2x1_ASAP7_75t_SL g26816 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_659),
    .Y(n_19043),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_627));
 XNOR2xp5_ASAP7_75t_SL g26817 (.A(n_12896),
    .B(n_12897),
    .Y(n_19044));
 XOR2xp5_ASAP7_75t_SL g26818 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_42),
    .Y(n_19045));
 XNOR2xp5_ASAP7_75t_SL g26822 (.A(n_9407),
    .B(n_9408),
    .Y(n_19049));
 XOR2x2_ASAP7_75t_SL g26823 (.A(n_18063),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_275),
    .Y(n_19050));
 INVx1_ASAP7_75t_SL g26825 (.A(n_19052),
    .Y(n_19053));
 OAI32xp33_ASAP7_75t_SL g26826 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_117),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_80),
    .B1(n_9375),
    .B2(n_9376),
    .Y(n_19052));
 AND3x1_ASAP7_75t_SL g26827 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_20464),
    .C(n_22164),
    .Y(n_19054));
 AND3x1_ASAP7_75t_SL g26828 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_20464),
    .C(n_12748),
    .Y(n_19055));
 AND3x1_ASAP7_75t_SL g26829 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_2525),
    .C(n_13030),
    .Y(n_19056));
 AND3x1_ASAP7_75t_SL g26830 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_2525),
    .C(n_20825),
    .Y(n_19057));
 AND3x1_ASAP7_75t_SL g26831 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_2945),
    .C(n_2160),
    .Y(n_19058));
 AND3x1_ASAP7_75t_SL g26832 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_20464),
    .C(n_2168),
    .Y(n_19059));
 AND3x1_ASAP7_75t_SL g26833 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(n_2525),
    .C(n_19370),
    .Y(n_19060));
 AND3x1_ASAP7_75t_SL g26834 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_2945),
    .C(n_2162),
    .Y(n_19061));
 AND3x1_ASAP7_75t_SL g26835 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_2945),
    .C(n_2165),
    .Y(n_19062));
 AND3x1_ASAP7_75t_SL g26836 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_20464),
    .C(n_2159),
    .Y(n_19063));
 AND3x1_ASAP7_75t_SL g26837 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(n_2525),
    .C(n_12781),
    .Y(n_19064));
 AND3x1_ASAP7_75t_SL g26838 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_2944),
    .C(n_19838),
    .Y(n_19065));
 FAx1_ASAP7_75t_SL g26840 (.SN(n_19067),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .B(n_19069),
    .CI(n_19071),
    .CON(UNCONNECTED));
 FAx1_ASAP7_75t_SL g26841 (.SN(n_19068),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .CON(UNCONNECTED0));
 FAx1_ASAP7_75t_SL g26842 (.SN(n_19069),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_671),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_799),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_n_639),
    .CON(UNCONNECTED1));
 FAx1_ASAP7_75t_SL g26843 (.SN(n_19070),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_573),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_n_701),
    .CON(UNCONNECTED2));
 FAx1_ASAP7_75t_SL g26844 (.SN(n_19071),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_767),
    .B(n_19064),
    .CI(n_19065),
    .CON(UNCONNECTED3));
 AO21x1_ASAP7_75t_SL g26845 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_91),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_144),
    .Y(n_19072));
 AO21x1_ASAP7_75t_SL g26846 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_142),
    .Y(n_19073));
 AO21x1_ASAP7_75t_SL g26848 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_168),
    .Y(n_19075));
 AO21x1_ASAP7_75t_SL g26849 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_51),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_164),
    .Y(n_19076));
 FAx1_ASAP7_75t_SL g26850 (.SN(n_19077),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_157),
    .CON(UNCONNECTED4));
 AO21x1_ASAP7_75t_SL g26851 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_49),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_162),
    .Y(n_19078));
 FAx1_ASAP7_75t_SL g26852 (.SN(n_19079),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_96),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_159),
    .CON(UNCONNECTED5));
 AO21x1_ASAP7_75t_SL g26853 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_168),
    .Y(n_19080));
 FAx1_ASAP7_75t_SL g26856 (.SN(n_19083),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .B(n_19084),
    .CI(n_26181),
    .CON(UNCONNECTED6));
 FAx1_ASAP7_75t_SL g26857 (.SN(n_19084),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_671),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_799),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_n_639),
    .CON(UNCONNECTED7));
 AO21x1_ASAP7_75t_SL g26858 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_91),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_144),
    .Y(n_19085));
 OAI21xp33_ASAP7_75t_SL g26859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_181),
    .A2(n_21210),
    .B(n_9883),
    .Y(n_19086));
 AO21x1_ASAP7_75t_SL g26861 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_142),
    .Y(n_19088));
 AO21x1_ASAP7_75t_SL g26862 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_168),
    .Y(n_19089));
 FAx1_ASAP7_75t_SL g26863 (.SN(n_19090),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_157),
    .CON(UNCONNECTED8));
 AO21x1_ASAP7_75t_SL g26864 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_49),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_162),
    .Y(n_19091));
 AO21x1_ASAP7_75t_SL g26866 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_142),
    .A2(n_13250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_167),
    .Y(n_19093));
 FAx1_ASAP7_75t_SL g26868 (.SN(n_19095),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .B(n_19097),
    .CI(n_19098),
    .CON(UNCONNECTED9));
 FAx1_ASAP7_75t_SL g26869 (.SN(n_19096),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .CON(UNCONNECTED10));
 FAx1_ASAP7_75t_SL g26870 (.SN(n_19097),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_671),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_799),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_n_639),
    .CON(UNCONNECTED11));
 FAx1_ASAP7_75t_SL g26871 (.SN(n_19098),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_767),
    .B(n_19060),
    .CI(n_19061),
    .CON(UNCONNECTED12));
 AO21x1_ASAP7_75t_SL g26872 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_91),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_144),
    .Y(n_19099));
 AO21x1_ASAP7_75t_SL g26874 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_142),
    .Y(n_19101));
 AO21x1_ASAP7_75t_SL g26875 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_168),
    .Y(n_19102));
 FAx1_ASAP7_75t_SL g26876 (.SN(n_19103),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_38),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_87),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_159),
    .CON(UNCONNECTED13));
 AO21x1_ASAP7_75t_SL g26877 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_51),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_164),
    .Y(n_19104));
 FAx1_ASAP7_75t_SL g26878 (.SN(n_19105),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_157),
    .CON(UNCONNECTED14));
 AO21x1_ASAP7_75t_SL g26879 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_49),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_162),
    .Y(n_19106));
 AO21x1_ASAP7_75t_SL g26881 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_168),
    .Y(n_19108));
 AO21x1_ASAP7_75t_SL g26882 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_142),
    .A2(n_13251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_167),
    .Y(n_19109));
 FAx1_ASAP7_75t_SL g26884 (.SN(n_19111),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .B(n_19113),
    .CI(n_19114),
    .CON(UNCONNECTED15));
 FAx1_ASAP7_75t_SL g26885 (.SN(n_19112),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .CON(UNCONNECTED16));
 FAx1_ASAP7_75t_SL g26886 (.SN(n_19113),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_671),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_799),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_n_639),
    .CON(UNCONNECTED17));
 FAx1_ASAP7_75t_SL g26887 (.SN(n_19114),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_767),
    .B(n_19056),
    .CI(n_19062),
    .CON(UNCONNECTED18));
 AO21x1_ASAP7_75t_SL g26888 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_91),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_144),
    .Y(n_19115));
 AO21x1_ASAP7_75t_SL g26890 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_142),
    .Y(n_19117));
 AO21x1_ASAP7_75t_SL g26893 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_51),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_164),
    .Y(n_19120));
 AO21x1_ASAP7_75t_SL g26895 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_49),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_162),
    .Y(n_19122));
 FAx1_ASAP7_75t_SL g26896 (.SN(n_19123),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_96),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_159),
    .CON(UNCONNECTED19));
 AO21x1_ASAP7_75t_SL g26897 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_139),
    .B(n_8974),
    .Y(n_19124));
 OAI22xp5_ASAP7_75t_SL g26899 (.A1(n_4031),
    .A2(n_5602),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_69),
    .B2(n_13723),
    .Y(n_19126));
 MAJIxp5_ASAP7_75t_SL g269 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_212),
    .B(n_6928),
    .C(n_6929),
    .Y(n_6930));
 AND3x1_ASAP7_75t_SL g26901 (.A(n_6144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_84),
    .Y(n_19128));
 XNOR2xp5_ASAP7_75t_SL g26902 (.A(n_6371),
    .B(n_18700),
    .Y(n_19129));
 MAJIxp5_ASAP7_75t_SL g26904 (.A(n_5536),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_115),
    .C(n_6439),
    .Y(n_19131));
 AOI21xp33_ASAP7_75t_SL g26905 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_274),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_270),
    .B(n_19734),
    .Y(n_19132));
 OAI21xp33_ASAP7_75t_SL g26906 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_181),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_214),
    .B(n_6655),
    .Y(n_19133));
 MAJx2_ASAP7_75t_SL g26907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_131),
    .C(n_6741),
    .Y(n_19134));
 MAJx2_ASAP7_75t_SL g26908 (.A(n_6754),
    .B(n_11361),
    .C(n_6751),
    .Y(n_19135));
 XNOR2xp5_ASAP7_75t_SL g26909 (.A(n_6862),
    .B(n_18710),
    .Y(n_19136));
 XNOR2xp5_ASAP7_75t_SL g26910 (.A(n_18719),
    .B(n_6894),
    .Y(n_19137));
 OAI22xp5_ASAP7_75t_SL g26911 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_73),
    .A2(n_6967),
    .B1(n_6969),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_72),
    .Y(n_19138));
 OAI22xp5_ASAP7_75t_SL g26914 (.A1(n_7082),
    .A2(n_3770),
    .B1(n_8836),
    .B2(n_8838),
    .Y(n_19141));
 OAI21xp33_ASAP7_75t_SL g26915 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_188),
    .A2(n_21462),
    .B(n_7169),
    .Y(n_19142));
 MAJx2_ASAP7_75t_SL g26916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_89),
    .B(n_15552),
    .C(n_9441),
    .Y(n_19143));
 XOR2xp5_ASAP7_75t_SL g26917 (.A(n_7256),
    .B(n_7257),
    .Y(n_19144));
 XNOR2xp5_ASAP7_75t_SL g26918 (.A(n_19531),
    .B(n_19207),
    .Y(n_19145));
 NOR3xp33_ASAP7_75t_SL g26919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_119),
    .C(n_2718),
    .Y(n_19146));
 OAI21xp33_ASAP7_75t_SL g26920 (.A1(n_19201),
    .A2(n_15185),
    .B(n_15187),
    .Y(n_19147));
 MAJIxp5_ASAP7_75t_SL g26921 (.A(n_4515),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_108),
    .C(n_19764),
    .Y(n_8573));
 MAJIxp5_ASAP7_75t_SL g26922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .Y(n_19149));
 MAJIxp5_ASAP7_75t_SL g26923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_759),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_631),
    .Y(n_19150));
 MAJIxp5_ASAP7_75t_SL g26927 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_26),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_62),
    .Y(n_12252));
 XNOR2xp5_ASAP7_75t_SL g26933 (.A(n_10122),
    .B(n_18707),
    .Y(n_19160));
 OAI21xp5_ASAP7_75t_SL g26937 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_99),
    .B(n_10073),
    .Y(n_19164));
 MAJIxp5_ASAP7_75t_SL g26938 (.A(n_10125),
    .B(n_18707),
    .C(n_9747),
    .Y(n_19165));
 XNOR2xp5_ASAP7_75t_SL g26941 (.A(n_10718),
    .B(n_10350),
    .Y(n_19168));
 MAJIxp5_ASAP7_75t_SL g26942 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_147),
    .B(n_15386),
    .C(n_10466),
    .Y(n_19169));
 OA211x2_ASAP7_75t_SL g26943 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_n_753),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_3),
    .B(n_10503),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_145),
    .Y(n_19170));
 XNOR2xp5_ASAP7_75t_SL g26944 (.A(n_10516),
    .B(n_18732),
    .Y(n_10520));
 XOR2xp5_ASAP7_75t_SL g26945 (.A(n_10635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_4),
    .Y(n_19172));
 OAI21xp5_ASAP7_75t_SL g26947 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_193),
    .B(n_2180),
    .Y(n_19174));
 OA211x2_ASAP7_75t_SL g26948 (.A1(n_11000),
    .A2(n_10902),
    .B(n_9503),
    .C(n_11872),
    .Y(n_19175));
 XNOR2xp5_ASAP7_75t_SL g26950 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_156),
    .B(n_11054),
    .Y(n_19177));
 XNOR2xp5_ASAP7_75t_SL g26954 (.A(n_18781),
    .B(n_18701),
    .Y(n_19181));
 OAI32xp33_ASAP7_75t_SL g26955 (.A1(n_9209),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_297),
    .A3(n_11480),
    .B1(n_12276),
    .B2(n_11481),
    .Y(n_19182));
 OAI21xp33_ASAP7_75t_SL g26956 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_17),
    .Y(n_19183));
 MAJIxp5_ASAP7_75t_SL g26958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_147),
    .C(n_12929),
    .Y(n_19185));
 MAJIxp5_ASAP7_75t_SL g26959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .Y(n_19186));
 XNOR2xp5_ASAP7_75t_SL g26960 (.A(n_12814),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .Y(n_19187));
 MAJIxp5_ASAP7_75t_SL g26961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_759),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_131),
    .Y(n_19188));
 MAJIxp5_ASAP7_75t_SL g26962 (.A(n_3963),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_190),
    .C(n_20314),
    .Y(n_19189));
 MAJx2_ASAP7_75t_SL g26963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_73),
    .C(n_15158),
    .Y(n_19190));
 MAJx2_ASAP7_75t_SL g26964 (.A(n_19444),
    .B(n_18726),
    .C(n_5988),
    .Y(n_19191));
 OAI21xp5_ASAP7_75t_SL g26966 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_65),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_167),
    .B(n_13030),
    .Y(n_19193));
 A2O1A1Ixp33_ASAP7_75t_SL g26967 (.A1(n_16557),
    .A2(n_9182),
    .B(n_9259),
    .C(n_8014),
    .Y(n_19194));
 XNOR2xp5_ASAP7_75t_SL g26968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_200),
    .B(n_22232),
    .Y(n_19195));
 XOR2xp5_ASAP7_75t_SL g26970 (.A(n_14153),
    .B(n_14158),
    .Y(n_19197));
 XNOR2xp5_ASAP7_75t_SL g26972 (.A(n_14815),
    .B(n_18799),
    .Y(n_19199));
 MAJIxp5_ASAP7_75t_SL g26973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_43),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_88),
    .C(n_14857),
    .Y(n_19200));
 MAJIxp5_ASAP7_75t_SL g26974 (.A(n_18091),
    .B(n_15171),
    .C(n_3729),
    .Y(n_19201));
 OAI22xp5_ASAP7_75t_SL g26978 (.A1(n_17651),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .B2(n_11550),
    .Y(n_19205));
 XNOR2xp5_ASAP7_75t_SL g26979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_133),
    .B(n_18175),
    .Y(n_19206));
 OA21x2_ASAP7_75t_SL g26980 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_254),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_14),
    .B(n_19534),
    .Y(n_19207));
 XOR2xp5_ASAP7_75t_SL g26981 (.A(n_11361),
    .B(n_6751),
    .Y(n_19208));
 AOI21xp5_ASAP7_75t_SL g26991 (.A1(n_19218),
    .A2(n_8626),
    .B(n_8638),
    .Y(n_19219));
 XOR2xp5_ASAP7_75t_SL g26992 (.A(n_8631),
    .B(n_22815),
    .Y(n_19218));
 XOR2x1_ASAP7_75t_SL g26996 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_148),
    .Y(n_19222),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_161));
 AO21x2_ASAP7_75t_SL g27 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_266),
    .A2(n_8304),
    .B(n_20077),
    .Y(n_20078));
 AOI21xp5_ASAP7_75t_SL g27001 (.A1(n_7906),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_217),
    .B(n_19228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_73));
 OAI21xp33_ASAP7_75t_SL g27002 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_70),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_191),
    .B(n_9661),
    .Y(n_19228));
 OAI21xp5_ASAP7_75t_SL g27004 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_70),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_191),
    .B(n_2179),
    .Y(n_19230));
 OAI21xp5_ASAP7_75t_SL g27006 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_193),
    .B(n_9662),
    .Y(n_19232));
 XOR2xp5_ASAP7_75t_SL g27007 (.A(n_19234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_220),
    .Y(n_19235));
 XOR2xp5_ASAP7_75t_SL g27008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_154),
    .Y(n_19234));
 HAxp5_ASAP7_75t_SL g27009 (.A(u_NV_NVDLA_cmac_dp2reg_done),
    .B(u_NV_NVDLA_cmac_u_reg_dp2reg_consumer),
    .CON(n_19237),
    .SN(n_19236));
 HAxp5_ASAP7_75t_SL g27011 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_266),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_265),
    .CON(n_19241),
    .SN(n_19240));
 HAxp5_ASAP7_75t_SL g27012 (.A(n_9202),
    .B(n_8145),
    .CON(n_19242),
    .SN(n_19243));
 NAND2xp5_ASAP7_75t_SL g27014 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(n_5529));
 MAJIxp5_ASAP7_75t_SL g27017 (.A(n_19248),
    .B(n_9860),
    .C(n_9862),
    .Y(n_19249));
 MAJx2_ASAP7_75t_SL g27018 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_140),
    .Y(n_19248));
 MAJIxp5_ASAP7_75t_SL g27021 (.A(n_19252),
    .B(n_19516),
    .C(n_26102),
    .Y(n_19253));
 NOR2xp67_ASAP7_75t_SL g27023 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_258),
    .B(n_23169),
    .Y(n_19254));
 XNOR2xp5_ASAP7_75t_SL g27028 (.A(n_19259),
    .B(n_24670),
    .Y(n_19261));
 AND2x2_ASAP7_75t_SL g27029 (.A(n_12975),
    .B(n_12978),
    .Y(n_19259));
 OAI21xp5_ASAP7_75t_SL g27031 (.A1(n_19263),
    .A2(n_10240),
    .B(n_10243),
    .Y(n_19264));
 AO21x1_ASAP7_75t_SL g27033 (.A1(n_12107),
    .A2(n_19263),
    .B(n_12108),
    .Y(n_19265));
 XNOR2xp5_ASAP7_75t_SL g27035 (.A(n_14064),
    .B(n_19269),
    .Y(n_19270));
 XNOR2xp5_ASAP7_75t_SL g27036 (.A(n_19267),
    .B(n_19268),
    .Y(n_19269));
 MAJIxp5_ASAP7_75t_SL g27037 (.A(n_21212),
    .B(n_9434),
    .C(n_18597),
    .Y(n_19267));
 MAJIxp5_ASAP7_75t_SL g27038 (.A(n_14064),
    .B(n_19271),
    .C(n_19272),
    .Y(n_19273));
 INVxp67_ASAP7_75t_SRAM g27039 (.A(n_19268),
    .Y(n_19271));
 HB1xp67_ASAP7_75t_SL g27040 (.A(n_19267),
    .Y(n_19272));
 HB1xp67_ASAP7_75t_SL g27053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_63),
    .Y(n_19304));
 NAND2x1_ASAP7_75t_SL g27056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109),
    .B(n_19305),
    .Y(n_19306));
 OR2x2_ASAP7_75t_SL g27057 (.A(n_13936),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_67),
    .Y(n_19305));
 MAJx2_ASAP7_75t_SL g27058 (.A(n_19307),
    .B(n_19308),
    .C(n_19309),
    .Y(n_19310));
 INVx1_ASAP7_75t_SL g27059 (.A(n_10421),
    .Y(n_19308));
 INVx1_ASAP7_75t_SL g27060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_63),
    .Y(n_19309));
 XOR2xp5_ASAP7_75t_SL g27068 (.A(n_20810),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_199),
    .Y(n_19323));
 MAJIxp5_ASAP7_75t_SL g27069 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_167),
    .B(n_8019),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_185),
    .Y(n_19324));
 HB1xp67_ASAP7_75t_SL g27070 (.A(n_19326),
    .Y(n_19327));
 XNOR2xp5_ASAP7_75t_SL g27071 (.A(n_22854),
    .B(n_23408),
    .Y(n_19330));
 AOI21xp5_ASAP7_75t_SL g27072 (.A1(n_19332),
    .A2(n_19336),
    .B(n_19338),
    .Y(n_19339));
 XNOR2xp5_ASAP7_75t_SL g27073 (.A(n_19331),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_15),
    .Y(n_19332));
 HB1xp67_ASAP7_75t_SL g27074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_33),
    .Y(n_19331));
 NAND2xp33_ASAP7_75t_SL g27075 (.A(n_19334),
    .B(n_19335),
    .Y(n_19336));
 INVxp33_ASAP7_75t_SL g27076 (.A(n_19333),
    .Y(n_19334));
 XNOR2x1_ASAP7_75t_SL g27077 (.B(n_10389),
    .Y(n_19333),
    .A(n_20297));
 MAJIxp5_ASAP7_75t_SL g27078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_140),
    .C(n_6795),
    .Y(n_19335));
 NOR2xp33_ASAP7_75t_SL g27079 (.A(n_19337),
    .B(n_19335),
    .Y(n_19338));
 INVx1_ASAP7_75t_SL g27080 (.A(n_19333),
    .Y(n_19337));
 NAND2xp67_ASAP7_75t_SL g27081 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .B(n_19340),
    .Y(n_19341));
 OAI21x1_ASAP7_75t_SL g27091 (.A1(n_19356),
    .A2(n_19358),
    .B(n_19359),
    .Y(n_19360));
 AND2x2_ASAP7_75t_SL g27092 (.A(n_19353),
    .B(n_19355),
    .Y(n_19356));
 XNOR2x2_ASAP7_75t_SL g27093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_20),
    .Y(n_19353));
 MAJIxp5_ASAP7_75t_SL g27094 (.A(n_7079),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_103),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_78),
    .Y(n_19354));
 XNOR2x1_ASAP7_75t_SL g27095 (.B(n_7681),
    .Y(n_19358),
    .A(n_19357));
 OR2x2_ASAP7_75t_SL g27097 (.A(n_19353),
    .B(n_19355),
    .Y(n_19359));
 XNOR2xp5_ASAP7_75t_SL g27099 (.A(n_19365),
    .B(n_19366),
    .Y(n_19367));
 XNOR2x1_ASAP7_75t_SL g27100 (.B(n_19363),
    .Y(n_19365),
    .A(n_26066));
 MAJx2_ASAP7_75t_SL g27103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_116),
    .C(n_7686),
    .Y(n_19363));
 NAND2x1_ASAP7_75t_SL g27104 (.A(n_19372),
    .B(n_19375),
    .Y(n_19376));
 AOI21xp5_ASAP7_75t_SL g27105 (.A1(n_19369),
    .A2(n_16563),
    .B(n_19371),
    .Y(n_19372));
 AND2x2_ASAP7_75t_SL g27106 (.A(n_19368),
    .B(n_16565),
    .Y(n_19369));
 OAI21xp5_ASAP7_75t_SL g27107 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_65),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_189),
    .Y(n_19368));
 OAI21xp5_ASAP7_75t_SL g27108 (.A1(n_19368),
    .A2(n_16565),
    .B(n_19370),
    .Y(n_19371));
 AND3x2_ASAP7_75t_L g27109 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[2]),
    .Y(n_19370));
 AOI22xp33_ASAP7_75t_SL g27110 (.A1(n_10136),
    .A2(n_19374),
    .B1(n_16564),
    .B2(n_19369),
    .Y(n_19375));
 NOR2xp33_ASAP7_75t_SL g27111 (.A(n_19368),
    .B(n_16563),
    .Y(n_19374));
 NAND3xp33_ASAP7_75t_SL g27112 (.A(n_19377),
    .B(n_19378),
    .C(n_10475),
    .Y(n_19380));
 NAND2x1_ASAP7_75t_SL g27113 (.A(n_12667),
    .B(n_12669),
    .Y(n_19377));
 OR2x2_ASAP7_75t_SL g27114 (.A(n_12672),
    .B(n_12674),
    .Y(n_19378));
 OA22x2_ASAP7_75t_SL g27115 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263),
    .B1(n_10533),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_264),
    .Y(n_10475));
 NOR2x1_ASAP7_75t_SL g27116 (.A(n_10533),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_264),
    .Y(n_19381));
 NOR2x1_ASAP7_75t_SL g27117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263),
    .Y(n_19382));
 INVxp67_ASAP7_75t_SL g27121 (.A(n_21988),
    .Y(n_19385));
 MAJIxp5_ASAP7_75t_SL g27123 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_42),
    .Y(n_19386));
 XNOR2xp5_ASAP7_75t_SL g27127 (.A(n_19398),
    .B(n_26097),
    .Y(n_19404));
 XOR2xp5_ASAP7_75t_SL g27128 (.A(n_9917),
    .B(n_10567),
    .Y(n_19398));
 XNOR2xp5_ASAP7_75t_SL g27132 (.A(n_11193),
    .B(n_8530),
    .Y(n_19400));
 AND2x2_ASAP7_75t_SL g27137 (.A(n_22019),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .Y(n_19407));
 NOR2x1p5_ASAP7_75t_SL g27139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_43),
    .B(n_4550),
    .Y(n_19408));
 XNOR2xp5_ASAP7_75t_SL g27154 (.A(n_19428),
    .B(n_19431),
    .Y(n_19432));
 MAJIxp5_ASAP7_75t_SL g27155 (.A(n_14643),
    .B(n_19553),
    .C(n_8283),
    .Y(n_19428));
 XNOR2x1_ASAP7_75t_SL g27156 (.B(n_19430),
    .Y(n_19431),
    .A(n_19429));
 NAND2x1_ASAP7_75t_SL g27157 (.A(n_2180),
    .B(n_11033),
    .Y(n_19429));
 NAND2x1_ASAP7_75t_SL g27158 (.A(n_2176),
    .B(n_7106),
    .Y(n_19430));
 XNOR2xp5_ASAP7_75t_SL g27159 (.A(n_19435),
    .B(n_19440),
    .Y(n_19441));
 OAI22xp5_ASAP7_75t_SL g27160 (.A1(n_19433),
    .A2(n_9797),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113),
    .B2(n_9799),
    .Y(n_19435));
 INVx1_ASAP7_75t_SL g27161 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113),
    .Y(n_19433));
 XNOR2xp5_ASAP7_75t_SL g27163 (.A(n_19437),
    .B(n_19439),
    .Y(n_19440));
 INVxp67_ASAP7_75t_SL g27164 (.A(n_19436),
    .Y(n_19437));
 NAND2xp5_ASAP7_75t_SL g27165 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(n_15192),
    .Y(n_19436));
 AOI21x1_ASAP7_75t_SL g27166 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_52),
    .B(n_19438),
    .Y(n_19439));
 AND2x2_ASAP7_75t_SL g27167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_85),
    .Y(n_19438));
 XOR2xp5_ASAP7_75t_SL g27169 (.A(n_19443),
    .B(n_19444),
    .Y(n_19445));
 XNOR2xp5_ASAP7_75t_SL g27170 (.A(n_18726),
    .B(n_5986),
    .Y(n_19443));
 XNOR2x1_ASAP7_75t_SL g27171 (.B(n_23550),
    .Y(n_19444),
    .A(n_19950));
 XOR2xp5_ASAP7_75t_SL g27172 (.A(n_19446),
    .B(n_19448),
    .Y(n_19449));
 NAND2xp5_ASAP7_75t_SL g27177 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_3374),
    .Y(n_19453));
 NAND2xp5_ASAP7_75t_SL g27178 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_121),
    .Y(n_19454));
 XNOR2xp5_ASAP7_75t_SL g27180 (.A(n_19457),
    .B(n_19461),
    .Y(n_19462));
 INVx1_ASAP7_75t_SL g27181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_131),
    .Y(n_19457));
 XNOR2x1_ASAP7_75t_SL g27190 (.B(n_19471),
    .Y(n_19472),
    .A(n_26100));
 AOI22xp5_ASAP7_75t_SL g27193 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_202),
    .A2(n_4224),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_25),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_190),
    .Y(n_19471));
 MAJx2_ASAP7_75t_SL g27197 (.A(n_23268),
    .B(n_7558),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_83),
    .Y(n_19478));
 INVx1_ASAP7_75t_SL g27199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_78),
    .Y(n_19480));
 XOR2x2_ASAP7_75t_SL g27201 (.A(n_19486),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_224),
    .Y(n_19487));
 XNOR2xp5_ASAP7_75t_SL g27202 (.A(n_6606),
    .B(n_19485),
    .Y(n_19486));
 MAJIxp5_ASAP7_75t_SL g27203 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_182),
    .B(n_21859),
    .C(n_6605),
    .Y(n_19485));
 XNOR2x1_ASAP7_75t_SL g27204 (.B(n_19489),
    .Y(n_19490),
    .A(n_19488));
 MAJx2_ASAP7_75t_SL g27205 (.A(n_10327),
    .B(n_24977),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_186),
    .Y(n_19488));
 XOR2x2_ASAP7_75t_SL g27206 (.A(n_10305),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_9),
    .Y(n_19489));
 XNOR2xp5_ASAP7_75t_SL g27207 (.A(n_19491),
    .B(n_19492),
    .Y(n_19493));
 NAND2xp5_ASAP7_75t_SL g27208 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(n_19491));
 NAND2xp5_ASAP7_75t_SL g27209 (.A(n_14987),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .Y(n_19492));
 INVxp67_ASAP7_75t_SL g27210 (.A(n_19491),
    .Y(n_19494));
 NAND2xp5_ASAP7_75t_SL g27218 (.A(n_19730),
    .B(n_19729),
    .Y(n_19515));
 XNOR2xp5_ASAP7_75t_SL g27221 (.A(n_19517),
    .B(n_26102),
    .Y(n_19522));
 INVx1_ASAP7_75t_SL g27222 (.A(n_19516),
    .Y(n_19517));
 OR2x2_ASAP7_75t_SL g27223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_100),
    .Y(n_19516));
 NOR2xp67_ASAP7_75t_SL g27227 (.A(n_19523),
    .B(n_20239),
    .Y(n_19525));
 XOR2x2_ASAP7_75t_SL g27229 (.A(n_26103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_545),
    .Y(n_19530));
 OA21x2_ASAP7_75t_SL g27235 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_305),
    .Y(n_19531));
 HB1xp67_ASAP7_75t_SL g27236 (.A(n_19532),
    .Y(n_19533));
 NOR2xp33_ASAP7_75t_SL g27237 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_14),
    .Y(n_19532));
 NAND2xp5_ASAP7_75t_SL g27238 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_14),
    .Y(n_19534));
 XOR2xp5_ASAP7_75t_SL g27239 (.A(n_23139),
    .B(n_20288),
    .Y(n_19538));
 OAI21x1_ASAP7_75t_SL g27242 (.A1(n_19539),
    .A2(n_19541),
    .B(n_19542),
    .Y(n_19543));
 INVx1_ASAP7_75t_SL g27243 (.A(n_19540),
    .Y(n_19541));
 OAI21xp5_ASAP7_75t_SL g27244 (.A1(n_4443),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_198),
    .Y(n_19540));
 XNOR2xp5_ASAP7_75t_SL g27251 (.A(n_19550),
    .B(n_19551),
    .Y(n_19552));
 NAND2x1_ASAP7_75t_SL g27252 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_774),
    .B(n_2158),
    .Y(n_19550));
 NAND2x1_ASAP7_75t_SL g27253 (.A(n_18577),
    .B(n_11236),
    .Y(n_19551));
 INVx1_ASAP7_75t_SL g27254 (.A(n_19550),
    .Y(n_19553));
 XNOR2x1_ASAP7_75t_SL g27255 (.B(n_19555),
    .Y(n_19556),
    .A(n_19554));
 OAI21xp5_ASAP7_75t_SL g27256 (.A1(n_12567),
    .A2(n_14327),
    .B(n_14330),
    .Y(n_19554));
 AND2x4_ASAP7_75t_SL g27257 (.A(n_12260),
    .B(n_2158),
    .Y(n_19555));
 XNOR2xp5_ASAP7_75t_SL g27258 (.A(n_19557),
    .B(n_19558),
    .Y(n_19559));
 NAND2x1_ASAP7_75t_SL g27259 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .Y(n_19557));
 NAND2x1_ASAP7_75t_SL g27260 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(n_19558));
 XNOR2x1_ASAP7_75t_SL g27264 (.B(n_19767),
    .Y(n_19566),
    .A(n_19565));
 XNOR2x1_ASAP7_75t_SL g27265 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_93),
    .Y(n_19565),
    .A(n_19564));
 INVx2_ASAP7_75t_SL g27266 (.A(n_19563),
    .Y(n_19564));
 NAND2x1p5_ASAP7_75t_SL g27267 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .B(n_16757),
    .Y(n_19563));
 XNOR2xp5_ASAP7_75t_SL g27268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_30),
    .B(n_19570),
    .Y(n_19571));
 INVx1_ASAP7_75t_SL g27269 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_40),
    .Y(n_19568));
 XNOR2xp5_ASAP7_75t_SL g27270 (.A(n_19573),
    .B(n_26213),
    .Y(n_19575));
 HB1xp67_ASAP7_75t_SL g27271 (.A(n_19572),
    .Y(n_19573));
 OAI21x1_ASAP7_75t_SL g27272 (.A1(n_8321),
    .A2(n_22222),
    .B(n_9263),
    .Y(n_19572));
 XNOR2xp5_ASAP7_75t_SL g27280 (.A(n_19582),
    .B(n_19583),
    .Y(n_19584));
 OAI21xp5_ASAP7_75t_SL g27281 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_191),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_217),
    .Y(n_19582));
 OAI21xp5_ASAP7_75t_SL g27282 (.A1(n_21961),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_288),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_297),
    .Y(n_19583));
 NAND2xp5_ASAP7_75t_SL g27289 (.A(n_22856),
    .B(n_19330),
    .Y(n_19595));
 XNOR2xp5_ASAP7_75t_SL g27290 (.A(n_19597),
    .B(n_19598),
    .Y(n_19599));
 MAJIxp5_ASAP7_75t_SL g27291 (.A(n_14299),
    .B(n_13701),
    .C(n_4245),
    .Y(n_19597));
 XNOR2x1_ASAP7_75t_SL g27292 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_178),
    .Y(n_19598),
    .A(n_7309));
 XNOR2xp5_ASAP7_75t_SL g27294 (.A(n_19602),
    .B(n_19604),
    .Y(n_19605));
 INVx1_ASAP7_75t_SL g27295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_190),
    .Y(n_19601));
 INVxp67_ASAP7_75t_SL g27296 (.A(n_20314),
    .Y(n_19604));
 NOR2xp67_ASAP7_75t_SL g273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_267),
    .B(n_10754),
    .Y(n_19594));
 XOR2xp5_ASAP7_75t_SL g27302 (.A(n_19612),
    .B(n_19613),
    .Y(n_19614));
 NAND2x1_ASAP7_75t_SL g27303 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(n_6861),
    .Y(n_19612));
 NAND2xp5_ASAP7_75t_SL g27304 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .Y(n_19613));
 INVxp67_ASAP7_75t_SL g27305 (.A(n_19613),
    .Y(n_19615));
 XOR2xp5_ASAP7_75t_SL g27310 (.A(n_19622),
    .B(n_10029),
    .Y(n_19625));
 XNOR2xp5_ASAP7_75t_SL g27311 (.A(n_7886),
    .B(n_11088),
    .Y(n_19622));
 NAND2xp5_ASAP7_75t_SL g27327 (.A(n_19645),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .Y(n_19646));
 XNOR2xp5_ASAP7_75t_SL g27331 (.A(n_19650),
    .B(n_26105),
    .Y(n_7925));
 INVxp67_ASAP7_75t_SL g27332 (.A(n_19649),
    .Y(n_19650));
 MAJIxp5_ASAP7_75t_SL g27333 (.A(n_7263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_150),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_146),
    .Y(n_19649));
 XNOR2x1_ASAP7_75t_SL g27335 (.B(n_19656),
    .Y(n_19657),
    .A(n_22794));
 NAND2x1_ASAP7_75t_SL g27337 (.A(n_2179),
    .B(n_14022),
    .Y(n_19656));
 INVx1_ASAP7_75t_SL g27338 (.A(n_19656),
    .Y(n_19658));
 XNOR2xp5_ASAP7_75t_SL g27340 (.A(n_19661),
    .B(n_19662),
    .Y(n_19663));
 HB1xp67_ASAP7_75t_SL g27341 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_115),
    .Y(n_19660));
 XNOR2xp5_ASAP7_75t_SL g27342 (.A(n_19665),
    .B(n_19666),
    .Y(n_19667));
 INVxp67_ASAP7_75t_SL g27343 (.A(n_19664),
    .Y(n_19665));
 MAJIxp5_ASAP7_75t_SL g27344 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_157),
    .B(n_10635),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_4),
    .Y(n_19664));
 OAI22xp5_ASAP7_75t_SL g27345 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_172),
    .A2(n_26168),
    .B1(n_23372),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_173),
    .Y(n_19666));
 INVxp67_ASAP7_75t_SL g27346 (.A(n_19669),
    .Y(n_19670));
 XNOR2xp5_ASAP7_75t_SL g27347 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_128),
    .Y(n_19669));
 MAJIxp5_ASAP7_75t_SL g27349 (.A(n_25999),
    .B(n_19672),
    .C(n_19673),
    .Y(n_19674));
 INVx1_ASAP7_75t_SL g27350 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_89),
    .Y(n_19672));
 XNOR2xp5_ASAP7_75t_SL g27351 (.A(n_12056),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_141),
    .Y(n_19675));
 XOR2xp5_ASAP7_75t_SL g27352 (.A(n_19679),
    .B(n_19680),
    .Y(n_19681));
 NAND2xp5_ASAP7_75t_SL g27353 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .Y(n_19679));
 NAND2x1p5_ASAP7_75t_SL g27354 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(n_14987),
    .Y(n_19680));
 XNOR2xp5_ASAP7_75t_SL g27355 (.A(n_19682),
    .B(n_26005),
    .Y(n_19685));
 NAND2x1_ASAP7_75t_SL g27356 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .B(n_9154),
    .Y(n_19682));
 XNOR2xp5_ASAP7_75t_SL g27359 (.A(n_19686),
    .B(n_21309),
    .Y(n_19688));
 XNOR2xp5_ASAP7_75t_SL g27360 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_4),
    .Y(n_19686));
 NOR2x1p5_ASAP7_75t_SL g27362 (.A(n_21283),
    .B(n_19695),
    .Y(n_19696));
 XOR2x2_ASAP7_75t_SL g27369 (.A(n_26040),
    .B(n_8500),
    .Y(n_19695));
 INVx1_ASAP7_75t_SL g27370 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_115),
    .Y(n_19697));
 INVx1_ASAP7_75t_SL g27371 (.A(n_21045),
    .Y(n_19698));
 NOR2xp33_ASAP7_75t_SL g27372 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_85),
    .Y(n_19699));
 OAI22xp5_ASAP7_75t_SL g27373 (.A1(n_21045),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_115),
    .B1(n_19697),
    .B2(n_19698),
    .Y(n_19701));
 XOR2xp5_ASAP7_75t_SL g27374 (.A(n_19702),
    .B(n_19704),
    .Y(n_19705));
 NAND2xp5_ASAP7_75t_SL g27375 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(n_3504),
    .Y(n_19702));
 INVx1_ASAP7_75t_SL g27376 (.A(n_19703),
    .Y(n_19704));
 NAND2xp5_ASAP7_75t_SL g27377 (.A(n_2307),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .Y(n_19703));
 INVx1_ASAP7_75t_SL g27378 (.A(n_19702),
    .Y(n_19706));
 XNOR2xp5_ASAP7_75t_SL g27379 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_131),
    .B(n_19711),
    .Y(n_19712));
 XOR2xp5_ASAP7_75t_SL g27380 (.A(n_26108),
    .B(n_19710),
    .Y(n_19711));
 INVx1_ASAP7_75t_SL g27384 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_74),
    .Y(n_19710));
 XNOR2x1_ASAP7_75t_SL g27387 (.B(n_19718),
    .Y(n_19719),
    .A(n_26109));
 XNOR2x1_ASAP7_75t_SL g27391 (.B(n_13505),
    .Y(n_19718),
    .A(n_9061));
 AOI22xp5_ASAP7_75t_SL g27395 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_85),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_16),
    .Y(n_19722));
 XNOR2x1_ASAP7_75t_SL g274 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_65),
    .Y(n_9704),
    .A(n_7657));
 NAND2xp5_ASAP7_75t_SL g27402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_273),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_269),
    .Y(n_19729));
 NAND2xp5_ASAP7_75t_SL g27403 (.A(n_12666),
    .B(n_8365),
    .Y(n_19730));
 INVxp33_ASAP7_75t_SRAM g27404 (.A(n_19729),
    .Y(n_19734));
 OAI22xp5_ASAP7_75t_SL g27407 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_135),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_120),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_134),
    .Y(n_19736));
 XNOR2x1_ASAP7_75t_SL g27408 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_91),
    .Y(n_19737),
    .A(n_8148));
 MAJIxp5_ASAP7_75t_SL g27412 (.A(n_20999),
    .B(n_20996),
    .C(n_20998),
    .Y(n_19746));
 XNOR2xp5_ASAP7_75t_SL g27419 (.A(n_19752),
    .B(n_19753),
    .Y(n_19754));
 NAND2xp5_ASAP7_75t_SL g27420 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .Y(n_19752));
 NAND2xp5_ASAP7_75t_SL g27421 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .Y(n_19753));
 AND2x2_ASAP7_75t_SL g27432 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(n_19764));
 NAND2xp33_ASAP7_75t_SL g27433 (.A(n_4275),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(n_4515));
 HB1xp67_ASAP7_75t_SL g27434 (.A(n_15163),
    .Y(n_19767));
 XNOR2x1_ASAP7_75t_SL g27435 (.B(n_19775),
    .Y(n_19776),
    .A(n_19774));
 NAND2x1_ASAP7_75t_SL g27436 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(n_12800),
    .Y(n_19774));
 AND2x2_ASAP7_75t_SL g27437 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .Y(n_19775));
 XNOR2x1_ASAP7_75t_SL g27439 (.B(n_26111),
    .Y(n_19783),
    .A(n_19779));
 XNOR2xp5_ASAP7_75t_SL g27440 (.A(n_19778),
    .B(n_10972),
    .Y(n_19779));
 INVx1_ASAP7_75t_SL g27441 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_136),
    .Y(n_19778));
 AOI21xp5_ASAP7_75t_SL g27445 (.A1(n_19785),
    .A2(n_19787),
    .B(n_19789),
    .Y(n_19790));
 XNOR2x1_ASAP7_75t_SL g27453 (.B(n_19795),
    .Y(n_19796),
    .A(n_26215));
 INVxp67_ASAP7_75t_SL g27455 (.A(n_21855),
    .Y(n_19795));
 XNOR2x1_ASAP7_75t_SL g27457 (.B(n_19801),
    .Y(n_19802),
    .A(n_19799));
 OAI22xp5_ASAP7_75t_SL g27458 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_23),
    .B1(n_19797),
    .B2(n_12281),
    .Y(n_19799));
 INVx1_ASAP7_75t_SL g27459 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_23),
    .Y(n_19797));
 XNOR2x1_ASAP7_75t_SL g27461 (.B(n_19800),
    .Y(n_19801),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_144));
 INVxp67_ASAP7_75t_SL g27462 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_56),
    .Y(n_19800));
 XNOR2xp5_ASAP7_75t_SL g27464 (.A(n_19804),
    .B(n_26112),
    .Y(n_19808));
 XNOR2xp5_ASAP7_75t_SL g27465 (.A(n_18748),
    .B(n_11852),
    .Y(n_19804));
 HB1xp67_ASAP7_75t_SL g27469 (.A(n_8150),
    .Y(n_19809));
 XNOR2x1_ASAP7_75t_SL g27471 (.B(n_19815),
    .Y(n_19816),
    .A(n_26113));
 XNOR2x1_ASAP7_75t_SL g27475 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_6),
    .Y(n_19815),
    .A(n_19814));
 INVx1_ASAP7_75t_SL g27476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_119),
    .Y(n_19814));
 MAJIxp5_ASAP7_75t_SL g27479 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_105),
    .B(n_19753),
    .C(n_19752),
    .Y(n_19820));
 NAND2xp67_ASAP7_75t_SL g27480 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_23),
    .Y(n_19821));
 XNOR2x1_ASAP7_75t_SL g27483 (.B(n_19826),
    .Y(n_19827),
    .A(n_19825));
 XNOR2xp5_ASAP7_75t_SL g27484 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_17),
    .B(n_20770),
    .Y(n_19825));
 XNOR2x1_ASAP7_75t_SL g27485 (.B(n_26196),
    .Y(n_19826),
    .A(n_5904));
 MAJIxp5_ASAP7_75t_SL g27486 (.A(n_19829),
    .B(n_19832),
    .C(n_19833),
    .Y(n_19834));
 INVx1_ASAP7_75t_SL g27489 (.A(n_10778),
    .Y(n_19830));
 INVx1_ASAP7_75t_SL g27490 (.A(n_13456),
    .Y(n_19831));
 MAJIxp5_ASAP7_75t_SL g27491 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_86),
    .Y(n_19833));
 OAI22xp5_ASAP7_75t_SL g27492 (.A1(n_13456),
    .A2(n_10778),
    .B1(n_19830),
    .B2(n_19831),
    .Y(n_19835));
 AND3x2_ASAP7_75t_SL g27496 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[3]),
    .Y(n_19838));
 INVxp33_ASAP7_75t_SL g27499 (.A(n_19838),
    .Y(n_19840));
 NAND2x1_ASAP7_75t_SL g275 (.A(n_21283),
    .B(n_19695),
    .Y(n_4286));
 AOI221xp5_ASAP7_75t_SL g27500 (.A1(n_19844),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_196),
    .B1(n_18957),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_195),
    .C(n_26216),
    .Y(n_19850));
 INVx1_ASAP7_75t_SL g27501 (.A(n_18957),
    .Y(n_19844));
 INVx1_ASAP7_75t_SL g27502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_196));
 OAI22xp33_ASAP7_75t_SL g27507 (.A1(n_18957),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_195),
    .B1(n_19844),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_196),
    .Y(n_19851));
 OAI22xp5_ASAP7_75t_SL g27511 (.A1(n_19857),
    .A2(n_19858),
    .B1(n_19859),
    .B2(n_19860),
    .Y(n_19861));
 INVx2_ASAP7_75t_SL g27512 (.A(n_19856),
    .Y(n_19857));
 XOR2x1_ASAP7_75t_SL g27513 (.A(n_18961),
    .Y(n_19856),
    .B(n_19855));
 INVxp67_ASAP7_75t_SL g27514 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_86),
    .Y(n_19855));
 XNOR2x2_ASAP7_75t_SL g27515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_30),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_114),
    .Y(n_19858));
 INVxp67_ASAP7_75t_SL g27516 (.A(n_19857),
    .Y(n_19859));
 INVx2_ASAP7_75t_SL g27517 (.A(n_19858),
    .Y(n_19860));
 OAI22xp5_ASAP7_75t_SL g27518 (.A1(n_19866),
    .A2(n_19867),
    .B1(n_19865),
    .B2(n_19868),
    .Y(n_19869));
 MAJx2_ASAP7_75t_SL g27520 (.A(n_19862),
    .B(n_19863),
    .C(n_19864),
    .Y(n_19865));
 INVx1_ASAP7_75t_SL g27521 (.A(n_9244),
    .Y(n_19862));
 INVx1_ASAP7_75t_SL g27522 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_577),
    .Y(n_19863));
 INVx1_ASAP7_75t_SL g27523 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_673),
    .Y(n_19864));
 XOR2x2_ASAP7_75t_L g27524 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_10),
    .B(n_13057),
    .Y(n_19867));
 XNOR2x1_ASAP7_75t_SL g27525 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_10),
    .Y(n_19868),
    .A(n_13057));
 INVx2_ASAP7_75t_SL g27526 (.A(n_19865),
    .Y(n_19866));
 XNOR2xp5_ASAP7_75t_SL g27529 (.A(n_19878),
    .B(n_26114),
    .Y(n_19882));
 XNOR2x1_ASAP7_75t_SL g27530 (.B(n_19877),
    .Y(n_19878),
    .A(n_19126));
 XNOR2x1_ASAP7_75t_SL g27536 (.B(n_26011),
    .Y(n_19890),
    .A(n_19886));
 OAI22x1_ASAP7_75t_SL g27537 (.A1(n_19884),
    .A2(n_10225),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_193),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_191),
    .Y(n_19886));
 INVx2_ASAP7_75t_SL g27538 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_191),
    .Y(n_19884));
 AND3x1_ASAP7_75t_SL g27545 (.A(n_19645),
    .B(n_19892),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .Y(n_19893));
 NAND2xp5_ASAP7_75t_SL g27546 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .Y(n_19892));
 AND2x2_ASAP7_75t_SL g27547 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(n_14975),
    .Y(n_19894));
 XOR2xp5_ASAP7_75t_SL g27550 (.A(n_19899),
    .B(n_19900),
    .Y(n_19901));
 MAJIxp5_ASAP7_75t_SL g27551 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_171),
    .B(n_9756),
    .C(n_23555),
    .Y(n_19898));
 XOR2xp5_ASAP7_75t_SL g27552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_148),
    .B(n_10303),
    .Y(n_19900));
 XNOR2xp5_ASAP7_75t_SL g27554 (.A(n_19905),
    .B(n_19908),
    .Y(n_19909));
 OAI21x1_ASAP7_75t_SL g27556 (.A1(n_12255),
    .A2(n_19903),
    .B(n_19904),
    .Y(n_19905));
 AND2x2_ASAP7_75t_SL g27557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_9),
    .Y(n_19903));
 OR2x2_ASAP7_75t_SL g27558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_9),
    .Y(n_19904));
 OAI22xp5_ASAP7_75t_SL g27559 (.A1(n_19907),
    .A2(n_10771),
    .B1(n_20311),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_216),
    .Y(n_19908));
 HB1xp67_ASAP7_75t_SL g27560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_215),
    .Y(n_19907));
 XNOR2xp5_ASAP7_75t_SL g27561 (.A(n_7620),
    .B(n_19911),
    .Y(n_19912));
 MAJIxp5_ASAP7_75t_SL g27562 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_203),
    .B(n_22413),
    .C(n_15003),
    .Y(n_19910));
 XNOR2xp5_ASAP7_75t_SL g27563 (.A(n_19913),
    .B(n_19914),
    .Y(n_19915));
 AOI22xp5_ASAP7_75t_SL g27564 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_17),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_89),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_90),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_74),
    .Y(n_19914));
 NOR2x1_ASAP7_75t_SL g27567 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252),
    .B(n_13196),
    .Y(n_19917));
 NAND2xp5_ASAP7_75t_SL g27568 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252),
    .B(n_13196),
    .Y(n_19918));
 NAND2xp5_ASAP7_75t_SL g27577 (.A(n_19928),
    .B(n_19929),
    .Y(n_19930));
 AOI21xp5_ASAP7_75t_SL g27578 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_445),
    .A2(n_23580),
    .B(n_4082),
    .Y(n_19928));
 AOI21xp33_ASAP7_75t_SL g27579 (.A1(n_14152),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .B(n_6039),
    .Y(n_19929));
 XNOR2xp5_ASAP7_75t_SL g27594 (.A(n_19821),
    .B(n_19820),
    .Y(n_19945));
 XNOR2x1_ASAP7_75t_SL g27596 (.B(n_19949),
    .Y(n_19950),
    .A(n_19948));
 BUFx2_ASAP7_75t_SL g27597 (.A(n_13475),
    .Y(n_19948));
 XNOR2xp5_ASAP7_75t_SL g27598 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .Y(n_19949));
 NOR2xp33_ASAP7_75t_SL g27599 (.A(n_19951),
    .B(n_13848),
    .Y(n_19952));
 XNOR2x2_ASAP7_75t_SL g276 (.A(n_18758),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_202),
    .Y(n_21036));
 XOR2x2_ASAP7_75t_SL g27600 (.A(n_10642),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_151),
    .Y(n_19951));
 NAND2xp5_ASAP7_75t_SL g27601 (.A(n_19951),
    .B(n_13848),
    .Y(n_19953));
 OAI22xp5_ASAP7_75t_SL g27602 (.A1(n_13848),
    .A2(n_19954),
    .B1(n_19951),
    .B2(n_19955),
    .Y(n_19956));
 INVx1_ASAP7_75t_SL g27603 (.A(n_19951),
    .Y(n_19954));
 INVx1_ASAP7_75t_SL g27604 (.A(n_13848),
    .Y(n_19955));
 NAND2xp5_ASAP7_75t_SL g27605 (.A(n_14445),
    .B(n_19957),
    .Y(n_19958));
 XNOR2xp5_ASAP7_75t_SL g27606 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_235),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_256),
    .Y(n_19957));
 NOR2xp67_ASAP7_75t_SL g27607 (.A(n_14445),
    .B(n_19957),
    .Y(n_19959));
 XNOR2xp5_ASAP7_75t_SL g27611 (.A(n_19963),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_149),
    .Y(n_19964));
 MAJx2_ASAP7_75t_SL g27612 (.A(n_14092),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_112),
    .C(n_10163),
    .Y(n_19963));
 MAJIxp5_ASAP7_75t_SL g27613 (.A(n_19965),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_22),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_21),
    .Y(n_19967));
 INVx1_ASAP7_75t_SL g27614 (.A(n_19963),
    .Y(n_19965));
 OAI22xp33_ASAP7_75t_SL g27616 (.A1(n_19969),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_293),
    .B1(n_20360),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_294),
    .Y(n_19970));
 INVx2_ASAP7_75t_SL g27617 (.A(n_20360),
    .Y(n_19969));
 OAI21xp5_ASAP7_75t_SL g27619 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_283),
    .A2(n_20360),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_281),
    .Y(n_19971));
 NAND2xp5_ASAP7_75t_SL g27629 (.A(n_19982),
    .B(n_4022),
    .Y(n_19983));
 INVxp67_ASAP7_75t_SRAM g27630 (.A(n_19981),
    .Y(n_19982));
 NOR2xp67_ASAP7_75t_SL g27631 (.A(n_10267),
    .B(n_11961),
    .Y(n_19981));
 HB1xp67_ASAP7_75t_SL g27633 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_191),
    .Y(n_19985));
 INVx1_ASAP7_75t_SL g27660 (.A(n_21505),
    .Y(n_20012));
 MAJIxp5_ASAP7_75t_SL g27662 (.A(n_20016),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_157),
    .Y(n_20017));
 XNOR2xp5_ASAP7_75t_SL g27663 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_4),
    .Y(n_20016));
 XNOR2xp5_ASAP7_75t_SL g27664 (.A(n_9089),
    .B(n_20016),
    .Y(n_20018));
 MAJIxp5_ASAP7_75t_SL g27668 (.A(n_20022),
    .B(n_13674),
    .C(n_2271),
    .Y(n_20023));
 MAJIxp5_ASAP7_75t_SL g27669 (.A(n_9107),
    .B(n_3766),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_205),
    .Y(n_20022));
 MAJIxp5_ASAP7_75t_SL g27671 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_224),
    .B(n_20025),
    .C(n_20029),
    .Y(n_20030));
 HB1xp67_ASAP7_75t_SL g27672 (.A(n_20096),
    .Y(n_20025));
 OAI22xp5_ASAP7_75t_SL g27673 (.A1(n_20026),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_195),
    .B1(n_20027),
    .B2(n_20028),
    .Y(n_20029));
 HB1xp67_ASAP7_75t_SL g27674 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_185),
    .Y(n_20026));
 INVx1_ASAP7_75t_SL g27675 (.A(n_20026),
    .Y(n_20027));
 INVx1_ASAP7_75t_SL g27676 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_195),
    .Y(n_20028));
 XNOR2xp5_ASAP7_75t_SL g27677 (.A(n_20028),
    .B(n_26117),
    .Y(n_20034));
 OAI21xp5_ASAP7_75t_SL g27681 (.A1(n_19969),
    .A2(n_20038),
    .B(n_20041),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_70));
 INVxp67_ASAP7_75t_SL g27682 (.A(n_20037),
    .Y(n_20038));
 NAND2xp5_ASAP7_75t_SL g27683 (.A(n_24102),
    .B(n_20035),
    .Y(n_20036));
 AOI21xp33_ASAP7_75t_SL g27684 (.A1(n_20039),
    .A2(n_20037),
    .B(n_20040),
    .Y(n_20041));
 INVxp67_ASAP7_75t_SL g27685 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_298),
    .Y(n_20039));
 NOR2xp33_ASAP7_75t_SL g27686 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_211),
    .B(n_20036),
    .Y(n_20040));
 NOR2xp67_ASAP7_75t_SL g27688 (.A(n_7075),
    .B(n_20043),
    .Y(n_20044));
 XNOR2xp5_ASAP7_75t_SL g27689 (.A(n_8380),
    .B(n_9295),
    .Y(n_20043));
 NAND2xp5_ASAP7_75t_SL g27690 (.A(n_20043),
    .B(n_7075),
    .Y(n_20046));
 XNOR2x1_ASAP7_75t_SL g27696 (.B(n_8576),
    .Y(n_20054),
    .A(n_26218));
 AOI21xp33_ASAP7_75t_SL g27709 (.A1(n_22439),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_466),
    .B(n_11320),
    .Y(n_20066));
 MAJIxp5_ASAP7_75t_SL g27712 (.A(n_10157),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_86),
    .C(n_20073),
    .Y(n_20074));
 HB1xp67_ASAP7_75t_SL g27713 (.A(n_20072),
    .Y(n_20073));
 MAJIxp5_ASAP7_75t_SL g27714 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_24),
    .B(n_4968),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_108),
    .Y(n_20072));
 OAI22xp5_ASAP7_75t_SL g27715 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_86),
    .A2(n_20072),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_85),
    .B2(n_20075),
    .Y(n_20076));
 INVx1_ASAP7_75t_SL g27716 (.A(n_20072),
    .Y(n_20075));
 NOR2xp33_ASAP7_75t_SL g27717 (.A(n_10888),
    .B(n_12576),
    .Y(n_20077));
 XNOR2xp5_ASAP7_75t_SL g27722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_157),
    .B(n_10326),
    .Y(n_20083));
 MAJIxp5_ASAP7_75t_SL g27725 (.A(n_8185),
    .B(n_20087),
    .C(n_25977),
    .Y(n_20088));
 INVxp67_ASAP7_75t_SL g27726 (.A(n_20083),
    .Y(n_20087));
 XOR2x2_ASAP7_75t_SL g27730 (.A(n_21219),
    .B(n_11067),
    .Y(n_20093));
 XNOR2xp5_ASAP7_75t_SL g27732 (.A(n_19705),
    .B(n_20094),
    .Y(n_20095));
 MAJIxp5_ASAP7_75t_SL g27733 (.A(n_22051),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_20),
    .C(n_25978),
    .Y(n_20094));
 MAJIxp5_ASAP7_75t_SL g27734 (.A(n_20094),
    .B(n_19703),
    .C(n_19706),
    .Y(n_20096));
 NOR2xp67_ASAP7_75t_SL g27735 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_253),
    .B(n_20097),
    .Y(n_20098));
 XNOR2xp5_ASAP7_75t_SL g27736 (.A(n_7876),
    .B(n_7879),
    .Y(n_20097));
 NAND2xp5_ASAP7_75t_SL g27737 (.A(n_20097),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_253),
    .Y(n_20099));
 XOR2xp5_ASAP7_75t_SL g27741 (.A(n_19044),
    .B(n_12895),
    .Y(n_20103));
 MAJIxp5_ASAP7_75t_SL g27743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_204),
    .B(n_20106),
    .C(n_20107),
    .Y(n_20108));
 HB1xp67_ASAP7_75t_SL g27744 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_150),
    .Y(n_20106));
 XOR2xp5_ASAP7_75t_SL g27745 (.A(n_20109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_319),
    .Y(n_20110));
 XNOR2x1_ASAP7_75t_SL g27746 (.B(n_14684),
    .Y(n_20109),
    .A(n_13397));
 MAJIxp5_ASAP7_75t_SL g27747 (.A(n_10483),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_319),
    .C(n_20109),
    .Y(n_20111));
 XNOR2x1_ASAP7_75t_SL g27748 (.B(n_20113),
    .Y(n_20114),
    .A(n_20112));
 OAI22xp5_ASAP7_75t_SL g27749 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_167),
    .A2(n_8130),
    .B1(n_9750),
    .B2(n_8129),
    .Y(n_20112));
 BUFx2_ASAP7_75t_SL g27750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_17),
    .Y(n_20113));
 MAJIxp5_ASAP7_75t_SL g27751 (.A(n_12644),
    .B(n_20115),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_118),
    .Y(n_20116));
 NAND2x1_ASAP7_75t_SL g27752 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .Y(n_20115));
 OAI22xp5_ASAP7_75t_SL g27753 (.A1(n_20115),
    .A2(n_12644),
    .B1(n_12643),
    .B2(n_20117),
    .Y(n_20118));
 INVx1_ASAP7_75t_SL g27754 (.A(n_20115),
    .Y(n_20117));
 XNOR2xp5_ASAP7_75t_SL g27755 (.A(n_8428),
    .B(n_20120),
    .Y(n_20121));
 XNOR2xp5_ASAP7_75t_SL g27756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_80),
    .B(n_11328),
    .Y(n_20120));
 AO21x1_ASAP7_75t_SL g27758 (.A1(n_20122),
    .A2(n_20120),
    .B(n_20123),
    .Y(n_20124));
 NAND2xp33_ASAP7_75t_SL g27759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_22),
    .Y(n_20122));
 NOR2xp33_ASAP7_75t_SL g27760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_22),
    .Y(n_20123));
 XNOR2x1_ASAP7_75t_SL g27761 (.B(n_19538),
    .Y(n_20128),
    .A(n_20127));
 AO22x2_ASAP7_75t_SL g27762 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_149),
    .A2(n_20125),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_163),
    .B2(n_20126),
    .Y(n_20127));
 INVx1_ASAP7_75t_SL g27763 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_163),
    .Y(n_20125));
 INVx1_ASAP7_75t_SL g27764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_149),
    .Y(n_20126));
 OAI21xp33_ASAP7_75t_SL g27765 (.A1(n_20127),
    .A2(n_20129),
    .B(n_20133),
    .Y(n_20134));
 INVxp67_ASAP7_75t_SL g27766 (.A(n_23139),
    .Y(n_20129));
 A2O1A1Ixp33_ASAP7_75t_SL g27767 (.A1(n_20130),
    .A2(n_20131),
    .B(n_20132),
    .C(n_11984),
    .Y(n_20133));
 INVxp67_ASAP7_75t_SL g27768 (.A(n_20125),
    .Y(n_20130));
 INVxp67_ASAP7_75t_SL g27769 (.A(n_20126),
    .Y(n_20131));
 OAI21xp5_ASAP7_75t_SL g27770 (.A1(n_20130),
    .A2(n_20131),
    .B(n_20129),
    .Y(n_20132));
 OAI22xp5_ASAP7_75t_SL g27771 (.A1(n_20135),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_30),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_158),
    .B2(n_20136),
    .Y(n_20137));
 MAJIxp5_ASAP7_75t_SL g27772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_65),
    .B(n_9327),
    .C(n_22839),
    .Y(n_20135));
 INVx1_ASAP7_75t_SL g27773 (.A(n_20135),
    .Y(n_20136));
 MAJIxp5_ASAP7_75t_SL g27774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_152),
    .B(n_20138),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_30),
    .Y(n_20139));
 INVxp67_ASAP7_75t_SL g27775 (.A(n_20135),
    .Y(n_20138));
 MAJx2_ASAP7_75t_SL g27776 (.A(n_18766),
    .B(n_20142),
    .C(n_19131),
    .Y(n_20143));
 INVxp67_ASAP7_75t_SL g27777 (.A(n_20140),
    .Y(n_20142));
 XNOR2xp5_ASAP7_75t_SL g27778 (.A(n_26012),
    .B(n_26120),
    .Y(n_20148));
 MAJx2_ASAP7_75t_SL g27783 (.A(n_20149),
    .B(n_26012),
    .C(n_20151),
    .Y(n_20152));
 INVx1_ASAP7_75t_SL g27784 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_134),
    .Y(n_20149));
 OAI21xp5_ASAP7_75t_SL g27788 (.A1(n_20156),
    .A2(n_20157),
    .B(n_5870),
    .Y(n_20158));
 INVx1_ASAP7_75t_SL g27789 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_445),
    .Y(n_20157));
 OAI21xp33_ASAP7_75t_SL g27790 (.A1(n_16256),
    .A2(n_20157),
    .B(n_5867),
    .Y(n_20160));
 INVxp67_ASAP7_75t_SL g27792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_298),
    .Y(n_20161));
 NOR2xp33_ASAP7_75t_SL g27793 (.A(n_20161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_317),
    .Y(n_20163));
 MAJIxp5_ASAP7_75t_SL g27823 (.A(n_20307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_172),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_33),
    .Y(n_20195));
 NOR2xp33_ASAP7_75t_SL g27825 (.A(n_22951),
    .B(n_22952),
    .Y(n_20198));
 NAND2xp33_ASAP7_75t_SL g27826 (.A(n_22952),
    .B(n_22951),
    .Y(n_20199));
 XOR2xp5_ASAP7_75t_SL g27827 (.A(n_20307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_172),
    .Y(n_20200));
 NAND2xp5_ASAP7_75t_SL g27838 (.A(n_2820),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .Y(n_20210));
 NAND2x1_ASAP7_75t_SL g27840 (.A(n_20210),
    .B(n_19607),
    .Y(n_20214));
 MAJIxp5_ASAP7_75t_SL g27841 (.A(n_20219),
    .B(n_20220),
    .C(n_14788),
    .Y(n_20221));
 XOR2x2_ASAP7_75t_SL g27842 (.A(n_20218),
    .B(n_22632),
    .Y(n_20219));
 OAI22xp5_ASAP7_75t_SL g27843 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_106),
    .A2(n_13794),
    .B1(n_20216),
    .B2(n_20217),
    .Y(n_20218));
 INVx1_ASAP7_75t_SL g27844 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_106),
    .Y(n_20216));
 HB1xp67_ASAP7_75t_SL g27845 (.A(n_3235),
    .Y(n_20220));
 XNOR2x1_ASAP7_75t_SL g27846 (.B(n_20219),
    .Y(n_20222),
    .A(n_14791));
 XNOR2xp5_ASAP7_75t_SL g27854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_177),
    .B(n_20232),
    .Y(n_20233));
 MAJIxp5_ASAP7_75t_SL g27856 (.A(n_23470),
    .B(n_5529),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_87),
    .Y(n_20231));
 MAJIxp5_ASAP7_75t_SL g27858 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_149),
    .B(n_20231),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_158),
    .Y(n_20234));
 XOR2xp5_ASAP7_75t_SL g27859 (.A(n_18835),
    .B(n_23470),
    .Y(n_20235));
 XOR2xp5_ASAP7_75t_SL g27860 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_243),
    .B(n_20237),
    .Y(n_20238));
 OAI21xp5_ASAP7_75t_SL g27861 (.A1(n_7507),
    .A2(n_20236),
    .B(n_7508),
    .Y(n_20237));
 OA21x2_ASAP7_75t_SL g27862 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_274),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_276),
    .Y(n_20236));
 OAI21x1_ASAP7_75t_SL g27863 (.A1(n_7515),
    .A2(n_20236),
    .B(n_7517),
    .Y(n_20239));
 OAI21xp5_ASAP7_75t_SL g27893 (.A1(n_9986),
    .A2(n_20275),
    .B(n_9987),
    .Y(n_20276));
 AOI21xp5_ASAP7_75t_SL g27894 (.A1(n_9494),
    .A2(n_22786),
    .B(n_20274),
    .Y(n_20275));
 NOR2xp67_ASAP7_75t_SL g27895 (.A(n_22785),
    .B(n_22780),
    .Y(n_20274));
 INVxp67_ASAP7_75t_SL g27897 (.A(n_20275),
    .Y(n_20277));
 NAND2xp5_ASAP7_75t_SL g27898 (.A(n_20279),
    .B(n_4024),
    .Y(n_20280));
 INVxp67_ASAP7_75t_SRAM g27899 (.A(n_20274),
    .Y(n_20279));
 INVxp67_ASAP7_75t_SL g279 (.A(n_21882),
    .Y(n_21883));
 HB1xp67_ASAP7_75t_SL g27900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_86),
    .Y(n_20281));
 MAJIxp5_ASAP7_75t_SL g27901 (.A(n_9762),
    .B(n_9763),
    .C(n_20282),
    .Y(n_20283));
 NAND2xp5_ASAP7_75t_SL g27902 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .Y(n_20282));
 INVx1_ASAP7_75t_SL g27903 (.A(n_20283),
    .Y(n_20285));
 XNOR2xp5_ASAP7_75t_SL g27904 (.A(n_20287),
    .B(n_13441),
    .Y(n_20288));
 INVxp67_ASAP7_75t_SL g27905 (.A(n_20282),
    .Y(n_20287));
 OAI21xp33_ASAP7_75t_SL g27906 (.A1(n_22440),
    .A2(n_11317),
    .B(n_20290),
    .Y(n_20291));
 AOI21xp5_ASAP7_75t_SL g27907 (.A1(n_11318),
    .A2(n_22440),
    .B(n_26015),
    .Y(n_20290));
 MAJIxp5_ASAP7_75t_SL g27909 (.A(n_20292),
    .B(n_20293),
    .C(n_20295),
    .Y(n_20296));
 INVx1_ASAP7_75t_SL g27910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_5),
    .Y(n_20292));
 INVx1_ASAP7_75t_SL g27911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_127),
    .Y(n_20293));
 MAJx2_ASAP7_75t_SL g27912 (.A(n_13712),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_20),
    .C(n_20294),
    .Y(n_20295));
 NAND2xp5_ASAP7_75t_SL g27913 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .Y(n_20294));
 XOR2xp5_ASAP7_75t_SL g27914 (.A(n_10387),
    .B(n_20295),
    .Y(n_20297));
 OAI22xp5_ASAP7_75t_SL g27917 (.A1(n_20302),
    .A2(n_11943),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_158),
    .B2(n_20303),
    .Y(n_20304));
 MAJIxp5_ASAP7_75t_SL g27918 (.A(n_15142),
    .B(n_15144),
    .C(n_20301),
    .Y(n_20302));
 INVx1_ASAP7_75t_SL g27919 (.A(n_20302),
    .Y(n_20303));
 MAJIxp5_ASAP7_75t_SL g27920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_152),
    .B(n_11943),
    .C(n_20305),
    .Y(n_20306));
 INVxp67_ASAP7_75t_SL g27921 (.A(n_20302),
    .Y(n_20305));
 XNOR2xp5_ASAP7_75t_SL g27922 (.A(n_20301),
    .B(n_15145),
    .Y(n_20307));
 XOR2x2_ASAP7_75t_SL g27923 (.A(n_20310),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_192),
    .Y(n_20311));
 XOR2xp5_ASAP7_75t_SL g27924 (.A(n_26016),
    .B(n_20309),
    .Y(n_20310));
 XNOR2xp5_ASAP7_75t_SL g27926 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_108),
    .B(n_20590),
    .Y(n_20309));
 MAJIxp5_ASAP7_75t_SL g27927 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_192),
    .B(n_20312),
    .C(n_20313),
    .Y(n_20314));
 INVxp67_ASAP7_75t_SL g27928 (.A(n_26016),
    .Y(n_20312));
 HB1xp67_ASAP7_75t_SL g27929 (.A(n_20309),
    .Y(n_20313));
 HB1xp67_ASAP7_75t_SL g27938 (.A(n_8228),
    .Y(n_20329));
 AO21x1_ASAP7_75t_SL g27939 (.A1(n_20333),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_212),
    .B(n_20334),
    .Y(n_20335));
 OR2x2_ASAP7_75t_SL g27940 (.A(n_20332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_203),
    .Y(n_20333));
 XNOR2x1_ASAP7_75t_SL g27941 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_133),
    .Y(n_20332),
    .A(n_20331));
 XNOR2xp5_ASAP7_75t_SL g27942 (.A(n_20330),
    .B(n_6243),
    .Y(n_20331));
 INVx1_ASAP7_75t_SL g27943 (.A(n_8228),
    .Y(n_20330));
 AND2x2_ASAP7_75t_SL g27944 (.A(n_20332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_203),
    .Y(n_20334));
 XNOR2x1_ASAP7_75t_SL g27945 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_203),
    .Y(n_20336),
    .A(n_20332));
 INVx1_ASAP7_75t_SL g27952 (.A(n_20344),
    .Y(n_20345));
 NAND2x1p5_ASAP7_75t_SL g27953 (.A(n_7052),
    .B(n_20343),
    .Y(n_20344));
 OA21x2_ASAP7_75t_SL g27954 (.A1(n_11781),
    .A2(n_7053),
    .B(n_23021),
    .Y(n_20343));
 AOI21xp5_ASAP7_75t_SL g27955 (.A1(n_20344),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_304),
    .B(n_5471),
    .Y(n_20346));
 AND2x2_ASAP7_75t_SL g27956 (.A(n_20344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_304),
    .Y(n_20347));
 XOR2xp5_ASAP7_75t_SL g27962 (.A(n_20354),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .Y(n_20355));
 OAI21xp5_ASAP7_75t_SL g27963 (.A1(n_20353),
    .A2(n_11998),
    .B(n_11026),
    .Y(n_20354));
 NOR2xp33_ASAP7_75t_SL g27964 (.A(n_11022),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_647),
    .Y(n_20353));
 MAJx2_ASAP7_75t_SL g27965 (.A(n_22716),
    .B(n_16247),
    .C(n_20356),
    .Y(n_20357));
 HB1xp67_ASAP7_75t_SL g27966 (.A(n_20354),
    .Y(n_20356));
 AOI21x1_ASAP7_75t_SL g27967 (.A1(n_14800),
    .A2(n_20359),
    .B(n_11768),
    .Y(n_20360));
 NOR2xp67_ASAP7_75t_SL g27968 (.A(n_20358),
    .B(n_19732),
    .Y(n_20359));
 NAND2xp5_ASAP7_75t_SL g27969 (.A(n_19729),
    .B(n_19730),
    .Y(n_20358));
 OAI21xp5_ASAP7_75t_SL g27970 (.A1(n_20363),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307),
    .B(n_20371),
    .Y(n_20372));
 INVxp67_ASAP7_75t_SL g27971 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_226),
    .Y(n_20361));
 INVxp67_ASAP7_75t_SL g27972 (.A(n_2159),
    .Y(n_20362));
 AOI21xp33_ASAP7_75t_SRAM g27974 (.A1(n_26123),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307),
    .B(n_20370),
    .Y(n_20371));
 NOR2xp33_ASAP7_75t_SL g27976 (.A(n_20362),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_226),
    .Y(n_20365));
 OAI21xp5_ASAP7_75t_SL g27977 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_288),
    .A2(n_20363),
    .B(n_20369),
    .Y(n_20370));
 NAND2xp5_ASAP7_75t_SL g27978 (.A(n_20365),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_291),
    .Y(n_20369));
 XOR2xp5_ASAP7_75t_SL g27979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_80),
    .B(n_20375),
    .Y(n_20376));
 OAI22xp5_ASAP7_75t_SL g27980 (.A1(n_20373),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_94),
    .B1(n_20374),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_93),
    .Y(n_20375));
 NAND2xp5_ASAP7_75t_SL g27981 (.A(n_4831),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .Y(n_20373));
 INVx1_ASAP7_75t_SL g27982 (.A(n_20373),
    .Y(n_20374));
 MAJIxp5_ASAP7_75t_SL g27983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_80),
    .C(n_20373),
    .Y(n_20377));
 XNOR2x1_ASAP7_75t_SL g27986 (.B(n_20379),
    .Y(n_20380),
    .A(n_26044));
 XOR2x2_ASAP7_75t_SL g27987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_127),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_75),
    .Y(n_20379));
 MAJIxp5_ASAP7_75t_SL g27989 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_213),
    .B(n_20383),
    .C(n_20384),
    .Y(n_20385));
 HB1xp67_ASAP7_75t_SL g27990 (.A(n_5781),
    .Y(n_20383));
 HB1xp67_ASAP7_75t_SL g27991 (.A(n_20380),
    .Y(n_20384));
 AOI21xp5_ASAP7_75t_SL g27998 (.A1(n_19254),
    .A2(n_11338),
    .B(n_5630),
    .Y(n_20390));
 NOR2x1_ASAP7_75t_SL g28 (.A(n_9058),
    .B(n_9059),
    .Y(n_9060));
 NOR2xp33_ASAP7_75t_SL g280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_362),
    .B(n_10264),
    .Y(n_21892));
 INVxp67_ASAP7_75t_SL g28000 (.A(n_20390),
    .Y(n_20393));
 INVxp67_ASAP7_75t_SL g281 (.A(n_8563),
    .Y(n_8572));
 NAND2xp5_ASAP7_75t_L g28136 (.A(n_2182),
    .B(n_21595),
    .Y(n_20588));
 XNOR2x1_ASAP7_75t_SL g28138 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_101),
    .Y(n_20590),
    .A(n_9534));
 NOR2xp33_ASAP7_75t_SL g28144 (.A(n_20645),
    .B(n_11869),
    .Y(n_20646));
 AOI221xp5_ASAP7_75t_SL g28145 (.A1(n_20641),
    .A2(n_20765),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_208),
    .B2(n_20642),
    .C(n_20644),
    .Y(n_20645));
 MAJIxp5_ASAP7_75t_SL g28146 (.A(n_3973),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_190),
    .C(n_20643),
    .Y(n_20644));
 HB1xp67_ASAP7_75t_SL g28147 (.A(n_20134),
    .Y(n_20643));
 OAI21x1_ASAP7_75t_SL g28149 (.A1(n_6008),
    .A2(n_20390),
    .B(n_11213),
    .Y(n_20650));
 NAND2xp5_ASAP7_75t_SL g28150 (.A(n_20644),
    .B(n_20652),
    .Y(n_20653));
 XNOR2xp5_ASAP7_75t_SL g28151 (.A(n_20642),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_208),
    .Y(n_20652));
 NOR2xp67_ASAP7_75t_SL g28154 (.A(n_20644),
    .B(n_20652),
    .Y(n_20659));
 NAND2xp5_ASAP7_75t_SL g28155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_193),
    .B(n_20638),
    .Y(n_20660));
 XOR2x2_ASAP7_75t_SL g28165 (.A(n_20671),
    .B(n_26004),
    .Y(n_20673));
 OAI21x1_ASAP7_75t_SL g28166 (.A1(n_13667),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .B(n_20670),
    .Y(n_20671));
 OR2x2_ASAP7_75t_SL g28167 (.A(n_20833),
    .B(n_6673),
    .Y(n_20670));
 NAND2x1_ASAP7_75t_SL g28171 (.A(n_3317),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .Y(n_20675));
 NOR2x1_ASAP7_75t_SL g28174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252),
    .B(n_13196),
    .Y(n_20680));
 XNOR2x1_ASAP7_75t_SL g28175 (.B(n_18956),
    .Y(n_13196),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_236));
 OR2x2_ASAP7_75t_SL g28177 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_269),
    .B(n_19533),
    .Y(n_20681));
 AND2x2_ASAP7_75t_SL g28179 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_269),
    .B(n_19534),
    .Y(n_20682));
 AO21x1_ASAP7_75t_SL g28180 (.A1(n_20682),
    .A2(n_19533),
    .B(n_20683),
    .Y(n_20684));
 NOR2xp33_ASAP7_75t_SL g28181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_269),
    .B(n_19534),
    .Y(n_20683));
 MAJIxp5_ASAP7_75t_SL g28182 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_140),
    .C(n_20688),
    .Y(n_20689));
 XNOR2x1_ASAP7_75t_SL g28183 (.B(n_17710),
    .Y(n_20688),
    .A(n_20687));
 HB1xp67_ASAP7_75t_SL g28184 (.A(n_17707),
    .Y(n_20687));
 AOI22xp5_ASAP7_75t_SL g28195 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_43),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_85),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_84),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_44),
    .Y(n_20700));
 NAND2xp5_ASAP7_75t_SL g282 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .B(n_3112),
    .Y(n_8563));
 XNOR2x1_ASAP7_75t_SL g28209 (.B(n_20718),
    .Y(n_20719),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_178));
 XNOR2xp5_ASAP7_75t_SL g28210 (.A(n_20716),
    .B(n_20717),
    .Y(n_20718));
 OAI21x1_ASAP7_75t_SL g28211 (.A1(n_8527),
    .A2(n_8522),
    .B(n_8528),
    .Y(n_20716));
 XNOR2xp5_ASAP7_75t_SL g28212 (.A(n_7938),
    .B(n_21795),
    .Y(n_20717));
 MAJIxp5_ASAP7_75t_SL g28215 (.A(n_18757),
    .B(n_20727),
    .C(n_9584),
    .Y(n_20728));
 HB1xp67_ASAP7_75t_SL g28216 (.A(n_20726),
    .Y(n_20727));
 XOR2x2_ASAP7_75t_SL g28217 (.A(n_20723),
    .B(n_20725),
    .Y(n_20726));
 XOR2xp5_ASAP7_75t_SL g28218 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_67),
    .Y(n_20723));
 INVxp67_ASAP7_75t_SL g28219 (.A(n_20724),
    .Y(n_20725));
 NAND2xp5_ASAP7_75t_SL g28220 (.A(n_14183),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .Y(n_20724));
 XNOR2x1_ASAP7_75t_SL g28221 (.B(n_9584),
    .Y(n_20729),
    .A(n_20726));
 MAJIxp5_ASAP7_75t_SL g28222 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_67),
    .C(n_20724),
    .Y(n_20730));
 NOR2xp67_ASAP7_75t_SL g28225 (.A(n_12088),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_400),
    .Y(n_20731));
 INVx1_ASAP7_75t_SL g28228 (.A(n_21322),
    .Y(n_10309));
 INVxp67_ASAP7_75t_SL g28229 (.A(n_22458),
    .Y(n_20737));
 OAI22xp33_ASAP7_75t_SL g28230 (.A1(n_22323),
    .A2(n_20740),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_488),
    .B2(n_20739),
    .Y(n_20741));
 INVxp67_ASAP7_75t_SL g28231 (.A(n_20739),
    .Y(n_20740));
 NOR2xp33_ASAP7_75t_SL g28232 (.A(n_20731),
    .B(n_23753),
    .Y(n_20739));
 INVxp33_ASAP7_75t_SRAM g28233 (.A(n_20731),
    .Y(n_20742));
 NOR2x1p5_ASAP7_75t_SL g28243 (.A(n_20752),
    .B(n_21098),
    .Y(n_20758));
 NAND2xp5_ASAP7_75t_SL g28249 (.A(n_21098),
    .B(n_22101),
    .Y(n_20759));
 MAJIxp5_ASAP7_75t_SL g28251 (.A(n_20764),
    .B(n_20281),
    .C(n_20283),
    .Y(n_20765));
 MAJIxp5_ASAP7_75t_SL g28258 (.A(n_20769),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_55),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_73),
    .Y(n_20770));
 NAND2xp5_ASAP7_75t_SL g28259 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .Y(n_20769));
 XNOR2xp5_ASAP7_75t_SL g28260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_55),
    .B(n_20769),
    .Y(n_20771));
 INVxp67_ASAP7_75t_SL g28266 (.A(n_2169),
    .Y(n_20776));
 NOR2xp33_ASAP7_75t_SL g28267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_193),
    .Y(n_20777));
 NOR2xp67_ASAP7_75t_SL g28268 (.A(n_20782),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_20783));
 INVx2_ASAP7_75t_SL g28269 (.A(n_23830),
    .Y(n_20782));
 NAND2xp5_ASAP7_75t_SL g28270 (.A(n_20782),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_20784));
 OR2x2_ASAP7_75t_SL g28271 (.A(n_20773),
    .B(n_20777),
    .Y(n_20785));
 XNOR2xp5_ASAP7_75t_SL g28273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_567),
    .B(n_20788),
    .Y(n_20789));
 XOR2xp5_ASAP7_75t_SL g28274 (.A(n_20787),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_599),
    .Y(n_20788));
 NAND2xp5_ASAP7_75t_SL g28275 (.A(n_20825),
    .B(n_6878),
    .Y(n_20787));
 MAJIxp5_ASAP7_75t_SL g28277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .B(n_20789),
    .C(n_20793),
    .Y(n_20794));
 HB1xp67_ASAP7_75t_SL g28278 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .Y(n_20793));
 MAJIxp5_ASAP7_75t_SL g28279 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_567),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_599),
    .C(n_20795),
    .Y(n_20796));
 INVxp67_ASAP7_75t_SL g28280 (.A(n_20787),
    .Y(n_20795));
 XNOR2xp5_ASAP7_75t_SL g28291 (.A(n_11835),
    .B(n_9261),
    .Y(n_20809));
 MAJx2_ASAP7_75t_SL g28292 (.A(n_20810),
    .B(n_20812),
    .C(n_20813),
    .Y(n_20814));
 MAJx2_ASAP7_75t_SL g28293 (.A(n_7874),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_140),
    .Y(n_20810));
 XOR2x2_ASAP7_75t_SL g28294 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_4),
    .B(n_20811),
    .Y(n_20812));
 INVxp67_ASAP7_75t_SL g28295 (.A(n_22628),
    .Y(n_20811));
 XOR2xp5_ASAP7_75t_SL g28296 (.A(n_19685),
    .B(n_6949),
    .Y(n_20813));
 HB1xp67_ASAP7_75t_SL g283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_121),
    .Y(n_23085));
 XNOR2x1_ASAP7_75t_SL g28300 (.B(n_20832),
    .Y(n_20833),
    .A(n_20824));
 XNOR2x1_ASAP7_75t_SL g28301 (.B(n_10595),
    .Y(n_20824),
    .A(n_20823));
 INVx1_ASAP7_75t_SL g28302 (.A(n_19264),
    .Y(n_20823));
 HB1xp67_ASAP7_75t_SL g28303 (.A(n_20831),
    .Y(n_20832));
 OAI21x1_ASAP7_75t_L g28304 (.A1(n_20828),
    .A2(n_4865),
    .B(n_20830),
    .Y(n_20831));
 OR2x2_ASAP7_75t_SL g28305 (.A(n_26226),
    .B(n_20979),
    .Y(n_20828));
 AND3x1_ASAP7_75t_SL g28307 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[2]),
    .Y(n_20825));
 INVx1_ASAP7_75t_SL g28309 (.A(n_20829),
    .Y(n_20830));
 OAI22xp5_ASAP7_75t_SL g28310 (.A1(n_20977),
    .A2(n_20828),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_189),
    .B2(n_26226),
    .Y(n_20829));
 XOR2xp5_ASAP7_75t_SL g28317 (.A(n_20841),
    .B(n_20844),
    .Y(n_20845));
 MAJx2_ASAP7_75t_SL g28318 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_172),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_186),
    .Y(n_20841));
 XNOR2xp5_ASAP7_75t_SL g28319 (.A(n_20842),
    .B(n_20843),
    .Y(n_20844));
 XOR2xp5_ASAP7_75t_SL g28320 (.A(n_20700),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_51),
    .Y(n_20842));
 OAI22xp5_ASAP7_75t_SL g28321 (.A1(n_21988),
    .A2(n_19387),
    .B1(n_19386),
    .B2(n_19385),
    .Y(n_20843));
 AOI22xp5_ASAP7_75t_SL g28322 (.A1(n_20849),
    .A2(n_20850),
    .B1(n_20851),
    .B2(n_20852),
    .Y(n_20853));
 NAND2xp33_ASAP7_75t_SL g28323 (.A(n_20847),
    .B(n_21064),
    .Y(n_20849));
 INVxp67_ASAP7_75t_SL g28324 (.A(n_21059),
    .Y(n_20847));
 XNOR2xp5_ASAP7_75t_SL g28327 (.A(n_13525),
    .B(n_19015),
    .Y(n_20850));
 INVxp67_ASAP7_75t_SL g28328 (.A(n_21064),
    .Y(n_20851));
 INVxp67_ASAP7_75t_SL g28329 (.A(n_20847),
    .Y(n_20852));
 XOR2xp5_ASAP7_75t_SL g28331 (.A(n_20855),
    .B(n_20856),
    .Y(n_20857));
 NAND2xp5_ASAP7_75t_SL g28332 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .Y(n_20855));
 NAND2x1_ASAP7_75t_SL g28333 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .B(n_11770),
    .Y(n_20856));
 INVxp33_ASAP7_75t_SL g28334 (.A(n_20855),
    .Y(n_20047));
 NAND2x1p5_ASAP7_75t_SL g28335 (.A(n_20863),
    .B(n_20867),
    .Y(n_20868));
 OAI21xp5_ASAP7_75t_SL g28336 (.A1(n_20233),
    .A2(n_20861),
    .B(n_20862),
    .Y(n_20863));
 NOR2xp67_ASAP7_75t_SL g28337 (.A(n_20859),
    .B(n_20860),
    .Y(n_20861));
 INVx1_ASAP7_75t_SL g28338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_194),
    .Y(n_20859));
 INVx2_ASAP7_75t_SL g28339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_9),
    .Y(n_20860));
 NAND2xp5_ASAP7_75t_SL g28340 (.A(n_20859),
    .B(n_20860),
    .Y(n_20862));
 XNOR2x2_ASAP7_75t_SL g28341 (.A(n_20865),
    .B(n_20866),
    .Y(n_20867));
 XOR2x1_ASAP7_75t_SL g28342 (.A(n_19222),
    .Y(n_20865),
    .B(n_20864));
 HB1xp67_ASAP7_75t_SL g28343 (.A(n_19834),
    .Y(n_20864));
 XNOR2xp5_ASAP7_75t_SL g28344 (.A(n_14143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_191),
    .Y(n_20866));
 XNOR2xp5_ASAP7_75t_SL g28345 (.A(n_20871),
    .B(n_20872),
    .Y(n_20873));
 XOR2xp5_ASAP7_75t_SL g28346 (.A(n_20869),
    .B(n_20870),
    .Y(n_20871));
 MAJIxp5_ASAP7_75t_SL g28347 (.A(n_25298),
    .B(n_25294),
    .C(n_23941),
    .Y(n_20869));
 XNOR2xp5_ASAP7_75t_SL g28348 (.A(n_6456),
    .B(n_23987),
    .Y(n_20870));
 XOR2x2_ASAP7_75t_SL g28349 (.A(n_21947),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_277),
    .Y(n_20872));
 XNOR2xp5_ASAP7_75t_SL g28350 (.A(n_20882),
    .B(n_20883),
    .Y(n_20884));
 NAND2x1_ASAP7_75t_SL g28351 (.A(n_20878),
    .B(n_20881),
    .Y(n_20882));
 OAI21xp5_ASAP7_75t_SL g28352 (.A1(n_20874),
    .A2(n_20875),
    .B(n_20877),
    .Y(n_20878));
 INVxp67_ASAP7_75t_SL g28353 (.A(n_4826),
    .Y(n_20874));
 INVxp67_ASAP7_75t_SL g28354 (.A(n_21861),
    .Y(n_20875));
 INVx1_ASAP7_75t_SL g28355 (.A(n_20876),
    .Y(n_20877));
 NAND2xp5_ASAP7_75t_SL g28356 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .Y(n_20876));
 NAND2xp5_ASAP7_75t_SL g28357 (.A(n_20876),
    .B(n_26021),
    .Y(n_20881));
 MAJIxp5_ASAP7_75t_SL g28359 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_41),
    .B(n_23400),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_44),
    .Y(n_20883));
 NAND2xp5_ASAP7_75t_SL g28362 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(n_20887));
 NAND2xp5_ASAP7_75t_SL g28363 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .Y(n_20888));
 INVx1_ASAP7_75t_SL g28366 (.A(n_20888),
    .Y(n_20893));
 XOR2xp5_ASAP7_75t_SL g28367 (.A(n_20897),
    .B(n_20899),
    .Y(n_20900));
 XOR2xp5_ASAP7_75t_SL g28368 (.A(n_20895),
    .B(n_20896),
    .Y(n_20897));
 XNOR2xp5_ASAP7_75t_SL g28369 (.A(n_20894),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_143),
    .Y(n_20895));
 INVx1_ASAP7_75t_SL g28370 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_99),
    .Y(n_20894));
 MAJx2_ASAP7_75t_SL g28371 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_44),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_51),
    .Y(n_20896));
 XNOR2xp5_ASAP7_75t_SL g28372 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_145),
    .Y(n_20898));
 MAJIxp5_ASAP7_75t_SL g28374 (.A(n_20905),
    .B(n_20909),
    .C(n_20912),
    .Y(n_20913));
 NOR2xp33_ASAP7_75t_SL g28375 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_144),
    .Y(n_20902));
 NOR2xp67_ASAP7_75t_SL g28376 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_160),
    .Y(n_20903));
 NAND2xp5_ASAP7_75t_SL g28377 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_160),
    .Y(n_20904));
 MAJIxp5_ASAP7_75t_SRAM g28378 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_45),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_29),
    .Y(n_20909));
 AO22x1_ASAP7_75t_SL g28381 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_162),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_158),
    .B1(n_20911),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_157),
    .Y(n_20912));
 INVxp67_ASAP7_75t_SL g28383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_162),
    .Y(n_20911));
 HB1xp67_ASAP7_75t_SL g28384 (.A(n_20913),
    .Y(n_20914));
 NOR2x1_ASAP7_75t_SL g28386 (.A(n_20916),
    .B(n_20921),
    .Y(n_20922));
 NOR3xp33_ASAP7_75t_SL g28387 (.A(n_2718),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_119),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_40),
    .Y(n_20916));
 XNOR2xp5_ASAP7_75t_SL g28388 (.A(n_20917),
    .B(n_26127),
    .Y(n_20921));
 AOI22xp5_ASAP7_75t_SL g28389 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_116),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_76),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_115),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_75),
    .Y(n_20917));
 XNOR2xp5_ASAP7_75t_SL g28393 (.A(n_20923),
    .B(n_20924),
    .Y(n_20925));
 NAND2xp5_ASAP7_75t_SL g28394 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(n_20923));
 NAND2xp5_ASAP7_75t_SL g28395 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .Y(n_20924));
 XNOR2xp5_ASAP7_75t_SL g28396 (.A(n_20926),
    .B(n_20927),
    .Y(n_20928));
 NAND2xp5_ASAP7_75t_SL g28397 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .Y(n_20926));
 NAND2xp5_ASAP7_75t_SL g28398 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .Y(n_20927));
 AOI21xp5_ASAP7_75t_SL g284 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_239),
    .A2(n_14038),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_240),
    .Y(n_12051));
 XNOR2xp5_ASAP7_75t_SL g28401 (.A(n_20933),
    .B(n_20934),
    .Y(n_20935));
 HB1xp67_ASAP7_75t_SL g28402 (.A(n_9154),
    .Y(n_20932));
 MAJIxp5_ASAP7_75t_SL g28406 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_675),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_547),
    .C(n_13544),
    .Y(n_20943));
 NAND2xp5_ASAP7_75t_SL g28407 (.A(n_20946),
    .B(n_20939),
    .Y(n_19792));
 OAI21xp5_ASAP7_75t_SL g28408 (.A1(n_10848),
    .A2(n_10847),
    .B(n_18774),
    .Y(n_19787));
 OAI21xp5_ASAP7_75t_SL g28409 (.A1(n_20954),
    .A2(n_20957),
    .B(n_20964),
    .Y(n_20965));
 NOR2xp33_ASAP7_75t_SL g28410 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_101),
    .Y(n_20949));
 NOR2xp33_ASAP7_75t_SL g28411 (.A(n_20949),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_138),
    .Y(n_20953));
 AND2x2_ASAP7_75t_SL g28413 (.A(n_25979),
    .B(n_20956),
    .Y(n_20957));
 INVxp67_ASAP7_75t_SL g28415 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_123),
    .Y(n_20956));
 AO21x1_ASAP7_75t_SL g28416 (.A1(n_20959),
    .A2(n_20961),
    .B(n_20963),
    .Y(n_20964));
 NAND2xp5_ASAP7_75t_SL g28417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_131),
    .Y(n_20959));
 NAND2xp5_ASAP7_75t_SL g28419 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_138),
    .B(n_20951),
    .Y(n_20961));
 INVx1_ASAP7_75t_SL g28421 (.A(n_20949),
    .Y(n_20963));
 AO21x1_ASAP7_75t_SL g28423 (.A1(n_20959),
    .A2(n_20961),
    .B(n_20963),
    .Y(n_20966));
 XNOR2xp5_ASAP7_75t_SL g28424 (.A(n_20969),
    .B(n_20973),
    .Y(n_20974));
 HB1xp67_ASAP7_75t_SL g28425 (.A(n_20968),
    .Y(n_20969));
 MAJIxp5_ASAP7_75t_SL g28426 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_184),
    .B(n_20967),
    .C(n_18758),
    .Y(n_20968));
 XOR2xp5_ASAP7_75t_SL g28428 (.A(n_20971),
    .B(n_20972),
    .Y(n_20973));
 INVxp67_ASAP7_75t_SL g28429 (.A(n_26227),
    .Y(n_20971));
 XNOR2x2_ASAP7_75t_SL g28431 (.A(n_6605),
    .B(n_21867),
    .Y(n_20972));
 XOR2xp5_ASAP7_75t_SL g28433 (.A(n_20981),
    .B(n_20982),
    .Y(n_20983));
 AOI21xp5_ASAP7_75t_SL g28434 (.A1(n_20976),
    .A2(n_20977),
    .B(n_20979),
    .Y(n_20981));
 OAI21x1_ASAP7_75t_SL g28435 (.A1(n_4861),
    .A2(n_7015),
    .B(n_7021),
    .Y(n_20976));
 OAI21xp5_ASAP7_75t_SL g28438 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_232),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_236),
    .Y(n_20979));
 OAI21xp33_ASAP7_75t_SL g28439 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_65),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_189),
    .Y(n_20982));
 AND2x2_ASAP7_75t_SL g28440 (.A(n_13030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_720),
    .Y(n_20984));
 XNOR2xp5_ASAP7_75t_SL g28441 (.A(n_20985),
    .B(n_20986),
    .Y(n_20987));
 NAND2x1_ASAP7_75t_SL g28442 (.A(n_2181),
    .B(n_23132),
    .Y(n_20985));
 NAND2x1_ASAP7_75t_SL g28443 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_784),
    .Y(n_20986));
 INVx1_ASAP7_75t_SL g28444 (.A(n_20986),
    .Y(n_20989));
 INVx1_ASAP7_75t_SL g28445 (.A(n_20985),
    .Y(n_20990));
 XOR2xp5_ASAP7_75t_SL g28448 (.A(n_22524),
    .B(n_20993),
    .Y(n_20994));
 MAJIxp5_ASAP7_75t_SL g28450 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_95),
    .B(n_9926),
    .C(n_5423),
    .Y(n_20993));
 HB1xp67_ASAP7_75t_SL g28452 (.A(n_20996),
    .Y(n_20997));
 MAJIxp5_ASAP7_75t_SL g28453 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_80),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_89),
    .Y(n_20996));
 XOR2xp5_ASAP7_75t_SL g28454 (.A(n_20998),
    .B(n_20999),
    .Y(n_21000));
 XNOR2xp5_ASAP7_75t_SL g28455 (.A(n_6905),
    .B(n_6910),
    .Y(n_20998));
 XNOR2xp5_ASAP7_75t_SL g28456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_128),
    .Y(n_20999));
 XNOR2xp5_ASAP7_75t_SL g28457 (.A(n_21002),
    .B(n_26129),
    .Y(n_21010));
 AO21x1_ASAP7_75t_SL g28458 (.A1(n_8377),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_148),
    .B(n_8378),
    .Y(n_21002));
 XOR2x2_ASAP7_75t_SL g28461 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_126),
    .B(n_25990),
    .Y(n_21004));
 MAJx2_ASAP7_75t_SL g28463 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_19),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_18),
    .Y(n_21007));
 HB1xp67_ASAP7_75t_SL g28468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_128),
    .Y(n_21013));
 AOI221x1_ASAP7_75t_SL g28469 (.A1(n_21016),
    .A2(n_26130),
    .B1(n_21015),
    .B2(n_21020),
    .C(n_26228),
    .Y(n_21025));
 INVx2_ASAP7_75t_SL g28470 (.A(n_21015),
    .Y(n_21016));
 XNOR2x2_ASAP7_75t_SL g28471 (.A(n_21014),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_125),
    .Y(n_21015));
 INVxp67_ASAP7_75t_SL g28472 (.A(n_22633),
    .Y(n_21014));
 INVx1_ASAP7_75t_SL g28474 (.A(n_26130),
    .Y(n_21020));
 OR2x2_ASAP7_75t_SL g28480 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_71),
    .B(n_22634),
    .Y(n_21023));
 OAI22xp5_ASAP7_75t_SL g28481 (.A1(n_21026),
    .A2(n_21015),
    .B1(n_26130),
    .B2(n_21016),
    .Y(n_21028));
 INVx1_ASAP7_75t_SL g28482 (.A(n_26130),
    .Y(n_21026));
 NOR2xp67_ASAP7_75t_SL g28491 (.A(n_21038),
    .B(n_26235),
    .Y(n_21042));
 XNOR2xp5_ASAP7_75t_SL g28492 (.A(n_21036),
    .B(n_26058),
    .Y(n_21038));
 XNOR2xp5_ASAP7_75t_SL g28496 (.A(n_21043),
    .B(n_21044),
    .Y(n_21045));
 NAND2xp5_ASAP7_75t_SL g28497 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(n_21043));
 NAND2xp5_ASAP7_75t_SL g28498 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .Y(n_21044));
 XNOR2x1_ASAP7_75t_SL g28499 (.B(n_21050),
    .Y(n_21051),
    .A(n_21047));
 XOR2xp5_ASAP7_75t_SL g285 (.A(n_4907),
    .B(n_14038),
    .Y(n_12050));
 INVxp67_ASAP7_75t_SL g28500 (.A(n_21046),
    .Y(n_21047));
 AOI21xp5_ASAP7_75t_SL g28501 (.A1(n_18983),
    .A2(n_11924),
    .B(n_11925),
    .Y(n_21046));
 XNOR2x1_ASAP7_75t_SL g28502 (.B(n_21049),
    .Y(n_21050),
    .A(n_21048));
 AND2x4_ASAP7_75t_SL g28503 (.A(n_2163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_552),
    .Y(n_21048));
 AND2x2_ASAP7_75t_SL g28504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_776),
    .B(n_2173),
    .Y(n_21049));
 XNOR2x1_ASAP7_75t_SL g28505 (.B(n_23015),
    .Y(n_21056),
    .A(n_21052));
 NAND2xp5_ASAP7_75t_SL g28508 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .Y(n_21058));
 OAI22xp5_ASAP7_75t_SL g28510 (.A1(n_21059),
    .A2(n_21064),
    .B1(n_21065),
    .B2(n_21066),
    .Y(n_21067));
 XNOR2xp5_ASAP7_75t_SL g28511 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_151),
    .B(n_20137),
    .Y(n_21059));
 MAJx2_ASAP7_75t_SL g28512 (.A(n_21203),
    .B(n_21061),
    .C(n_21204),
    .Y(n_21064));
 AOI21xp5_ASAP7_75t_SL g28514 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_128),
    .Y(n_21061));
 INVxp67_ASAP7_75t_SL g28516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_26),
    .Y(n_21062));
 INVx1_ASAP7_75t_SL g28517 (.A(n_21059),
    .Y(n_21065));
 INVx1_ASAP7_75t_SL g28518 (.A(n_21064),
    .Y(n_21066));
 NAND2x1_ASAP7_75t_SL g28519 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .Y(n_21069));
 OAI21x1_ASAP7_75t_SL g28523 (.A1(n_21071),
    .A2(n_21078),
    .B(n_21082),
    .Y(n_21083));
 NOR2xp33_ASAP7_75t_SL g28524 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_162),
    .Y(n_21071));
 OAI22xp5_ASAP7_75t_SL g28525 (.A1(n_21074),
    .A2(n_21075),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120),
    .B2(n_21077),
    .Y(n_21078));
 NAND2xp5_ASAP7_75t_SL g28526 (.A(n_21072),
    .B(n_21073),
    .Y(n_21074));
 OR2x2_ASAP7_75t_SL g28527 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_60),
    .Y(n_21072));
 INVx1_ASAP7_75t_SL g28528 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2),
    .Y(n_21073));
 NAND2xp5_ASAP7_75t_SL g28531 (.A(n_21072),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2),
    .Y(n_21077));
 AO21x1_ASAP7_75t_SL g28532 (.A1(n_21080),
    .A2(n_21081),
    .B(n_21072),
    .Y(n_21082));
 NAND2xp5_ASAP7_75t_SL g28533 (.A(n_21079),
    .B(n_21073),
    .Y(n_21080));
 NAND2xp33_ASAP7_75t_SL g28534 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2),
    .Y(n_21081));
 XNOR2x1_ASAP7_75t_SL g28540 (.B(n_21097),
    .Y(n_21098),
    .A(n_25303));
 NOR2xp33_ASAP7_75t_SL g28544 (.A(n_21091),
    .B(n_21092),
    .Y(n_21093));
 INVxp67_ASAP7_75t_SL g28545 (.A(n_9344),
    .Y(n_21091));
 XNOR2x1_ASAP7_75t_SL g28548 (.B(n_23664),
    .Y(n_21097),
    .A(n_5961));
 HB1xp67_ASAP7_75t_SL g28560 (.A(n_12948),
    .Y(n_21110));
 NAND2xp5_ASAP7_75t_SL g28561 (.A(n_21111),
    .B(n_21117),
    .Y(n_21118));
 MAJIxp5_ASAP7_75t_SL g28562 (.A(n_14880),
    .B(n_14881),
    .C(n_14887),
    .Y(n_21111));
 XNOR2xp5_ASAP7_75t_SL g28563 (.A(n_21113),
    .B(n_26131),
    .Y(n_21117));
 INVxp67_ASAP7_75t_SL g28564 (.A(n_21112),
    .Y(n_21113));
 MAJIxp5_ASAP7_75t_SL g28565 (.A(n_5744),
    .B(n_22159),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_145),
    .Y(n_21112));
 HB1xp67_ASAP7_75t_SL g28576 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_227),
    .Y(n_21129));
 XNOR2x1_ASAP7_75t_SL g28577 (.B(n_26132),
    .Y(n_21134),
    .A(n_21130));
 INVxp67_ASAP7_75t_SL g28578 (.A(n_15651),
    .Y(n_21130));
 MAJIxp5_ASAP7_75t_SL g28581 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_227),
    .Y(n_21131));
 XOR2xp5_ASAP7_75t_SL g28582 (.A(n_21135),
    .B(n_21136),
    .Y(n_21137));
 NAND2x1_ASAP7_75t_SL g28583 (.A(n_2173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_780),
    .Y(n_21135));
 NAND2xp5_ASAP7_75t_SL g28584 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_556),
    .B(n_2163),
    .Y(n_21136));
 XOR2xp5_ASAP7_75t_SL g28585 (.A(n_22178),
    .B(n_21141),
    .Y(n_21142));
 OAI21x1_ASAP7_75t_SL g28587 (.A1(n_21139),
    .A2(n_17019),
    .B(n_21140),
    .Y(n_21141));
 AND2x2_ASAP7_75t_SL g28588 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_589),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_685),
    .Y(n_21139));
 OR2x2_ASAP7_75t_SL g28589 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_589),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_685),
    .Y(n_21140));
 OAI21x1_ASAP7_75t_SL g28590 (.A1(n_21143),
    .A2(n_21148),
    .B(n_21151),
    .Y(n_21152));
 AND2x2_ASAP7_75t_SL g28591 (.A(n_20825),
    .B(n_4866),
    .Y(n_21143));
 NOR2x1_ASAP7_75t_SL g28592 (.A(n_7040),
    .B(n_21147),
    .Y(n_21148));
 INVx4_ASAP7_75t_SL g28593 (.A(n_21144),
    .Y(n_7040));
 AND2x4_ASAP7_75t_SL g28594 (.A(n_2163),
    .B(n_21663),
    .Y(n_21144));
 INVx2_ASAP7_75t_SL g28595 (.A(n_21146),
    .Y(n_21147));
 AND2x4_ASAP7_75t_SL g28596 (.A(n_2173),
    .B(n_19261),
    .Y(n_21146));
 NAND2xp5_ASAP7_75t_SL g28597 (.A(n_21147),
    .B(n_7040),
    .Y(n_21151));
 XNOR2xp5_ASAP7_75t_SL g286 (.A(n_10414),
    .B(n_20140),
    .Y(n_20141));
 XOR2x2_ASAP7_75t_SL g28605 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_167),
    .Y(n_21159));
 XOR2xp5_ASAP7_75t_SL g28606 (.A(n_21162),
    .B(n_21163),
    .Y(n_21164));
 XNOR2xp5_ASAP7_75t_SL g28607 (.A(n_21161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_143),
    .Y(n_21162));
 INVx1_ASAP7_75t_SL g28608 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_99),
    .Y(n_21161));
 MAJx2_ASAP7_75t_SL g28609 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_44),
    .Y(n_21163));
 MAJIxp5_ASAP7_75t_SL g28610 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_693),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_597),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_757),
    .Y(n_21165));
 XNOR2x1_ASAP7_75t_SL g28611 (.B(n_21166),
    .Y(n_21167),
    .A(n_16228));
 INVx2_ASAP7_75t_SL g28612 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_723),
    .Y(n_21166));
 INVxp67_ASAP7_75t_SL g28613 (.A(n_21167),
    .Y(n_21169));
 INVx1_ASAP7_75t_SL g28614 (.A(n_21165),
    .Y(n_21170));
 XNOR2x1_ASAP7_75t_SL g28616 (.B(n_26024),
    .Y(n_21177),
    .A(n_26133));
 NAND2xp5_ASAP7_75t_SL g28626 (.A(n_21183),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .Y(n_21184));
 OAI21xp33_ASAP7_75t_SL g28633 (.A1(n_21191),
    .A2(n_21192),
    .B(n_24176),
    .Y(n_21197));
 NAND2xp33_ASAP7_75t_SL g28634 (.A(n_5349),
    .B(n_5348),
    .Y(n_21191));
 AOI21xp33_ASAP7_75t_SL g28635 (.A1(n_23580),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_466),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_473),
    .Y(n_21192));
 XOR2xp5_ASAP7_75t_SL g28640 (.A(n_21198),
    .B(n_21199),
    .Y(n_21200));
 NAND2x1_ASAP7_75t_SL g28641 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .B(n_14523),
    .Y(n_21198));
 AND2x2_ASAP7_75t_SL g28642 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .Y(n_21199));
 INVx1_ASAP7_75t_SL g28643 (.A(n_21198),
    .Y(n_21201));
 XOR2xp5_ASAP7_75t_SL g28644 (.A(n_21203),
    .B(n_21204),
    .Y(n_21205));
 XNOR2x1_ASAP7_75t_SL g28645 (.B(n_9997),
    .Y(n_21203),
    .A(n_21202));
 HB1xp67_ASAP7_75t_SL g28646 (.A(n_22839),
    .Y(n_21202));
 XOR2xp5_ASAP7_75t_SL g28647 (.A(n_21062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_0),
    .Y(n_21204));
 XNOR2xp5_ASAP7_75t_SL g28649 (.A(n_21207),
    .B(n_25921),
    .Y(n_21210));
 OA22x2_ASAP7_75t_SL g28650 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_138),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_131),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_130),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_139),
    .Y(n_21207));
 NAND2x1p5_ASAP7_75t_SL g28654 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(n_3868),
    .Y(n_21212));
 OAI22xp5_ASAP7_75t_SL g28655 (.A1(n_9434),
    .A2(n_9432),
    .B1(n_18597),
    .B2(n_21214),
    .Y(n_21215));
 INVx1_ASAP7_75t_SL g28657 (.A(n_9434),
    .Y(n_21214));
 XNOR2xp5_ASAP7_75t_SL g28658 (.A(n_21217),
    .B(n_21218),
    .Y(n_21219));
 NAND2xp5_ASAP7_75t_SL g28659 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .Y(n_21217));
 NAND2x1_ASAP7_75t_SL g28660 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .B(n_2825),
    .Y(n_21218));
 INVx1_ASAP7_75t_SL g28661 (.A(n_21217),
    .Y(n_21220));
 NOR2xp67_ASAP7_75t_SL g28665 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_17),
    .Y(n_21222));
 NAND2xp5_ASAP7_75t_SL g28666 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_17),
    .Y(n_21224));
 XNOR2xp5_ASAP7_75t_SL g28667 (.A(n_26134),
    .B(n_21229),
    .Y(n_21230));
 MAJx2_ASAP7_75t_SL g28671 (.A(n_8498),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_172),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_186),
    .Y(n_21229));
 OAI22xp5_ASAP7_75t_SL g28681 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_54),
    .A2(n_21240),
    .B1(n_21241),
    .B2(n_8315),
    .Y(n_21242));
 NAND2x1_ASAP7_75t_SL g28682 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(n_22019),
    .Y(n_21240));
 INVx1_ASAP7_75t_SL g28683 (.A(n_21240),
    .Y(n_21241));
 MAJIxp5_ASAP7_75t_SL g28684 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_54),
    .B(n_21241),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_100),
    .Y(n_21243));
 MAJx2_ASAP7_75t_SL g28685 (.A(n_21245),
    .B(n_8959),
    .C(n_13678),
    .Y(n_21246));
 XNOR2x1_ASAP7_75t_SL g28686 (.B(n_21244),
    .Y(n_21245),
    .A(n_18929));
 HB1xp67_ASAP7_75t_SL g28687 (.A(n_9525),
    .Y(n_21244));
 XNOR2xp5_ASAP7_75t_SL g28688 (.A(n_21245),
    .B(n_16149),
    .Y(n_21247));
 MAJIxp5_ASAP7_75t_SL g28689 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_141),
    .B(n_21249),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_5),
    .Y(n_21250));
 INVx1_ASAP7_75t_SL g28690 (.A(n_21248),
    .Y(n_21249));
 NOR2x1_ASAP7_75t_SL g28691 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_62),
    .Y(n_21248));
 OAI22xp5_ASAP7_75t_SL g28692 (.A1(n_21249),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_128),
    .B1(n_21248),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_5),
    .Y(n_21251));
 NAND2xp5_ASAP7_75t_SL g28695 (.A(n_21254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_248),
    .Y(n_21255));
 HB1xp67_ASAP7_75t_SL g28696 (.A(n_24913),
    .Y(n_21254));
 OAI21xp33_ASAP7_75t_SL g28697 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_274),
    .A2(n_6354),
    .B(n_21254),
    .Y(n_21256));
 OAI21xp5_ASAP7_75t_SL g28698 (.A1(n_9200),
    .A2(n_9201),
    .B(n_21257),
    .Y(n_21258));
 AOI32xp33_ASAP7_75t_SL g28699 (.A1(n_9199),
    .A2(n_14355),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253),
    .B1(n_8145),
    .B2(n_9202),
    .Y(n_21257));
 INVxp67_ASAP7_75t_SL g287 (.A(n_19252),
    .Y(n_7487));
 AND2x2_ASAP7_75t_SL g28706 (.A(n_23975),
    .B(n_24684),
    .Y(n_21266));
 OAI22xp5_ASAP7_75t_SL g28707 (.A1(n_21267),
    .A2(n_9172),
    .B1(n_21268),
    .B2(n_21269),
    .Y(n_21270));
 NAND2xp5_ASAP7_75t_SL g28708 (.A(n_19645),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .Y(n_21267));
 INVx1_ASAP7_75t_SL g28709 (.A(n_21267),
    .Y(n_21268));
 INVx1_ASAP7_75t_SL g28710 (.A(n_9172),
    .Y(n_21269));
 MAJIxp5_ASAP7_75t_SL g28711 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_91),
    .B(n_21267),
    .C(n_9172),
    .Y(n_9584));
 OAI22xp5_ASAP7_75t_SL g28713 (.A1(n_21322),
    .A2(n_21277),
    .B1(n_10309),
    .B2(n_21276),
    .Y(n_21278));
 OAI21x1_ASAP7_75t_SL g28715 (.A1(n_26010),
    .A2(n_21282),
    .B(n_26107),
    .Y(n_21283));
 XNOR2xp5_ASAP7_75t_SL g28720 (.A(n_18930),
    .B(n_26135),
    .Y(n_21284));
 OAI22xp5_ASAP7_75t_SL g28721 (.A1(n_21285),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_201),
    .B1(n_21286),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_200),
    .Y(n_21287));
 XNOR2xp5_ASAP7_75t_SL g28722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_172),
    .B(n_10866),
    .Y(n_21285));
 MAJIxp5_ASAP7_75t_SL g28724 (.A(n_21288),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_201),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_210),
    .Y(n_21289));
 MAJIxp5_ASAP7_75t_SL g28726 (.A(n_19688),
    .B(n_21291),
    .C(n_12575),
    .Y(n_21293));
 INVx2_ASAP7_75t_SL g28727 (.A(n_21290),
    .Y(n_21291));
 MAJx2_ASAP7_75t_SL g28728 (.A(n_26098),
    .B(n_19453),
    .C(n_19454),
    .Y(n_21290));
 OAI22xp5_ASAP7_75t_SL g28730 (.A1(n_21291),
    .A2(n_21294),
    .B1(n_12575),
    .B2(n_21290),
    .Y(n_21295));
 INVx1_ASAP7_75t_SL g28731 (.A(n_12575),
    .Y(n_21294));
 OAI22xp5_ASAP7_75t_SL g28738 (.A1(n_21306),
    .A2(n_21307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_140),
    .B2(n_21308),
    .Y(n_21309));
 HB1xp67_ASAP7_75t_SL g28739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_3),
    .Y(n_21306));
 MAJIxp5_ASAP7_75t_SL g28740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_95),
    .B(n_15156),
    .C(n_9514),
    .Y(n_21307));
 MAJIxp5_ASAP7_75t_SL g28742 (.A(n_19686),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_140),
    .C(n_21308),
    .Y(n_21311));
 INVx1_ASAP7_75t_SL g28743 (.A(n_21307),
    .Y(n_21308));
 OAI21xp33_ASAP7_75t_SL g28749 (.A1(n_21317),
    .A2(n_22458),
    .B(n_13567),
    .Y(n_21318));
 NAND2xp5_ASAP7_75t_SL g28750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .B(n_8197),
    .Y(n_21317));
 NOR2xp33_ASAP7_75t_SL g28751 (.A(n_10311),
    .B(n_21317),
    .Y(n_21319));
 MAJx2_ASAP7_75t_SL g28754 (.A(n_9111),
    .B(n_22044),
    .C(n_13069),
    .Y(n_21322));
 XNOR2xp5_ASAP7_75t_SL g28763 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_153),
    .B(n_21331),
    .Y(n_21332));
 XNOR2xp5_ASAP7_75t_SL g28764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_61),
    .B(n_21200),
    .Y(n_21331));
 MAJIxp5_ASAP7_75t_SL g28765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_212),
    .B(n_21333),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_153),
    .Y(n_21334));
 INVxp67_ASAP7_75t_SRAM g28766 (.A(n_21331),
    .Y(n_21333));
 HB1xp67_ASAP7_75t_SL g28767 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_118),
    .Y(n_21335));
 MAJIxp5_ASAP7_75t_SL g28768 (.A(n_21338),
    .B(n_8573),
    .C(n_8572),
    .Y(n_21339));
 INVx1_ASAP7_75t_SL g28769 (.A(n_21337),
    .Y(n_21338));
 XNOR2xp5_ASAP7_75t_SL g28770 (.A(n_21336),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_148),
    .Y(n_21337));
 INVx1_ASAP7_75t_SL g28771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_118),
    .Y(n_21336));
 OAI22xp5_ASAP7_75t_SL g28772 (.A1(n_8567),
    .A2(n_21338),
    .B1(n_21337),
    .B2(n_8568),
    .Y(n_21340));
 XOR2x2_ASAP7_75t_SL g28782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_151),
    .B(n_21350),
    .Y(n_21351));
 XOR2xp5_ASAP7_75t_SL g28783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_41),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_86),
    .Y(n_21350));
 OAI22xp5_ASAP7_75t_SL g28784 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .A2(n_21354),
    .B1(n_21353),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_314),
    .Y(n_21355));
 INVx2_ASAP7_75t_SL g28785 (.A(n_21353),
    .Y(n_21354));
 XNOR2x1_ASAP7_75t_SL g28786 (.B(n_11916),
    .Y(n_21353),
    .A(n_21352));
 INVxp67_ASAP7_75t_SL g28787 (.A(n_17024),
    .Y(n_21352));
 MAJIxp5_ASAP7_75t_SL g28788 (.A(n_6453),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .C(n_21353),
    .Y(n_21357));
 AO21x2_ASAP7_75t_SL g28795 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_256),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_22),
    .B(n_21363),
    .Y(n_21364));
 NOR2xp33_ASAP7_75t_SL g28796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255),
    .Y(n_21363));
 AOI22xp33_ASAP7_75t_SL g28797 (.A1(n_21365),
    .A2(n_21367),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231),
    .Y(n_21368));
 INVxp67_ASAP7_75t_SL g28798 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231),
    .Y(n_21365));
 OAI21xp5_ASAP7_75t_SL g288 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_69),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113),
    .Y(n_7990));
 MAJIxp5_ASAP7_75t_SL g28800 (.A(n_21369),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_140),
    .C(n_7821),
    .Y(n_21370));
 XNOR2xp5_ASAP7_75t_SL g28801 (.A(n_6880),
    .B(n_6888),
    .Y(n_21369));
 XNOR2xp5_ASAP7_75t_SL g28802 (.A(n_21371),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_24),
    .Y(n_21372));
 INVxp67_ASAP7_75t_SL g28803 (.A(n_21369),
    .Y(n_21371));
 AO22x2_ASAP7_75t_SL g28804 (.A1(n_21374),
    .A2(n_22155),
    .B1(n_21375),
    .B2(n_21376),
    .Y(n_21377));
 NOR2xp33_ASAP7_75t_SL g28805 (.A(n_21373),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_280),
    .Y(n_21374));
 INVx1_ASAP7_75t_SL g28806 (.A(n_21789),
    .Y(n_21373));
 AND2x2_ASAP7_75t_SL g28807 (.A(n_21789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_280),
    .Y(n_21375));
 INVxp67_ASAP7_75t_SL g28808 (.A(n_22155),
    .Y(n_21376));
 XNOR2xp5_ASAP7_75t_SL g28809 (.A(n_21380),
    .B(n_21381),
    .Y(n_21382));
 AOI22xp5_ASAP7_75t_SL g28810 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110),
    .A2(n_21378),
    .B1(n_21379),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_154),
    .Y(n_21380));
 INVx1_ASAP7_75t_SL g28811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_154),
    .Y(n_21378));
 INVx1_ASAP7_75t_SL g28812 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110),
    .Y(n_21379));
 INVx1_ASAP7_75t_SL g28813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_143),
    .Y(n_21381));
 MAJIxp5_ASAP7_75t_SL g28814 (.A(n_21383),
    .B(n_21384),
    .C(n_21339),
    .Y(n_21385));
 OAI22xp5_ASAP7_75t_SL g28815 (.A1(n_21379),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_143),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110),
    .B2(n_21381),
    .Y(n_21383));
 HB1xp67_ASAP7_75t_SL g28816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_154),
    .Y(n_21384));
 XOR2xp5_ASAP7_75t_SL g28817 (.A(n_11638),
    .B(n_21390),
    .Y(n_21391));
 OAI22x1_ASAP7_75t_SL g28818 (.A1(n_7197),
    .A2(n_21386),
    .B1(n_21387),
    .B2(n_21388),
    .Y(n_21389));
 AND2x2_ASAP7_75t_SL g28819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_234),
    .B(n_7190),
    .Y(n_21386));
 HB1xp67_ASAP7_75t_SL g28821 (.A(n_7190),
    .Y(n_21388));
 NOR2x1_ASAP7_75t_SL g28822 (.A(n_11638),
    .B(n_21389),
    .Y(n_21392));
 NAND2xp5_ASAP7_75t_SL g28823 (.A(n_21389),
    .B(n_11638),
    .Y(n_21393));
 MAJIxp5_ASAP7_75t_SL g28824 (.A(n_20047),
    .B(n_20767),
    .C(n_21394),
    .Y(n_21395));
 NAND2xp67_ASAP7_75t_SL g28825 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .B(n_19411),
    .Y(n_21394));
 AOI22xp33_ASAP7_75t_SL g28828 (.A1(n_21398),
    .A2(n_21399),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_255),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_231),
    .Y(n_21400));
 INVxp67_ASAP7_75t_SL g28829 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_255),
    .Y(n_21398));
 INVx1_ASAP7_75t_SL g28830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_231),
    .Y(n_21399));
 AO22x2_ASAP7_75t_SL g28831 (.A1(n_21399),
    .A2(n_21398),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_256),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_22),
    .Y(n_21401));
 INVxp67_ASAP7_75t_SL g28833 (.A(n_22318),
    .Y(n_21404));
 INVx2_ASAP7_75t_SL g28838 (.A(n_22318),
    .Y(n_21407));
 OAI21xp5_ASAP7_75t_SL g28840 (.A1(n_21409),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_200),
    .Y(n_21410));
 NOR2xp67_ASAP7_75t_SL g28841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_168),
    .Y(n_21409));
 XOR2xp5_ASAP7_75t_SL g28842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_212),
    .B(n_21409),
    .Y(n_21413));
 XOR2x2_ASAP7_75t_SL g28845 (.A(n_21215),
    .B(n_21414),
    .Y(n_21415));
 INVx1_ASAP7_75t_SL g28846 (.A(n_21212),
    .Y(n_21414));
 MAJIxp5_ASAP7_75t_SL g28849 (.A(n_21419),
    .B(n_21420),
    .C(n_21421),
    .Y(n_21422));
 INVxp67_ASAP7_75t_SL g28850 (.A(n_22525),
    .Y(n_21420));
 MAJx2_ASAP7_75t_SL g28851 (.A(n_25426),
    .B(n_25427),
    .C(n_25425),
    .Y(n_21421));
 INVxp67_ASAP7_75t_SL g28852 (.A(n_21421),
    .Y(n_21423));
 NAND2xp5_ASAP7_75t_SL g28853 (.A(n_21425),
    .B(n_6758),
    .Y(n_21426));
 XNOR2xp5_ASAP7_75t_SL g28854 (.A(n_6896),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_250),
    .Y(n_21425));
 AOI221xp5_ASAP7_75t_SL g28855 (.A1(n_21427),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_233),
    .B1(n_6896),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_250),
    .C(n_6758),
    .Y(n_21429));
 NOR2x1_ASAP7_75t_SL g28862 (.A(n_9832),
    .B(n_24152),
    .Y(n_21434));
 OAI21xp5_ASAP7_75t_SL g28863 (.A1(n_20833),
    .A2(n_21436),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_84),
    .Y(n_21437));
 NOR2xp33_ASAP7_75t_SL g28864 (.A(n_21435),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_21436));
 OAI21xp5_ASAP7_75t_SL g28866 (.A1(n_23423),
    .A2(n_21438),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_84),
    .Y(n_21439));
 NOR2xp33_ASAP7_75t_SL g28867 (.A(n_21435),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .Y(n_21438));
 XNOR2xp5_ASAP7_75t_SL g28874 (.A(n_21447),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_143),
    .Y(n_21448));
 XNOR2xp5_ASAP7_75t_SL g28875 (.A(n_21446),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_154),
    .Y(n_21447));
 INVx1_ASAP7_75t_SL g28876 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_110),
    .Y(n_21446));
 MAJIxp5_ASAP7_75t_SL g28877 (.A(n_21450),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_223),
    .Y(n_21452));
 OAI22xp5_ASAP7_75t_SL g28878 (.A1(n_21446),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_143),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_110),
    .B2(n_21449),
    .Y(n_21450));
 INVxp67_ASAP7_75t_SL g28879 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_143),
    .Y(n_21449));
 MAJx2_ASAP7_75t_SL g28884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_81),
    .C(n_7269),
    .Y(n_21454));
 NOR2xp33_ASAP7_75t_SL g28886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_113),
    .B(n_21454),
    .Y(n_21458));
 NAND2xp33_ASAP7_75t_SRAM g28887 (.A(n_21454),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_113),
    .Y(n_21459));
 XNOR2x1_ASAP7_75t_SL g28888 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_189),
    .Y(n_21462),
    .A(n_21461));
 XNOR2x1_ASAP7_75t_SL g28889 (.B(n_22028),
    .Y(n_21461),
    .A(n_21460));
 INVxp67_ASAP7_75t_SL g28890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_104),
    .Y(n_21460));
 MAJIxp5_ASAP7_75t_SL g28891 (.A(n_21463),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_132),
    .Y(n_21464));
 INVx1_ASAP7_75t_SL g28892 (.A(n_21461),
    .Y(n_21463));
 MAJx2_ASAP7_75t_SL g28893 (.A(n_21918),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_118),
    .C(n_21467),
    .Y(n_21469));
 MAJIxp5_ASAP7_75t_SL g28897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_93),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_63),
    .Y(n_21467));
 MAJIxp5_ASAP7_75t_SL g289 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_207),
    .B(n_18701),
    .C(n_11444),
    .Y(n_20140));
 NOR3xp33_ASAP7_75t_SL g28900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_286),
    .B(n_11869),
    .C(n_11343),
    .Y(n_21471));
 INVxp67_ASAP7_75t_SL g28901 (.A(n_21473),
    .Y(n_21474));
 NAND2x1_ASAP7_75t_SL g28902 (.A(n_7489),
    .B(n_11120),
    .Y(n_21473));
 OAI21xp5_ASAP7_75t_SL g28903 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302),
    .A2(n_7491),
    .B(n_21475),
    .Y(n_21476));
 HB1xp67_ASAP7_75t_SL g28904 (.A(n_21473),
    .Y(n_21475));
 OAI21xp5_ASAP7_75t_SL g28905 (.A1(n_21473),
    .A2(n_19917),
    .B(n_19918),
    .Y(n_21477));
 NAND2xp5_ASAP7_75t_SL g28906 (.A(n_21478),
    .B(n_19191),
    .Y(n_21479));
 XNOR2xp5_ASAP7_75t_SL g28907 (.A(n_23549),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_377),
    .Y(n_21478));
 NOR2xp67_ASAP7_75t_SL g28908 (.A(n_19191),
    .B(n_21478),
    .Y(n_21480));
 AOI21xp5_ASAP7_75t_SL g28909 (.A1(n_21481),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_243),
    .Y(n_21482));
 XOR2x1_ASAP7_75t_SL g28910 (.A(n_18945),
    .Y(n_21481),
    .B(n_9041));
 XNOR2xp5_ASAP7_75t_SL g28911 (.A(n_9605),
    .B(n_21481),
    .Y(n_21483));
 XOR2xp5_ASAP7_75t_SL g28912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_231),
    .B(n_21485),
    .Y(n_21486));
 HB1xp67_ASAP7_75t_SL g28913 (.A(n_21484),
    .Y(n_21485));
 MAJIxp5_ASAP7_75t_SL g28914 (.A(n_10520),
    .B(n_6871),
    .C(n_6872),
    .Y(n_21484));
 OAI21x1_ASAP7_75t_SL g28916 (.A1(n_21484),
    .A2(n_6479),
    .B(n_6480),
    .Y(n_21487));
 XNOR2xp5_ASAP7_75t_SL g28918 (.A(n_11243),
    .B(n_9893),
    .Y(n_21489));
 HB1xp67_ASAP7_75t_SL g28921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_118),
    .Y(n_21493));
 XNOR2xp5_ASAP7_75t_SL g28922 (.A(n_11771),
    .B(n_21496),
    .Y(n_21497));
 OAI22xp5_ASAP7_75t_SL g28923 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_118),
    .A2(n_12278),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_55),
    .B2(n_21495),
    .Y(n_21496));
 INVx1_ASAP7_75t_SL g28925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_118),
    .Y(n_21495));
 XOR2xp5_ASAP7_75t_SL g28930 (.A(n_14106),
    .B(n_22948),
    .Y(n_21503));
 XOR2x2_ASAP7_75t_SL g28932 (.A(n_21504),
    .B(n_13233),
    .Y(n_21505));
 OAI22xp5_ASAP7_75t_SL g28933 (.A1(n_19407),
    .A2(n_9818),
    .B1(n_19408),
    .B2(n_20008),
    .Y(n_21504));
 A2O1A1O1Ixp25_ASAP7_75t_SL g28934 (.A1(n_21506),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_273),
    .C(n_11966),
    .D(n_11968),
    .Y(n_21507));
 NAND2xp5_ASAP7_75t_SL g28935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_242),
    .Y(n_21506));
 AOI21x1_ASAP7_75t_SL g28936 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_290),
    .A2(n_21506),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_273),
    .Y(n_21508));
 NAND2xp5_ASAP7_75t_SL g28937 (.A(n_21506),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_274),
    .Y(n_21509));
 MAJIxp5_ASAP7_75t_SL g28938 (.A(n_12286),
    .B(n_12039),
    .C(n_21510),
    .Y(n_21511));
 NAND2xp5_ASAP7_75t_SL g28939 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .Y(n_21510));
 XNOR2xp5_ASAP7_75t_SL g28940 (.A(n_21512),
    .B(n_12285),
    .Y(n_21513));
 INVxp67_ASAP7_75t_SL g28941 (.A(n_21510),
    .Y(n_21512));
 AO21x2_ASAP7_75t_SL g28942 (.A1(n_21516),
    .A2(n_21517),
    .B(n_21518),
    .Y(n_21519));
 NOR2xp33_ASAP7_75t_SL g28943 (.A(n_21515),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_301),
    .Y(n_21516));
 NAND2xp5_ASAP7_75t_SL g28944 (.A(n_18577),
    .B(n_21514),
    .Y(n_21515));
 INVxp67_ASAP7_75t_SL g28945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_213),
    .Y(n_21514));
 INVxp67_ASAP7_75t_SRAM g28946 (.A(n_11235),
    .Y(n_21517));
 OAI32xp33_ASAP7_75t_SL g28947 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_298),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_301),
    .A3(n_21515),
    .B1(n_21515),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_211),
    .Y(n_21518));
 XNOR2xp5_ASAP7_75t_SL g28949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_112),
    .B(n_26139),
    .Y(n_21524));
 AOI21x1_ASAP7_75t_SL g28953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_309),
    .A2(n_21830),
    .B(n_21526),
    .Y(n_21527));
 INVxp67_ASAP7_75t_SL g28954 (.A(n_21847),
    .Y(n_21526));
 XNOR2xp5_ASAP7_75t_SL g28957 (.A(n_8418),
    .B(n_21529),
    .Y(n_21530));
 XOR2xp5_ASAP7_75t_SL g28958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_168),
    .B(n_12516),
    .Y(n_21529));
 MAJx2_ASAP7_75t_SL g28959 (.A(n_21531),
    .B(n_21532),
    .C(n_12520),
    .Y(n_21534));
 INVxp67_ASAP7_75t_SRAM g28960 (.A(n_21529),
    .Y(n_21531));
 INVx1_ASAP7_75t_SL g28961 (.A(n_12518),
    .Y(n_21532));
 NAND2xp5_ASAP7_75t_SL g28968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_296),
    .B(n_21827),
    .Y(n_21541));
 OAI22xp5_ASAP7_75t_SL g28971 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_86),
    .A2(n_21544),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_85),
    .B2(n_21543),
    .Y(n_21545));
 MAJx2_ASAP7_75t_SL g28973 (.A(n_9535),
    .B(n_20591),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_108),
    .Y(n_21543));
 NAND2xp5_ASAP7_75t_SL g28979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_229),
    .B(n_21551),
    .Y(n_21552));
 XNOR2x2_ASAP7_75t_SL g28980 (.A(n_14880),
    .B(n_14883),
    .Y(n_21551));
 NOR2xp67_ASAP7_75t_SL g28982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_229),
    .B(n_21551),
    .Y(n_21554));
 AOI21xp5_ASAP7_75t_SL g28984 (.A1(n_21556),
    .A2(n_21557),
    .B(n_7117),
    .Y(n_21559));
 NAND2xp5_ASAP7_75t_SL g28985 (.A(n_7746),
    .B(n_7523),
    .Y(n_21556));
 OR2x2_ASAP7_75t_SL g28986 (.A(n_7746),
    .B(n_7523),
    .Y(n_21557));
 NAND3xp33_ASAP7_75t_SL g28988 (.A(n_21557),
    .B(n_21556),
    .C(n_7117),
    .Y(n_21560));
 OAI22xp5_ASAP7_75t_SL g28998 (.A1(n_21570),
    .A2(n_9675),
    .B1(n_21571),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_54),
    .Y(n_21572));
 NAND2xp5_ASAP7_75t_SL g28999 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .Y(n_21570));
 XOR2xp5_ASAP7_75t_SL g29 (.A(n_12580),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_171),
    .Y(n_5339));
 XNOR2xp5_ASAP7_75t_SL g290 (.A(n_5811),
    .B(n_18848),
    .Y(n_5815));
 INVx1_ASAP7_75t_SL g29000 (.A(n_21570),
    .Y(n_21571));
 MAJIxp5_ASAP7_75t_SL g29001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_54),
    .B(n_21571),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_100),
    .Y(n_21573));
 AOI21x1_ASAP7_75t_SL g29005 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_290),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_273),
    .Y(n_21577));
 OAI22xp5_ASAP7_75t_SL g29006 (.A1(n_21578),
    .A2(n_12649),
    .B1(n_12648),
    .B2(n_21579),
    .Y(n_21580));
 XNOR2x1_ASAP7_75t_SL g29007 (.B(n_11108),
    .Y(n_21578),
    .A(n_26175));
 INVx1_ASAP7_75t_SL g29008 (.A(n_21578),
    .Y(n_21579));
 NAND2xp33_ASAP7_75t_SL g29009 (.A(n_21578),
    .B(n_12648),
    .Y(n_21581));
 NOR2xp33_ASAP7_75t_SL g29010 (.A(n_21578),
    .B(n_12648),
    .Y(n_21582));
 NAND2x1_ASAP7_75t_SL g29013 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(n_2922),
    .Y(n_21583));
 MAJIxp5_ASAP7_75t_SL g29016 (.A(n_22733),
    .B(n_21583),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_99),
    .Y(n_21588));
 AOI21x1_ASAP7_75t_SL g29022 (.A1(n_9456),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_319),
    .B(n_11178),
    .Y(n_21593));
 XNOR2xp5_ASAP7_75t_SL g29023 (.A(n_18716),
    .B(n_21593),
    .Y(n_21595));
 HB1xp67_ASAP7_75t_SL g29025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_281),
    .Y(n_21596));
 OAI22xp5_ASAP7_75t_SL g29026 (.A1(n_26224),
    .A2(n_21599),
    .B1(n_21600),
    .B2(n_21598),
    .Y(n_21601));
 INVx1_ASAP7_75t_SL g29027 (.A(n_21598),
    .Y(n_21599));
 MAJx2_ASAP7_75t_SL g29028 (.A(n_10355),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_13),
    .C(n_9549),
    .Y(n_21598));
 INVx2_ASAP7_75t_SL g29032 (.A(n_26224),
    .Y(n_21600));
 MAJIxp5_ASAP7_75t_SL g29034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_64),
    .B(n_21606),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_35),
    .Y(n_21607));
 NAND2xp5_ASAP7_75t_SL g29035 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .Y(n_21606));
 XNOR2xp5_ASAP7_75t_SL g29039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_188),
    .B(n_21611),
    .Y(n_21612));
 XNOR2xp5_ASAP7_75t_SL g29040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_124),
    .Y(n_21611));
 MAJIxp5_ASAP7_75t_SL g29041 (.A(n_21611),
    .B(n_13021),
    .C(n_13023),
    .Y(n_21613));
 XNOR2xp5_ASAP7_75t_SL g29043 (.A(n_26128),
    .B(n_26141),
    .Y(n_21617));
 XNOR2x1_ASAP7_75t_SL g29047 (.B(n_21620),
    .Y(n_21621),
    .A(n_21619));
 XNOR2x1_ASAP7_75t_SL g29048 (.B(n_9862),
    .Y(n_21619),
    .A(n_9860));
 INVx1_ASAP7_75t_SL g29049 (.A(n_19248),
    .Y(n_21620));
 OAI21xp5_ASAP7_75t_SL g29051 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_252),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_251),
    .B(n_21623),
    .Y(n_21624));
 NAND2xp5_ASAP7_75t_SL g29052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_236),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_207),
    .Y(n_21623));
 NAND2xp5_ASAP7_75t_SL g29053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_253),
    .B(n_21625),
    .Y(n_21626));
 HB1xp67_ASAP7_75t_SL g29054 (.A(n_21623),
    .Y(n_21625));
 MAJIxp5_ASAP7_75t_SL g29055 (.A(n_21628),
    .B(n_21629),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_131),
    .Y(n_21630));
 INVx1_ASAP7_75t_SL g29056 (.A(n_21627),
    .Y(n_21628));
 XNOR2x1_ASAP7_75t_SL g29057 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_8),
    .Y(n_21627),
    .A(n_13637));
 HB1xp67_ASAP7_75t_SL g29058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_147),
    .Y(n_21629));
 XNOR2xp5_ASAP7_75t_SL g29059 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_181),
    .B(n_21627),
    .Y(n_21631));
 OAI22xp5_ASAP7_75t_SL g29060 (.A1(n_21632),
    .A2(n_13036),
    .B1(n_21633),
    .B2(n_13038),
    .Y(n_21634));
 MAJIxp5_ASAP7_75t_SL g29061 (.A(n_12956),
    .B(n_19190),
    .C(n_14383),
    .Y(n_21632));
 INVx1_ASAP7_75t_SL g29062 (.A(n_21632),
    .Y(n_21633));
 OAI21xp5_ASAP7_75t_SL g29063 (.A1(n_21635),
    .A2(n_13034),
    .B(n_21636),
    .Y(n_21637));
 AND2x2_ASAP7_75t_SL g29064 (.A(n_21632),
    .B(n_13038),
    .Y(n_21635));
 OR2x2_ASAP7_75t_SL g29065 (.A(n_21632),
    .B(n_13038),
    .Y(n_21636));
 MAJx2_ASAP7_75t_SL g29068 (.A(n_21643),
    .B(n_11726),
    .C(n_5641),
    .Y(n_21644));
 XNOR2xp5_ASAP7_75t_SL g29069 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_747),
    .B(n_26142),
    .Y(n_21643));
 XOR2xp5_ASAP7_75t_SL g29073 (.A(n_21645),
    .B(n_6141),
    .Y(n_21646));
 HB1xp67_ASAP7_75t_SL g29074 (.A(n_21643),
    .Y(n_21645));
 XNOR2xp5_ASAP7_75t_SL g29078 (.A(n_22034),
    .B(n_21650),
    .Y(n_21651));
 AOI22xp5_ASAP7_75t_SL g29079 (.A1(n_18843),
    .A2(n_21648),
    .B1(n_21649),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_19),
    .Y(n_21650));
 INVx1_ASAP7_75t_SL g29080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_19),
    .Y(n_21648));
 AND2x2_ASAP7_75t_SL g29082 (.A(n_21651),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_243),
    .Y(n_21654));
 HB1xp67_ASAP7_75t_SL g29083 (.A(n_21666),
    .Y(n_21667));
 OAI22xp5_ASAP7_75t_SL g29084 (.A1(n_21664),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_157),
    .B1(n_21665),
    .B2(n_23423),
    .Y(n_21666));
 XOR2x2_ASAP7_75t_SL g29085 (.A(n_26252),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_609),
    .Y(n_21664));
 XNOR2xp5_ASAP7_75t_SL g29086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_42),
    .B(n_21666),
    .Y(n_21669));
 OAI22xp5_ASAP7_75t_SL g29089 (.A1(n_21664),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_162),
    .B1(n_20833),
    .B2(n_21665),
    .Y(n_21673));
 XNOR2x1_ASAP7_75t_SL g29090 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_207),
    .Y(n_21678),
    .A(n_21677));
 OAI22xp5_ASAP7_75t_SL g29091 (.A1(n_21676),
    .A2(n_10982),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_156),
    .B2(n_21675),
    .Y(n_21677));
 XNOR2xp5_ASAP7_75t_SL g29093 (.A(n_25978),
    .B(n_22052),
    .Y(n_21675));
 MAJx2_ASAP7_75t_SL g29096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_207),
    .B(n_21685),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_156),
    .Y(n_21686));
 INVxp67_ASAP7_75t_SL g29097 (.A(n_21684),
    .Y(n_21685));
 XNOR2xp5_ASAP7_75t_SL g29098 (.A(n_25984),
    .B(n_26143),
    .Y(n_21684));
 MAJIxp5_ASAP7_75t_SL g291 (.A(n_23461),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_75),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_76),
    .Y(n_23467));
 OAI21xp5_ASAP7_75t_SL g29104 (.A1(n_21684),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_156),
    .B(n_21689),
    .Y(n_21690));
 NAND2xp5_ASAP7_75t_L g29105 (.A(n_21684),
    .B(n_21688),
    .Y(n_21689));
 INVxp67_ASAP7_75t_SL g29106 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_155),
    .Y(n_21688));
 OAI22xp5_ASAP7_75t_SL g29108 (.A1(n_20625),
    .A2(n_21691),
    .B1(n_20624),
    .B2(n_20621),
    .Y(n_21692));
 NOR2xp33_ASAP7_75t_SL g29109 (.A(n_3681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .Y(n_21691));
 NAND2x1_ASAP7_75t_SL g29110 (.A(n_2181),
    .B(n_21696),
    .Y(n_21697));
 XNOR2xp5_ASAP7_75t_SL g29111 (.A(n_21694),
    .B(n_23124),
    .Y(n_21696));
 INVxp67_ASAP7_75t_SL g29112 (.A(n_11216),
    .Y(n_21694));
 OAI21xp5_ASAP7_75t_SL g29114 (.A1(n_21698),
    .A2(n_23124),
    .B(n_11215),
    .Y(n_21699));
 HB1xp67_ASAP7_75t_SL g29115 (.A(n_11869),
    .Y(n_21698));
 MAJx2_ASAP7_75t_SL g292 (.A(n_21913),
    .B(n_20589),
    .C(n_22499),
    .Y(n_23461));
 AND3x4_ASAP7_75t_SL g29200 (.A(n_2146),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .C(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[1]),
    .Y(n_21789));
 MAJIxp5_ASAP7_75t_SL g29201 (.A(n_13031),
    .B(n_7932),
    .C(n_25971),
    .Y(n_21793));
 XOR2xp5_ASAP7_75t_SL g29205 (.A(n_25971),
    .B(n_13031),
    .Y(n_21795));
 XNOR2x1_ASAP7_75t_SL g29206 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_194),
    .Y(n_21796),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_9));
 AND2x2_ASAP7_75t_L g29207 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_6965),
    .Y(n_21797));
 XNOR2x1_ASAP7_75t_SL g29212 (.B(n_15720),
    .Y(n_21802),
    .A(n_12834));
 XOR2xp5_ASAP7_75t_SL g29213 (.A(n_21803),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_114),
    .Y(n_21804));
 INVx2_ASAP7_75t_SL g29232 (.A(n_21829),
    .Y(n_21830));
 AOI21x1_ASAP7_75t_SL g29233 (.A1(n_21826),
    .A2(n_21827),
    .B(n_21828),
    .Y(n_21829));
 AO21x1_ASAP7_75t_SL g29234 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_266),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_277),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_264),
    .Y(n_21826));
 NAND2x1_ASAP7_75t_SL g29235 (.A(n_3246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_248),
    .Y(n_21827));
 MAJIxp5_ASAP7_75t_SL g29240 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_234),
    .B(n_2939),
    .C(n_3547),
    .Y(n_21832));
 NAND2xp5_ASAP7_75t_SL g29241 (.A(n_21835),
    .B(n_21836),
    .Y(n_21837));
 NAND2xp5_ASAP7_75t_SL g29242 (.A(n_10472),
    .B(n_21482),
    .Y(n_21835));
 NAND2xp5_ASAP7_75t_SL g29243 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_258),
    .B(n_21483),
    .Y(n_21836));
 OAI21xp5_ASAP7_75t_SL g29244 (.A1(n_21838),
    .A2(n_21839),
    .B(n_21840),
    .Y(n_21841));
 AOI21xp5_ASAP7_75t_SL g29245 (.A1(n_14059),
    .A2(n_14061),
    .B(n_14067),
    .Y(n_21838));
 NOR2xp33_ASAP7_75t_SL g29246 (.A(n_14061),
    .B(n_14059),
    .Y(n_21839));
 OAI21xp5_ASAP7_75t_SL g29247 (.A1(n_22335),
    .A2(n_21847),
    .B(n_21852),
    .Y(n_21853));
 AOI21xp5_ASAP7_75t_SL g29249 (.A1(n_21845),
    .A2(n_21835),
    .B(n_21846),
    .Y(n_21847));
 NOR2xp67_ASAP7_75t_SL g29250 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_258),
    .B(n_21483),
    .Y(n_21845));
 NOR2xp67_ASAP7_75t_SL g29251 (.A(n_21482),
    .B(n_10472),
    .Y(n_21846));
 AOI31xp33_ASAP7_75t_SL g29252 (.A1(n_21841),
    .A2(n_21848),
    .A3(n_21849),
    .B(n_21851),
    .Y(n_21852));
 INVx1_ASAP7_75t_SL g29254 (.A(n_21832),
    .Y(n_21849));
 NOR3xp33_ASAP7_75t_SL g29255 (.A(n_21840),
    .B(n_21838),
    .C(n_21850),
    .Y(n_21851));
 XNOR2xp5_ASAP7_75t_SL g29256 (.A(n_21859),
    .B(n_21866),
    .Y(n_21867));
 MAJIxp5_ASAP7_75t_SL g29257 (.A(n_21855),
    .B(n_21856),
    .C(n_21858),
    .Y(n_21859));
 NAND2xp5_ASAP7_75t_SL g29258 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .B(n_15201),
    .Y(n_21855));
 NAND2x1_ASAP7_75t_SL g29259 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(n_18039),
    .Y(n_21856));
 INVx1_ASAP7_75t_SL g29260 (.A(n_21857),
    .Y(n_21858));
 NAND2x1p5_ASAP7_75t_SL g29261 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .B(n_3218),
    .Y(n_21857));
 XNOR2xp5_ASAP7_75t_SL g29262 (.A(n_21862),
    .B(n_21865),
    .Y(n_21866));
 NAND2xp33_ASAP7_75t_SL g29263 (.A(n_21861),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(n_21862));
 XNOR2xp5_ASAP7_75t_SL g29265 (.A(n_21863),
    .B(n_21864),
    .Y(n_21865));
 NAND2x1_ASAP7_75t_SL g29266 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .B(n_18031),
    .Y(n_21863));
 NAND2x1_ASAP7_75t_SL g29267 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(n_4831),
    .Y(n_21864));
 INVxp67_ASAP7_75t_SL g29268 (.A(n_21863),
    .Y(n_21869));
 INVx1_ASAP7_75t_SL g29272 (.A(n_22739),
    .Y(n_21873));
 NOR3x1_ASAP7_75t_SL g29277 (.A(n_25128),
    .B(n_4843),
    .C(n_17443),
    .Y(n_21875));
 OAI21xp5_ASAP7_75t_SL g29278 (.A1(n_10627),
    .A2(n_25128),
    .B(n_25881),
    .Y(n_21876));
 NAND2xp5_ASAP7_75t_SL g29281 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_362),
    .B(n_10264),
    .Y(n_21880));
 NOR2xp33_ASAP7_75t_SL g29282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_362),
    .B(n_10264),
    .Y(n_21882));
 INVxp67_ASAP7_75t_SL g293 (.A(n_14733),
    .Y(n_14734));
 XNOR2xp5_ASAP7_75t_SL g29304 (.A(n_21911),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_18),
    .Y(n_21912));
 NAND2xp5_ASAP7_75t_SL g29305 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_3317),
    .Y(n_21911));
 AND2x2_ASAP7_75t_SL g29307 (.A(n_19370),
    .B(n_10141),
    .Y(n_21913));
 XOR2xp5_ASAP7_75t_SL g29308 (.A(n_26145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_26),
    .Y(n_21918));
 XNOR2x1_ASAP7_75t_SL g29313 (.B(n_21919),
    .Y(n_21920),
    .A(n_5784));
 INVx2_ASAP7_75t_SL g29314 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_743),
    .Y(n_21919));
 OAI22xp5_ASAP7_75t_SL g29315 (.A1(n_21922),
    .A2(n_21923),
    .B1(n_12750),
    .B2(n_21924),
    .Y(n_21925));
 AND2x2_ASAP7_75t_SL g29316 (.A(n_7638),
    .B(n_7637),
    .Y(n_21922));
 OR2x2_ASAP7_75t_SL g29317 (.A(n_12752),
    .B(n_7644),
    .Y(n_21923));
 AOI21xp5_ASAP7_75t_SL g29318 (.A1(n_7637),
    .A2(n_7638),
    .B(n_7644),
    .Y(n_21924));
 OAI21xp5_ASAP7_75t_SL g29320 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_196),
    .A2(n_21926),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_200),
    .Y(n_21927));
 NOR2xp67_ASAP7_75t_SL g29321 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_122),
    .B(n_10212),
    .Y(n_21926));
 XNOR2xp5_ASAP7_75t_SL g29322 (.A(n_21929),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_18),
    .Y(n_21930));
 NAND2x1_ASAP7_75t_SL g29323 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(n_3317),
    .Y(n_21929));
 MAJIxp5_ASAP7_75t_SL g29324 (.A(n_3806),
    .B(n_21931),
    .C(n_18720),
    .Y(n_21932));
 NAND2xp5_ASAP7_75t_SL g29325 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .Y(n_21931));
 XNOR2xp5_ASAP7_75t_SL g29329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_106),
    .B(n_21936),
    .Y(n_21937));
 NAND2xp5_ASAP7_75t_L g29330 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .Y(n_21936));
 AND2x2_ASAP7_75t_SL g29333 (.A(n_19866),
    .B(n_6323),
    .Y(n_21939));
 OAI21xp5_ASAP7_75t_SL g29334 (.A1(n_21941),
    .A2(n_8945),
    .B(n_21943),
    .Y(n_21944));
 AND2x2_ASAP7_75t_SL g29335 (.A(n_6576),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .Y(n_21941));
 NAND2xp5_ASAP7_75t_SL g29336 (.A(n_21942),
    .B(n_21941),
    .Y(n_21943));
 INVx1_ASAP7_75t_SL g29337 (.A(n_8943),
    .Y(n_21942));
 MAJIxp5_ASAP7_75t_SL g29338 (.A(n_21946),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_145),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_188),
    .Y(n_21947));
 HB1xp67_ASAP7_75t_SL g29339 (.A(n_21945),
    .Y(n_21946));
 XNOR2xp5_ASAP7_75t_SL g29340 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_721),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_8),
    .Y(n_21945));
 NAND2xp5_ASAP7_75t_SL g29342 (.A(n_21948),
    .B(n_21357),
    .Y(n_21949));
 XNOR2xp5_ASAP7_75t_SL g29343 (.A(n_12077),
    .B(n_14452),
    .Y(n_21948));
 XNOR2xp5_ASAP7_75t_SL g29345 (.A(n_21952),
    .B(n_26080),
    .Y(n_21956));
 INVx1_ASAP7_75t_SL g29346 (.A(n_4487),
    .Y(n_21952));
 AOI21x1_ASAP7_75t_SL g29353 (.A1(n_21960),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_310),
    .B(n_13953),
    .Y(n_21961));
 AND2x2_ASAP7_75t_SL g29354 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_304),
    .B(n_19281),
    .Y(n_21960));
 AND2x2_ASAP7_75t_SL g29355 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_314),
    .B(n_18769),
    .Y(n_21962));
 XNOR2xp5_ASAP7_75t_SL g29356 (.A(n_21967),
    .B(n_8951),
    .Y(n_21968));
 OAI21x1_ASAP7_75t_SL g29357 (.A1(n_10618),
    .A2(n_21965),
    .B(n_21966),
    .Y(n_21967));
 AND2x2_ASAP7_75t_SL g29358 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115),
    .B(n_4341),
    .Y(n_21965));
 OR2x2_ASAP7_75t_SL g29360 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115),
    .B(n_4341),
    .Y(n_21966));
 XNOR2xp5_ASAP7_75t_SL g29362 (.A(n_21970),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_167),
    .Y(n_21971));
 XOR2xp5_ASAP7_75t_SL g29363 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_38),
    .Y(n_21970));
 XOR2xp5_ASAP7_75t_SL g29364 (.A(n_21973),
    .B(n_26041),
    .Y(n_21974));
 INVxp67_ASAP7_75t_SL g29365 (.A(n_21972),
    .Y(n_21973));
 MAJIxp5_ASAP7_75t_SL g29366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_141),
    .C(n_8852),
    .Y(n_21972));
 MAJIxp5_ASAP7_75t_SL g29368 (.A(n_21977),
    .B(n_13590),
    .C(n_20413),
    .Y(n_21978));
 AND2x2_ASAP7_75t_SL g29369 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_610),
    .B(n_9661),
    .Y(n_21977));
 OAI21x1_ASAP7_75t_SL g29370 (.A1(n_21979),
    .A2(n_8975),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_200),
    .Y(n_21980));
 NOR2xp67_ASAP7_75t_SL g29371 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_179),
    .Y(n_21979));
 NOR2xp67_ASAP7_75t_SL g29374 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_231),
    .B(n_21983),
    .Y(n_21984));
 XNOR2xp5_ASAP7_75t_SL g29375 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_10),
    .B(n_20400),
    .Y(n_21983));
 MAJIxp5_ASAP7_75t_SL g29376 (.A(n_21985),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_206),
    .C(n_10086),
    .Y(n_21986));
 XNOR2x1_ASAP7_75t_SL g29377 (.B(n_21000),
    .Y(n_21985),
    .A(n_20997));
 NAND2x1_ASAP7_75t_SL g29378 (.A(n_21987),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_71),
    .Y(n_21988));
 NAND2xp5_ASAP7_75t_SL g29379 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(n_14987),
    .Y(n_21987));
 NAND2x1_ASAP7_75t_SL g29380 (.A(n_21990),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .Y(n_21991));
 MAJIxp5_ASAP7_75t_L g29383_dup (.A(n_22712),
    .B(n_22713),
    .C(n_22714),
    .Y(n_22717));
 XNOR2xp5_ASAP7_75t_SL g29386 (.A(n_21621),
    .B(n_21995),
    .Y(n_21996));
 XNOR2xp5_ASAP7_75t_SL g29387 (.A(n_23665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_24),
    .Y(n_21995));
 MAJx2_ASAP7_75t_SL g29388 (.A(n_21997),
    .B(n_21998),
    .C(n_21999),
    .Y(n_22000));
 INVx1_ASAP7_75t_SL g29389 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_653),
    .Y(n_21997));
 MAJIxp5_ASAP7_75t_SL g29390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_783),
    .B(n_6114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_559),
    .Y(n_21998));
 MAJIxp5_ASAP7_75t_SL g29392 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_779),
    .B(n_5800),
    .C(n_22001),
    .Y(n_22002));
 AND2x2_ASAP7_75t_SL g29393 (.A(n_12781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_714),
    .Y(n_22001));
 XOR2xp5_ASAP7_75t_SL g29394 (.A(n_22004),
    .B(n_4480),
    .Y(n_22005));
 XNOR2xp5_ASAP7_75t_SL g29395 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_5),
    .B(n_22003),
    .Y(n_22004));
 INVx1_ASAP7_75t_SL g29396 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_127),
    .Y(n_22003));
 XOR2xp5_ASAP7_75t_SL g294 (.A(n_24678),
    .B(n_24679),
    .Y(n_24680));
 NAND2xp5_ASAP7_75t_SL g29402 (.A(n_22011),
    .B(n_21880),
    .Y(n_22012));
 NAND2xp5_ASAP7_75t_SL g29403 (.A(n_11961),
    .B(n_10267),
    .Y(n_22011));
 XNOR2x1_ASAP7_75t_SL g29404 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_153),
    .Y(n_22016),
    .A(n_13597));
 XNOR2x1_ASAP7_75t_SL g29405 (.B(n_13593),
    .Y(n_13597),
    .A(n_22732));
 AND2x2_ASAP7_75t_SL g29408 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_714),
    .B(n_13030),
    .Y(n_22017));
 NAND2x1_ASAP7_75t_SL g29409 (.A(n_22019),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .Y(n_22020));
 XNOR2xp5_ASAP7_75t_SL g29411 (.A(n_13025),
    .B(n_22021),
    .Y(n_22022));
 XOR2xp5_ASAP7_75t_SL g29412 (.A(n_7389),
    .B(n_7390),
    .Y(n_22021));
 OAI21x1_ASAP7_75t_SL g29414 (.A1(n_22024),
    .A2(n_22026),
    .B(n_22027),
    .Y(n_22028));
 NAND2xp5_ASAP7_75t_SL g29415 (.A(n_11201),
    .B(n_11197),
    .Y(n_22025));
 NAND3xp33_ASAP7_75t_SL g29416 (.A(n_22024),
    .B(n_11197),
    .C(n_11201),
    .Y(n_22027));
 XNOR2x1_ASAP7_75t_SL g29419 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_186),
    .Y(n_22034),
    .A(n_26146));
 MAJIxp5_ASAP7_75t_SL g29422 (.A(n_23549),
    .B(n_6179),
    .C(n_22036),
    .Y(n_22037));
 HB1xp67_ASAP7_75t_SL g29423 (.A(n_22035),
    .Y(n_22036));
 XNOR2xp5_ASAP7_75t_SL g29424 (.A(n_13476),
    .B(n_11896),
    .Y(n_22035));
 OAI21xp5_ASAP7_75t_SL g29426 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_198),
    .A2(n_22040),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_201),
    .Y(n_22041));
 NOR2xp67_ASAP7_75t_SL g29428 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_180),
    .Y(n_22040));
 XOR2x1_ASAP7_75t_SL g29429 (.A(n_22042),
    .Y(n_22043),
    .B(n_11904));
 AND2x2_ASAP7_75t_SL g29430 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_592),
    .Y(n_22042));
 XNOR2x1_ASAP7_75t_SL g29431 (.B(n_13067),
    .Y(n_22045),
    .A(n_22044));
 MAJx2_ASAP7_75t_SL g29432 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(n_21051),
    .C(n_8495),
    .Y(n_22044));
 HB1xp67_ASAP7_75t_SL g29433 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_167),
    .Y(n_22046));
 XNOR2xp5_ASAP7_75t_SL g29434 (.A(n_22049),
    .B(n_6999),
    .Y(n_22050));
 OAI22xp5_ASAP7_75t_SL g29435 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_7),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_167),
    .B1(n_22047),
    .B2(n_22048),
    .Y(n_22049));
 INVx1_ASAP7_75t_SL g29436 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_7),
    .Y(n_22047));
 INVx1_ASAP7_75t_SL g29437 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_167),
    .Y(n_22048));
 XOR2xp5_ASAP7_75t_SL g29438 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_20),
    .B(n_22051),
    .Y(n_22052));
 NAND2x1_ASAP7_75t_SL g29439 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(n_14987),
    .Y(n_22051));
 OAI22x1_ASAP7_75t_SL g29440 (.A1(n_6675),
    .A2(n_22053),
    .B1(n_20673),
    .B2(n_22054),
    .Y(n_22055));
 OAI22x1_ASAP7_75t_SL g29441 (.A1(n_22892),
    .A2(n_15001),
    .B1(n_6676),
    .B2(n_21437),
    .Y(n_22053));
 INVx1_ASAP7_75t_SL g29442 (.A(n_22053),
    .Y(n_22054));
 MAJIxp5_ASAP7_75t_SL g29443 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_71),
    .C(n_22056),
    .Y(n_22057));
 NAND2xp5_ASAP7_75t_SL g29444 (.A(n_6965),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .Y(n_22056));
 NOR2xp67_ASAP7_75t_SL g29445 (.A(n_7471),
    .B(n_26147),
    .Y(n_22061));
 XNOR2xp5_ASAP7_75t_SL g29449 (.A(n_22062),
    .B(n_22063),
    .Y(n_22064));
 INVx1_ASAP7_75t_SL g29450 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_81),
    .Y(n_22062));
 AOI22xp5_ASAP7_75t_SL g29451 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_45),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_103),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_102),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_46),
    .Y(n_22063));
 XOR2x2_ASAP7_75t_SL g29452 (.A(n_22066),
    .B(n_11972),
    .Y(n_22068));
 XOR2xp5_ASAP7_75t_SL g29453 (.A(n_26003),
    .B(n_13709),
    .Y(n_22066));
 XNOR2x1_ASAP7_75t_SL g29456 (.B(n_22072),
    .Y(n_22073),
    .A(n_22071));
 INVxp67_ASAP7_75t_SL g29459 (.A(n_22621),
    .Y(n_22072));
 XOR2xp5_ASAP7_75t_SL g29460 (.A(n_22443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_120),
    .Y(n_22076));
 XNOR2xp5_ASAP7_75t_SL g29462 (.A(n_9299),
    .B(n_22077),
    .Y(n_22078));
 XNOR2x1_ASAP7_75t_SL g29463 (.B(n_19190),
    .Y(n_22077),
    .A(n_14386));
 NOR2xp33_ASAP7_75t_SL g29464 (.A(n_13130),
    .B(n_22080),
    .Y(n_22081));
 NAND2xp5_ASAP7_75t_SL g29465 (.A(n_22295),
    .B(n_13129),
    .Y(n_22079));
 INVx1_ASAP7_75t_SL g29468 (.A(n_22083),
    .Y(n_22084));
 XNOR2xp5_ASAP7_75t_SL g29469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_104),
    .B(n_13539),
    .Y(n_22083));
 AOI21xp5_ASAP7_75t_SL g29472 (.A1(n_16559),
    .A2(n_16558),
    .B(n_17663),
    .Y(n_22087));
 XNOR2xp5_ASAP7_75t_SL g29473 (.A(n_22089),
    .B(n_14832),
    .Y(n_22090));
 OAI22xp5_ASAP7_75t_SL g29474 (.A1(n_6128),
    .A2(n_6131),
    .B1(n_23431),
    .B2(n_18858),
    .Y(n_22089));
 OAI21xp33_ASAP7_75t_SL g29475 (.A1(n_5941),
    .A2(n_5936),
    .B(n_25448),
    .Y(n_22092));
 OAI21x1_ASAP7_75t_SL g29478 (.A1(n_22094),
    .A2(n_7907),
    .B(n_22096),
    .Y(n_22097));
 NAND2xp5_ASAP7_75t_SL g29479 (.A(n_9661),
    .B(n_22093),
    .Y(n_22094));
 INVxp67_ASAP7_75t_SL g29480 (.A(n_7909),
    .Y(n_22093));
 NAND2xp5_ASAP7_75t_SL g29481 (.A(n_22095),
    .B(n_7907),
    .Y(n_22096));
 AND2x2_ASAP7_75t_SL g29482 (.A(n_9661),
    .B(n_7909),
    .Y(n_22095));
 MAJIxp5_ASAP7_75t_SL g29483 (.A(n_22100),
    .B(n_3615),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_7),
    .Y(n_22101));
 XNOR2x1_ASAP7_75t_SL g29484 (.B(n_22099),
    .Y(n_22100),
    .A(n_18826));
 XNOR2x1_ASAP7_75t_SL g29485 (.B(n_5664),
    .Y(n_22099),
    .A(n_13508));
 XNOR2xp5_ASAP7_75t_SL g29486 (.A(n_8522),
    .B(n_22103),
    .Y(n_22104));
 XNOR2xp5_ASAP7_75t_SL g29487 (.A(n_4645),
    .B(n_22290),
    .Y(n_22103));
 HB1xp67_ASAP7_75t_SL g29489 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_81),
    .Y(n_22105));
 XNOR2x1_ASAP7_75t_SL g29492 (.B(n_26026),
    .Y(n_22112),
    .A(n_22110));
 XOR2x2_ASAP7_75t_SL g29493 (.A(n_26148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_50),
    .Y(n_22110));
 INVxp67_ASAP7_75t_SL g295 (.A(n_22242),
    .Y(n_8213));
 NAND2xp5_ASAP7_75t_SL g29501 (.A(n_5780),
    .B(n_22121),
    .Y(n_11596));
 INVxp67_ASAP7_75t_SL g29502 (.A(n_22120),
    .Y(n_22121));
 MAJIxp5_ASAP7_75t_SL g29503 (.A(n_26149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_18),
    .C(n_10569),
    .Y(n_22120));
 INVx1_ASAP7_75t_SL g29506 (.A(n_26149),
    .Y(n_22123));
 OAI21x1_ASAP7_75t_SL g29513 (.A1(n_22099),
    .A2(n_21093),
    .B(n_22128),
    .Y(n_22129));
 NAND2xp5_ASAP7_75t_SL g29514 (.A(n_21092),
    .B(n_21091),
    .Y(n_22128));
 BUFx2_ASAP7_75t_SL g29521 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_283),
    .Y(n_22138));
 NOR2x1_ASAP7_75t_SL g29527 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_263),
    .B(n_22138),
    .Y(n_22142));
 OAI21xp5_ASAP7_75t_SL g29529 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_263),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_267),
    .Y(n_22143));
 OAI21xp5_ASAP7_75t_SL g29533 (.A1(n_10723),
    .A2(n_22141),
    .B(n_22153),
    .Y(n_22154));
 AOI21xp5_ASAP7_75t_SL g29534 (.A1(n_22151),
    .A2(n_22152),
    .B(n_10725),
    .Y(n_22153));
 NOR2xp67_ASAP7_75t_SL g29535 (.A(n_10721),
    .B(n_22143),
    .Y(n_22151));
 INVx1_ASAP7_75t_SL g29536 (.A(n_22142),
    .Y(n_22152));
 OAI21xp33_ASAP7_75t_SL g29537 (.A1(n_23228),
    .A2(n_22138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_281),
    .Y(n_22155));
 MAJIxp5_ASAP7_75t_SL g29538 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_76),
    .B(n_22158),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_95),
    .Y(n_22159));
 NAND2xp5_ASAP7_75t_SL g29540 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .Y(n_22157));
 NOR2xp33_ASAP7_75t_SL g29541 (.A(n_99),
    .B(n_22161),
    .Y(n_22162));
 AND3x2_ASAP7_75t_SL g29545 (.A(n_17869),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .C(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[6]),
    .Y(n_22164));
 AO21x2_ASAP7_75t_SL g29547 (.A1(n_26028),
    .A2(n_4787),
    .B(n_22166),
    .Y(n_22167));
 OAI21xp5_ASAP7_75t_SL g29549 (.A1(n_26028),
    .A2(n_4787),
    .B(n_22164),
    .Y(n_22166));
 NOR2xp33_ASAP7_75t_SL g29550 (.A(n_22167),
    .B(n_11289),
    .Y(n_22169));
 NAND2xp5_ASAP7_75t_SL g29551 (.A(n_22167),
    .B(n_11289),
    .Y(n_22170));
 MAJIxp5_ASAP7_75t_SL g29552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_97),
    .B(n_22171),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_105),
    .Y(n_22172));
 NAND2xp5_ASAP7_75t_SL g29553 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .Y(n_22171));
 OAI22xp5_ASAP7_75t_SL g29554 (.A1(n_22171),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_97),
    .B1(n_22173),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_96),
    .Y(n_22174));
 INVx1_ASAP7_75t_SL g29555 (.A(n_22171),
    .Y(n_22173));
 XNOR2x1_ASAP7_75t_SL g29556 (.B(n_22177),
    .Y(n_22178),
    .A(n_8702));
 XNOR2xp5_ASAP7_75t_SL g29557 (.A(n_22176),
    .B(n_22175),
    .Y(n_22177));
 NAND2x1_ASAP7_75t_SL g29558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_778),
    .B(n_2173),
    .Y(n_22175));
 AND2x2_ASAP7_75t_SL g29559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_554),
    .B(n_2163),
    .Y(n_22176));
 MAJIxp5_ASAP7_75t_SL g29560 (.A(n_8702),
    .B(n_22179),
    .C(n_22176),
    .Y(n_22180));
 INVx1_ASAP7_75t_SL g29561 (.A(n_22175),
    .Y(n_22179));
 MAJIxp5_ASAP7_75t_SL g29562 (.A(n_18776),
    .B(n_22182),
    .C(n_22187),
    .Y(n_22188));
 INVxp67_ASAP7_75t_SL g29563 (.A(n_26247),
    .Y(n_22182));
 INVxp67_ASAP7_75t_SL g29565 (.A(n_22186),
    .Y(n_22187));
 XNOR2x1_ASAP7_75t_SL g29566 (.B(n_22185),
    .Y(n_22186),
    .A(n_22183));
 NAND2x1_ASAP7_75t_SL g29567 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(n_9154),
    .Y(n_22183));
 AOI22xp5_ASAP7_75t_SL g29568 (.A1(n_13766),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_45),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_64),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_46),
    .Y(n_22185));
 MAJIxp5_ASAP7_75t_SL g29571 (.A(n_13766),
    .B(n_22183),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_46),
    .Y(n_22190));
 XOR2xp5_ASAP7_75t_SL g29595 (.A(n_22215),
    .B(n_22220),
    .Y(n_22221));
 MAJx2_ASAP7_75t_SL g29596 (.A(n_8322),
    .B(n_22214),
    .C(n_8329),
    .Y(n_22215));
 AOI22xp5_ASAP7_75t_SL g29598 (.A1(n_22217),
    .A2(n_22219),
    .B1(n_22216),
    .B2(n_22218),
    .Y(n_22220));
 INVx1_ASAP7_75t_SL g29599 (.A(n_22216),
    .Y(n_22217));
 NAND2xp5_ASAP7_75t_SL g296 (.A(n_13770),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_67),
    .Y(n_24678));
 XNOR2x1_ASAP7_75t_SL g29600 (.B(n_21242),
    .Y(n_22216),
    .A(n_8312));
 INVx1_ASAP7_75t_SL g29601 (.A(n_22218),
    .Y(n_22219));
 MAJx2_ASAP7_75t_SL g29602 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_25),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_93),
    .Y(n_22218));
 MAJIxp5_ASAP7_75t_SL g29603 (.A(n_8322),
    .B(n_22214),
    .C(n_8329),
    .Y(n_22222));
 XNOR2x1_ASAP7_75t_SL g29605 (.B(n_22231),
    .Y(n_22232),
    .A(n_22224));
 XNOR2x1_ASAP7_75t_SL g29606 (.B(n_6304),
    .Y(n_22224),
    .A(n_13578));
 XNOR2xp5_ASAP7_75t_SL g29608 (.A(n_26151),
    .B(n_22229),
    .Y(n_22230));
 MAJIxp5_ASAP7_75t_SL g29611 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_37),
    .C(n_6145),
    .Y(n_22229));
 XNOR2xp5_ASAP7_75t_SL g29613 (.A(n_22234),
    .B(n_22241),
    .Y(n_22242));
 MAJIxp5_ASAP7_75t_SL g29614 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_46),
    .B(n_22883),
    .C(n_20512),
    .Y(n_22234));
 XNOR2xp5_ASAP7_75t_SL g29615 (.A(n_22236),
    .B(n_26152),
    .Y(n_22241));
 INVx1_ASAP7_75t_SL g29616 (.A(n_22235),
    .Y(n_22236));
 OR2x2_ASAP7_75t_SL g29617 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_100),
    .Y(n_22235));
 XNOR2xp5_ASAP7_75t_SL g29622 (.A(n_22243),
    .B(n_22246),
    .Y(n_22247));
 MAJIxp5_ASAP7_75t_SL g29623 (.A(n_22017),
    .B(n_13417),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_779),
    .Y(n_22243));
 XOR2xp5_ASAP7_75t_SL g29624 (.A(n_22244),
    .B(n_22245),
    .Y(n_22246));
 NAND2xp5_ASAP7_75t_SL g29625 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_616),
    .B(n_2179),
    .Y(n_22244));
 NAND2x1_ASAP7_75t_SL g29626 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_648),
    .B(n_2169),
    .Y(n_22245));
 INVxp67_ASAP7_75t_SL g29627 (.A(n_22245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_74));
 XNOR2xp5_ASAP7_75t_SL g29629 (.A(n_22250),
    .B(n_22251),
    .Y(n_22252));
 NAND2x1_ASAP7_75t_SL g29630 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .Y(n_22250));
 NAND2x1_ASAP7_75t_SL g29631 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .B(n_13231),
    .Y(n_22251));
 XNOR2xp5_ASAP7_75t_SL g29632 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_148),
    .B(n_11357),
    .Y(n_11121));
 MAJIxp5_ASAP7_75t_SL g29633 (.A(n_22256),
    .B(n_22257),
    .C(n_22259),
    .Y(n_22260));
 OAI21x1_ASAP7_75t_SL g29654 (.A1(n_22287),
    .A2(n_20681),
    .B(n_26239),
    .Y(n_22290));
 MAJx2_ASAP7_75t_SL g29657 (.A(n_22294),
    .B(n_7284),
    .C(n_19442),
    .Y(n_22295));
 XNOR2x1_ASAP7_75t_SL g29658 (.B(n_22293),
    .Y(n_22294),
    .A(n_22292));
 XNOR2xp5_ASAP7_75t_SL g29659 (.A(n_22291),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_183),
    .Y(n_22292));
 INVx1_ASAP7_75t_SL g29660 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_21),
    .Y(n_22291));
 INVx2_ASAP7_75t_SL g29661 (.A(n_10356),
    .Y(n_22293));
 XNOR2xp5_ASAP7_75t_SL g29662 (.A(n_18881),
    .B(n_22294),
    .Y(n_22296));
 AO21x1_ASAP7_75t_SL g29670 (.A1(n_26029),
    .A2(n_22309),
    .B(n_22311),
    .Y(n_22312));
 INVx2_ASAP7_75t_SL g29673 (.A(n_22306),
    .Y(n_22307));
 OA21x2_ASAP7_75t_SL g29674 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_304),
    .A2(n_12562),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_305),
    .Y(n_22306));
 INVx1_ASAP7_75t_SL g29675 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270),
    .Y(n_22308));
 O2A1O1Ixp33_ASAP7_75t_SRAM g29676 (.A1(n_14176),
    .A2(n_22306),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270),
    .C(n_26030),
    .Y(n_22311));
 OAI21xp33_ASAP7_75t_SL g29678 (.A1(n_22306),
    .A2(n_26031),
    .B(n_22314),
    .Y(n_22315));
 NAND2xp5_ASAP7_75t_SL g29679 (.A(n_22306),
    .B(n_26031),
    .Y(n_22314));
 XNOR2x1_ASAP7_75t_SL g29681 (.B(n_22317),
    .Y(n_22318),
    .A(n_22084));
 XNOR2x1_ASAP7_75t_SL g29682 (.B(n_22316),
    .Y(n_22317),
    .A(n_9966));
 XNOR2x1_ASAP7_75t_SL g29683 (.B(n_12787),
    .Y(n_22316),
    .A(n_7121));
 MAJIxp5_ASAP7_75t_SL g29684 (.A(n_22083),
    .B(n_9966),
    .C(n_22319),
    .Y(n_22320));
 INVx1_ASAP7_75t_SL g29685 (.A(n_22316),
    .Y(n_22319));
 AO21x2_ASAP7_75t_SL g29686 (.A1(n_24169),
    .A2(n_24029),
    .B(n_24028),
    .Y(n_22323));
 OR2x2_ASAP7_75t_SL g29688 (.A(n_21357),
    .B(n_21948),
    .Y(n_22321));
 NAND2xp5_ASAP7_75t_SL g29689 (.A(n_24021),
    .B(n_22325),
    .Y(n_22326));
 INVx1_ASAP7_75t_SL g29690 (.A(n_22324),
    .Y(n_22325));
 INVxp67_ASAP7_75t_SL g29691 (.A(n_22321),
    .Y(n_22324));
 NAND2xp5_ASAP7_75t_SL g29696 (.A(n_22331),
    .B(n_10657),
    .Y(n_22332));
 INVxp67_ASAP7_75t_SRAM g29697 (.A(n_23367),
    .Y(n_22331));
 OAI21xp5_ASAP7_75t_SL g29698 (.A1(n_22333),
    .A2(n_21527),
    .B(n_10657),
    .Y(n_22334));
 INVxp67_ASAP7_75t_SL g29699 (.A(n_22331),
    .Y(n_22333));
 NAND2xp5_ASAP7_75t_SL g29700 (.A(n_23366),
    .B(n_21841),
    .Y(n_22335));
 AO21x1_ASAP7_75t_SL g29745 (.A1(n_23820),
    .A2(n_21875),
    .B(n_21876),
    .Y(n_22379));
 XNOR2x1_ASAP7_75t_SL g29774 (.B(n_22418),
    .Y(n_22419),
    .A(n_22417));
 AOI22x1_ASAP7_75t_SL g29775 (.A1(n_22414),
    .A2(n_22416),
    .B1(n_22413),
    .B2(n_15003),
    .Y(n_22417));
 INVx2_ASAP7_75t_SL g29776 (.A(n_22413),
    .Y(n_22414));
 XNOR2x1_ASAP7_75t_SL g29777 (.B(n_22412),
    .Y(n_22413),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_132));
 INVxp67_ASAP7_75t_SL g29778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_47),
    .Y(n_22412));
 HB1xp67_ASAP7_75t_SL g29780 (.A(n_22521),
    .Y(n_22418));
 OAI21xp5_ASAP7_75t_SL g29782 (.A1(n_22426),
    .A2(n_4430),
    .B(n_13142),
    .Y(n_22427));
 OAI31xp33_ASAP7_75t_SL g29783 (.A1(n_13138),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_119),
    .A3(n_22422),
    .B(n_22425),
    .Y(n_22426));
 AO22x2_ASAP7_75t_SL g29784 (.A1(n_22420),
    .A2(n_22421),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_57),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_53),
    .Y(n_22422));
 INVx1_ASAP7_75t_SL g29785 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_53),
    .Y(n_22420));
 INVx1_ASAP7_75t_SL g29786 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_57),
    .Y(n_22421));
 NAND3xp33_ASAP7_75t_SL g29787 (.A(n_22423),
    .B(n_22424),
    .C(n_22422),
    .Y(n_22425));
 INVxp67_ASAP7_75t_SL g29789 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_119),
    .Y(n_22424));
 AOI21xp5_ASAP7_75t_SL g29790 (.A1(n_22430),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_310),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_313),
    .Y(n_22431));
 AND2x2_ASAP7_75t_SL g29791 (.A(n_9695),
    .B(n_22429),
    .Y(n_22430));
 OAI21x1_ASAP7_75t_SL g29792 (.A1(n_14941),
    .A2(n_11124),
    .B(n_10445),
    .Y(n_22429));
 AOI21x1_ASAP7_75t_SL g29796 (.A1(n_22436),
    .A2(n_5880),
    .B(n_5881),
    .Y(n_22437));
 OR2x2_ASAP7_75t_SL g29797 (.A(n_22435),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_204),
    .Y(n_22436));
 AO21x1_ASAP7_75t_SL g29798 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_268),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_270),
    .Y(n_22435));
 AOI21x1_ASAP7_75t_SL g29799 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_445),
    .A2(n_22439),
    .B(n_4087),
    .Y(n_22440));
 NOR2xp33_ASAP7_75t_SL g298 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_135),
    .Y(n_6528));
 AO21x2_ASAP7_75t_SL g29800 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .A2(n_22438),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_478),
    .Y(n_22439));
 NOR2xp33_ASAP7_75t_SL g29801 (.A(n_22611),
    .B(n_21126),
    .Y(n_22438));
 XNOR2xp5_ASAP7_75t_SL g29802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_713),
    .B(n_22442),
    .Y(n_22443));
 XOR2xp5_ASAP7_75t_SL g29803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_553),
    .B(n_22441),
    .Y(n_22442));
 AND2x2_ASAP7_75t_SL g29804 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_776),
    .B(n_2158),
    .Y(n_22441));
 XNOR2xp5_ASAP7_75t_SL g29808 (.A(n_22448),
    .B(n_26241),
    .Y(n_22451));
 INVx1_ASAP7_75t_SL g29809 (.A(n_8185),
    .Y(n_22448));
 AOI22xp5_ASAP7_75t_SL g29813 (.A1(n_22457),
    .A2(n_20731),
    .B1(n_21359),
    .B2(n_10309),
    .Y(n_22458));
 NAND2xp5_ASAP7_75t_SL g29814 (.A(n_22456),
    .B(n_21322),
    .Y(n_22457));
 XNOR2xp5_ASAP7_75t_SL g29815 (.A(n_20022),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_377),
    .Y(n_22456));
 XNOR2x1_ASAP7_75t_SL g29816 (.B(n_22462),
    .Y(n_22463),
    .A(n_21415));
 XNOR2x1_ASAP7_75t_SL g29817 (.B(n_22461),
    .Y(n_22462),
    .A(n_22459));
 MAJx2_ASAP7_75t_SL g29818 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_113),
    .C(n_15585),
    .Y(n_22459));
 BUFx2_ASAP7_75t_SL g29819 (.A(n_22460),
    .Y(n_22461));
 NAND2xp5_ASAP7_75t_SL g29820 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_23),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_83),
    .Y(n_22460));
 MAJIxp5_ASAP7_75t_SL g29821 (.A(n_21415),
    .B(n_22461),
    .C(n_22464),
    .Y(n_22465));
 INVxp67_ASAP7_75t_SL g29822 (.A(n_22459),
    .Y(n_22464));
 OAI22xp5_ASAP7_75t_SL g29834 (.A1(n_22478),
    .A2(n_13186),
    .B1(n_19882),
    .B2(n_22479),
    .Y(n_22480));
 MAJIxp5_ASAP7_75t_SL g29835 (.A(n_22477),
    .B(n_13387),
    .C(n_13502),
    .Y(n_22478));
 XOR2x2_ASAP7_75t_SL g29836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_126),
    .Y(n_22477));
 INVx1_ASAP7_75t_SL g29837 (.A(n_22478),
    .Y(n_22479));
 MAJIxp5_ASAP7_75t_SL g29838 (.A(n_22221),
    .B(n_13185),
    .C(n_22481),
    .Y(n_22482));
 HB1xp67_ASAP7_75t_SL g29839 (.A(n_22479),
    .Y(n_22481));
 NOR2xp67_ASAP7_75t_SL g29842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_258),
    .B(n_22486),
    .Y(n_22487));
 XNOR2xp5_ASAP7_75t_SL g29843 (.A(n_18838),
    .B(n_22485),
    .Y(n_22486));
 XNOR2xp5_ASAP7_75t_SL g29844 (.A(n_5570),
    .B(n_26083),
    .Y(n_22485));
 NAND2xp5_ASAP7_75t_SL g29845 (.A(n_22486),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_258),
    .Y(n_22488));
 AOI21xp5_ASAP7_75t_SL g29846 (.A1(n_22485),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_243),
    .Y(n_22489));
 OR2x2_ASAP7_75t_SL g29847 (.A(n_22495),
    .B(n_21968),
    .Y(n_22496));
 INVx1_ASAP7_75t_SL g29848 (.A(n_22494),
    .Y(n_22495));
 XNOR2xp5_ASAP7_75t_SL g29849 (.A(n_22490),
    .B(n_26159),
    .Y(n_22494));
 INVx1_ASAP7_75t_SL g29850 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_197),
    .Y(n_22490));
 NAND2xp5_ASAP7_75t_SL g29854 (.A(n_22495),
    .B(n_21968),
    .Y(n_22497));
 INVx1_ASAP7_75t_SL g29855 (.A(n_22496),
    .Y(n_22498));
 OAI22x1_ASAP7_75t_SL g29857 (.A1(n_22499),
    .A2(n_20588),
    .B1(n_20589),
    .B2(n_15549),
    .Y(n_22500));
 AND2x2_ASAP7_75t_SL g29858 (.A(n_19970),
    .B(n_24102),
    .Y(n_22499));
 NAND2xp33_ASAP7_75t_SL g29860 (.A(n_22506),
    .B(n_22510),
    .Y(n_22511));
 OAI221xp5_ASAP7_75t_SL g29861 (.A1(n_11502),
    .A2(n_22503),
    .B1(n_22504),
    .B2(n_11501),
    .C(n_20221),
    .Y(n_22506));
 XNOR2x1_ASAP7_75t_SL g29862 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_147),
    .Y(n_22503),
    .A(n_11509));
 INVxp67_ASAP7_75t_SL g29863 (.A(n_22503),
    .Y(n_22504));
 INVx1_ASAP7_75t_SL g29865 (.A(n_22509),
    .Y(n_22510));
 O2A1O1Ixp33_ASAP7_75t_SL g29866 (.A1(n_11502),
    .A2(n_22503),
    .B(n_22508),
    .C(n_20221),
    .Y(n_22509));
 NAND2xp5_ASAP7_75t_SL g29867 (.A(n_11502),
    .B(n_22503),
    .Y(n_22508));
 AO21x2_ASAP7_75t_SL g29869 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_250),
    .A2(n_22506),
    .B(n_22509),
    .Y(n_22512));
 XNOR2x1_ASAP7_75t_SL g29871 (.B(n_22518),
    .Y(n_22519),
    .A(n_22517));
 OAI21xp5_ASAP7_75t_SL g29872 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_144),
    .A2(n_22514),
    .B(n_22516),
    .Y(n_22517));
 OA21x2_ASAP7_75t_SL g29873 (.A1(n_13771),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109),
    .Y(n_22514));
 NAND2xp5_ASAP7_75t_SL g29874 (.A(n_22514),
    .B(n_22515),
    .Y(n_22516));
 INVxp67_ASAP7_75t_SL g29875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_143),
    .Y(n_22515));
 INVx1_ASAP7_75t_SL g29876 (.A(n_11783),
    .Y(n_22518));
 MAJIxp5_ASAP7_75t_SL g29877 (.A(n_22520),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_149),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_144),
    .Y(n_22521));
 INVx1_ASAP7_75t_SL g29878 (.A(n_22514),
    .Y(n_22520));
 AO22x2_ASAP7_75t_SL g29879 (.A1(n_22523),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_80),
    .B1(n_22522),
    .B2(n_8895),
    .Y(n_22524));
 INVxp67_ASAP7_75t_SL g29880 (.A(n_22522),
    .Y(n_22523));
 NAND2x1_ASAP7_75t_SL g29881 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(n_22522));
 NOR2xp67_ASAP7_75t_SL g29882 (.A(n_22522),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_80),
    .Y(n_22525));
 XNOR2x1_ASAP7_75t_SL g29890 (.B(n_15233),
    .Y(n_22540),
    .A(n_22539));
 XOR2xp5_ASAP7_75t_SL g29891 (.A(n_22537),
    .B(n_22538),
    .Y(n_22539));
 XNOR2x1_ASAP7_75t_SL g29892 (.B(n_22536),
    .Y(n_22537),
    .A(n_22533));
 XNOR2x1_ASAP7_75t_SL g29893 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_643),
    .Y(n_22533),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_739));
 AOI21x1_ASAP7_75t_SL g29894 (.A1(n_22534),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_n_709),
    .B(n_22535),
    .Y(n_22536));
 OR2x2_ASAP7_75t_SL g29895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_549),
    .B(n_21377),
    .Y(n_22534));
 AND2x2_ASAP7_75t_SL g29896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_549),
    .B(n_21377),
    .Y(n_22535));
 MAJIxp5_ASAP7_75t_SL g29897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_156),
    .B(n_19658),
    .C(n_22606),
    .Y(n_22538));
 MAJx2_ASAP7_75t_SL g29898 (.A(n_9671),
    .B(n_22537),
    .C(n_22538),
    .Y(n_22541));
 NAND2xp33_ASAP7_75t_L g299 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_135),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121),
    .Y(n_6527));
 NAND2xp5_ASAP7_75t_SL g29900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_643),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_739),
    .Y(n_22542));
 NOR2xp33_ASAP7_75t_SL g29901 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_739),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_643),
    .Y(n_22543));
 NAND2xp33_ASAP7_75t_SL g29914 (.A(n_22564),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_248),
    .Y(n_22565));
 NAND2xp5_ASAP7_75t_SL g29915 (.A(n_22561),
    .B(n_23086),
    .Y(n_22564));
 XNOR2xp5_ASAP7_75t_SL g29916 (.A(n_22557),
    .B(n_22560),
    .Y(n_22561));
 XNOR2x1_ASAP7_75t_SL g29917 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_6),
    .Y(n_22557),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_119));
 AOI22xp5_ASAP7_75t_SL g29918 (.A1(n_22558),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_154),
    .B1(n_22559),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_177),
    .Y(n_22560));
 INVx1_ASAP7_75t_SL g29919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_177),
    .Y(n_22558));
 INVx1_ASAP7_75t_SL g29920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_154),
    .Y(n_22559));
 HB1xp67_ASAP7_75t_SL g29922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_135),
    .Y(n_22562));
 OAI21xp5_ASAP7_75t_SL g29923 (.A1(n_22566),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_31),
    .B(n_22564),
    .Y(n_22567));
 NOR2xp67_ASAP7_75t_SL g29924 (.A(n_23086),
    .B(n_22561),
    .Y(n_22566));
 MAJIxp5_ASAP7_75t_SL g29925 (.A(n_2877),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_154),
    .C(n_22557),
    .Y(n_22568));
 XNOR2xp5_ASAP7_75t_SL g29955 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .B(n_12288),
    .Y(n_22608));
 MAJIxp5_ASAP7_75t_SL g29956 (.A(n_10417),
    .B(n_22975),
    .C(n_21404),
    .Y(n_22609));
 NAND2xp5_ASAP7_75t_SL g29957 (.A(n_22610),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_62),
    .Y(n_22611));
 NAND2xp5_ASAP7_75t_SL g29973 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(n_22616),
    .Y(n_22626));
 HB1xp67_ASAP7_75t_SRAM g29985 (.A(n_22616),
    .Y(n_22637));
 XOR2xp5_ASAP7_75t_SL g3 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_17),
    .Y(n_21803));
 OAI31xp33_ASAP7_75t_SL g30 (.A1(n_7514),
    .A2(n_7516),
    .A3(n_19193),
    .B(n_19013),
    .Y(n_24711));
 INVxp67_ASAP7_75t_SL g300 (.A(n_6523),
    .Y(n_6524));
 AND2x2_ASAP7_75t_SL g30061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_584),
    .B(n_12748),
    .Y(n_22713));
 MAJIxp5_ASAP7_75t_SL g30063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .B(n_22715),
    .C(n_21920),
    .Y(n_22716));
 MAJIxp5_ASAP7_75t_L g30064 (.A(n_22712),
    .B(n_22713),
    .C(n_22714),
    .Y(n_22715));
 OAI22xp5_ASAP7_75t_SL g30068 (.A1(n_22721),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_129),
    .B1(n_26032),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .Y(n_22724));
 MAJx2_ASAP7_75t_SL g30072 (.A(n_7316),
    .B(n_7315),
    .C(n_7313),
    .Y(n_22726));
 XNOR2x1_ASAP7_75t_SL g30073 (.B(n_9849),
    .Y(n_22727),
    .A(n_9848));
 XNOR2xp5_ASAP7_75t_SL g30077 (.A(n_21583),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_92),
    .Y(n_22732));
 XNOR2xp5_ASAP7_75t_L g30079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_187),
    .Y(n_22734));
 XOR2xp5_ASAP7_75t_SL g30081 (.A(n_10078),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_209),
    .Y(n_22736));
 XNOR2xp5_ASAP7_75t_SL g30084 (.A(n_22739),
    .B(n_22740),
    .Y(n_22741));
 NAND2x1_ASAP7_75t_SL g30085 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .Y(n_22739));
 NAND2xp5_ASAP7_75t_SL g30086 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(n_22740));
 NAND2xp5_ASAP7_75t_SL g30087 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .B(n_22743),
    .Y(n_22744));
 XNOR2xp5_ASAP7_75t_SL g30091 (.A(n_18665),
    .B(n_26243),
    .Y(n_22779));
 NAND2xp5_ASAP7_75t_SL g30096 (.A(n_22780),
    .B(n_22785),
    .Y(n_22786));
 XNOR2xp5_ASAP7_75t_SL g30097 (.A(n_15939),
    .B(n_8615),
    .Y(n_22780));
 AO21x1_ASAP7_75t_SL g30098 (.A1(n_22783),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_340),
    .B(n_22784),
    .Y(n_22785));
 NAND2xp5_ASAP7_75t_SL g30099 (.A(n_22781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_256),
    .Y(n_22783));
 NAND2xp5_ASAP7_75t_SL g301 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(n_3190),
    .Y(n_6523));
 INVx1_ASAP7_75t_SL g30100 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_309),
    .Y(n_22781));
 NOR2xp33_ASAP7_75t_SL g30102 (.A(n_22781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_256),
    .Y(n_22784));
 NAND2x1_ASAP7_75t_SL g30103 (.A(n_26244),
    .B(n_22793),
    .Y(n_22794));
 NAND2xp5_ASAP7_75t_SL g30104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_263),
    .Y(n_22787));
 NOR2xp33_ASAP7_75t_SL g30105 (.A(n_22787),
    .B(n_13629),
    .Y(n_22790));
 INVxp67_ASAP7_75t_SL g30106 (.A(n_15561),
    .Y(n_22791));
 OAI21xp5_ASAP7_75t_SL g30107 (.A1(n_9866),
    .A2(n_22787),
    .B(n_2169),
    .Y(n_22792));
 A2O1A1O1Ixp25_ASAP7_75t_SL g30108 (.A1(n_22795),
    .A2(n_22797),
    .B(n_22798),
    .C(n_22799),
    .D(n_22801),
    .Y(n_22802));
 NOR2xp33_ASAP7_75t_SL g30109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_257),
    .B(n_9481),
    .Y(n_22795));
 INVx2_ASAP7_75t_SL g30110 (.A(n_22796),
    .Y(n_22797));
 OA21x2_ASAP7_75t_SL g30111 (.A1(n_21508),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_305),
    .Y(n_22796));
 OAI21xp5_ASAP7_75t_SL g30112 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_257),
    .A2(n_9483),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_260),
    .Y(n_22798));
 NAND2xp5_ASAP7_75t_SL g30113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_70),
    .Y(n_22799));
 NAND2xp5_ASAP7_75t_SL g30114 (.A(n_2165),
    .B(n_22800),
    .Y(n_22801));
 OR2x2_ASAP7_75t_SL g30115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_193),
    .Y(n_22800));
 OAI21xp5_ASAP7_75t_SL g30116 (.A1(n_22803),
    .A2(n_22796),
    .B(n_22804),
    .Y(n_22805));
 INVxp67_ASAP7_75t_SL g30117 (.A(n_22795),
    .Y(n_22803));
 INVx1_ASAP7_75t_SL g30118 (.A(n_22798),
    .Y(n_22804));
 OAI21x1_ASAP7_75t_SL g30119 (.A1(n_9481),
    .A2(n_22796),
    .B(n_9483),
    .Y(n_22807));
 XOR2xp5_ASAP7_75t_SL g30120 (.A(n_9700),
    .B(n_22814),
    .Y(n_22815));
 XOR2x2_ASAP7_75t_SL g30121 (.A(n_9704),
    .B(n_22813),
    .Y(n_22814));
 AOI21x1_ASAP7_75t_SL g30122 (.A1(n_26164),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_118),
    .B(n_22812),
    .Y(n_22813));
 AND2x2_ASAP7_75t_SL g30126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_75),
    .Y(n_22812));
 XNOR2xp5_ASAP7_75t_SL g30127 (.A(n_8069),
    .B(n_22818),
    .Y(n_22819));
 OAI22xp5_ASAP7_75t_SL g30128 (.A1(n_22816),
    .A2(n_22814),
    .B1(n_9700),
    .B2(n_22817),
    .Y(n_22818));
 INVx1_ASAP7_75t_SL g30129 (.A(n_9700),
    .Y(n_22816));
 INVx1_ASAP7_75t_SL g30130 (.A(n_22814),
    .Y(n_22817));
 MAJIxp5_ASAP7_75t_SL g30131 (.A(n_22815),
    .B(n_8072),
    .C(n_8071),
    .Y(n_22820));
 OAI21x1_ASAP7_75t_SL g30132 (.A1(n_22816),
    .A2(n_22822),
    .B(n_22824),
    .Y(n_22825));
 NOR2xp33_ASAP7_75t_SL g30133 (.A(n_22821),
    .B(n_9704),
    .Y(n_22822));
 INVxp67_ASAP7_75t_SL g30134 (.A(n_22813),
    .Y(n_22821));
 NAND2xp5_ASAP7_75t_SL g30135 (.A(n_22823),
    .B(n_9704),
    .Y(n_22824));
 INVxp67_ASAP7_75t_SL g30136 (.A(n_22813),
    .Y(n_22823));
 XOR2xp5_ASAP7_75t_SL g30154 (.A(n_9708),
    .B(n_9709),
    .Y(n_22842));
 HB1xp67_ASAP7_75t_SRAM g30156 (.A(n_22843),
    .Y(n_22845));
 XNOR2xp5_ASAP7_75t_SL g30158 (.A(n_6062),
    .B(n_10842),
    .Y(n_22848));
 MAJIxp5_ASAP7_75t_SL g30159 (.A(n_9237),
    .B(n_2566),
    .C(n_11892),
    .Y(n_22849));
 OR2x2_ASAP7_75t_SL g30161 (.A(n_22848),
    .B(n_22849),
    .Y(n_22850));
 NAND2xp5_ASAP7_75t_SL g30162 (.A(n_18605),
    .B(n_22852),
    .Y(n_22853));
 HB1xp67_ASAP7_75t_SRAM g30163 (.A(n_22850),
    .Y(n_22852));
 XNOR2x1_ASAP7_75t_SL g30164 (.B(n_20814),
    .Y(n_22854),
    .A(n_20809));
 MAJIxp5_ASAP7_75t_SL g30166 (.A(n_19323),
    .B(n_19325),
    .C(n_19327),
    .Y(n_22856));
 HB1xp67_ASAP7_75t_SRAM g30168 (.A(n_22859),
    .Y(n_22860));
 AOI221xp5_ASAP7_75t_SL g30169 (.A1(n_22854),
    .A2(n_23408),
    .B1(n_12114),
    .B2(n_22858),
    .C(n_22856),
    .Y(n_22859));
 INVxp67_ASAP7_75t_SL g30171 (.A(n_22854),
    .Y(n_22858));
 OAI21xp5_ASAP7_75t_SL g30172 (.A1(n_22859),
    .A2(n_19594),
    .B(n_19595),
    .Y(n_22862));
 NAND2xp5_ASAP7_75t_SL g30173 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .B(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[6]),
    .Y(n_22863));
 INVxp67_ASAP7_75t_SL g30175 (.A(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[50]),
    .Y(n_22864));
 AND2x2_ASAP7_75t_SL g30183 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22873));
 NAND2x1_ASAP7_75t_SL g30186 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .Y(n_22876));
 INVxp33_ASAP7_75t_L g30190 (.A(n_22879),
    .Y(n_22880));
 OAI21xp5_ASAP7_75t_SL g30198 (.A1(n_22889),
    .A2(n_21664),
    .B(n_22891),
    .Y(n_22892));
 INVx2_ASAP7_75t_SL g30199 (.A(n_22888),
    .Y(n_22889));
 INVx1_ASAP7_75t_SL g302 (.A(n_20883),
    .Y(n_20885));
 MAJx2_ASAP7_75t_SL g30200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_71),
    .B(n_20831),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_70),
    .Y(n_22888));
 NAND2xp5_ASAP7_75t_SL g30201 (.A(n_21664),
    .B(n_22890),
    .Y(n_22891));
 INVx2_ASAP7_75t_L g30202 (.A(n_22888),
    .Y(n_22890));
 XOR2xp5_ASAP7_75t_SL g30203 (.A(n_22889),
    .B(n_11830),
    .Y(n_22893));
 MAJx2_ASAP7_75t_SL g30206 (.A(n_21673),
    .B(n_22890),
    .C(n_4367),
    .Y(n_22896));
 XOR2xp5_ASAP7_75t_SL g30258 (.A(n_22242),
    .B(n_11469),
    .Y(n_22948));
 XOR2xp5_ASAP7_75t_SL g30260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_218),
    .B(n_20195),
    .Y(n_22950));
 INVx1_ASAP7_75t_SL g30261 (.A(n_20195),
    .Y(n_22951));
 AND2x2_ASAP7_75t_SL g30263 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .Y(n_22953));
 NAND2xp5_ASAP7_75t_SL g30264 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .Y(n_22954));
 OA21x2_ASAP7_75t_SL g30265 (.A1(n_6223),
    .A2(n_6220),
    .B(n_6225),
    .Y(n_22955));
 OAI21xp5_ASAP7_75t_SL g30266 (.A1(n_6223),
    .A2(n_6220),
    .B(n_6225),
    .Y(n_22956));
 XOR2x2_ASAP7_75t_SL g30268 (.A(n_9076),
    .B(n_18968),
    .Y(n_22958));
 OA31x2_ASAP7_75t_SL g30269 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_286),
    .A2(n_13635),
    .A3(n_15561),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_295),
    .Y(n_22959));
 OAI31xp67_ASAP7_75t_SL g30270 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_286),
    .A2(n_13635),
    .A3(n_15561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_295),
    .Y(n_22960));
 NAND2xp5_ASAP7_75t_SL g30273 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .Y(n_22962));
 XOR2xp5_ASAP7_75t_SL g30276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_234),
    .B(n_22966),
    .Y(n_22967));
 XNOR2xp5_ASAP7_75t_SL g30277 (.A(n_7195),
    .B(n_7200),
    .Y(n_22966));
 OAI21xp5_ASAP7_75t_SL g30278 (.A1(n_22968),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_286),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_295),
    .Y(n_22969));
 AOI21xp5_ASAP7_75t_SL g30279 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_310),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_308),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_311),
    .Y(n_22968));
 OAI21xp33_ASAP7_75t_SL g30280 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .A2(n_6382),
    .B(n_22970),
    .Y(n_22971));
 AOI21xp33_ASAP7_75t_SL g30281 (.A1(n_6384),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_500),
    .B(n_6385),
    .Y(n_22970));
 MAJIxp5_ASAP7_75t_SL g30282 (.A(n_22972),
    .B(n_17398),
    .C(n_17404),
    .Y(n_22973));
 MAJIxp5_ASAP7_75t_SL g30283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_227),
    .Y(n_22972));
 OAI22xp5_ASAP7_75t_SL g30285 (.A1(n_22318),
    .A2(n_22975),
    .B1(n_22976),
    .B2(n_21407),
    .Y(n_22977));
 MAJx2_ASAP7_75t_SL g30286 (.A(n_13476),
    .B(n_15334),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_243),
    .Y(n_22975));
 INVx1_ASAP7_75t_SL g30287 (.A(n_22975),
    .Y(n_22976));
 HB1xp67_ASAP7_75t_SL g30288 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_129),
    .Y(n_22978));
 OA21x2_ASAP7_75t_SL g30290 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_123),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_142),
    .B(n_22979),
    .Y(n_22980));
 INVxp67_ASAP7_75t_SL g30291 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_129),
    .Y(n_22979));
 AOI21xp5_ASAP7_75t_SL g30294 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_298),
    .A2(n_19969),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_301),
    .Y(n_22983));
 XNOR2xp5_ASAP7_75t_SL g30297 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_194),
    .B(n_22988),
    .Y(n_22989));
 XNOR2xp5_ASAP7_75t_SL g30298 (.A(n_22987),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_125),
    .Y(n_22988));
 INVx1_ASAP7_75t_SL g30299 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_81),
    .Y(n_22987));
 INVx1_ASAP7_75t_SL g303 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_181),
    .Y(n_6519));
 XOR2xp5_ASAP7_75t_SL g30303 (.A(n_18933),
    .B(n_6298),
    .Y(n_22994));
 MAJIxp5_ASAP7_75t_SL g30304 (.A(n_20372),
    .B(n_11800),
    .C(n_4957),
    .Y(n_6298));
 XNOR2x1_ASAP7_75t_SL g30308 (.B(n_6524),
    .Y(n_23000),
    .A(n_26063));
 XNOR2xp5_ASAP7_75t_SL g30311 (.A(n_12584),
    .B(n_23001),
    .Y(n_23002));
 AOI22xp5_ASAP7_75t_SL g30312 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_42),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_69),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_68),
    .B2(n_22878),
    .Y(n_23001));
 XNOR2x1_ASAP7_75t_SL g30318 (.B(n_23014),
    .Y(n_23015),
    .A(n_23445));
 AOI21x1_ASAP7_75t_SL g30319 (.A1(n_23010),
    .A2(n_23012),
    .B(n_12990),
    .Y(n_23014));
 NAND2xp5_ASAP7_75t_SL g30320 (.A(n_23009),
    .B(n_19971),
    .Y(n_23010));
 INVxp67_ASAP7_75t_SL g30321 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_280),
    .Y(n_23009));
 NAND2xp5_ASAP7_75t_SL g30322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_280),
    .B(n_23011),
    .Y(n_23012));
 INVx1_ASAP7_75t_SL g30323 (.A(n_19971),
    .Y(n_23011));
 INVx1_ASAP7_75t_SL g30324 (.A(n_24102),
    .Y(n_12990));
 NAND2xp5_ASAP7_75t_SL g30327 (.A(n_23020),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_242),
    .Y(n_23021));
 INVxp67_ASAP7_75t_SL g30328 (.A(n_23019),
    .Y(n_23020));
 XNOR2xp5_ASAP7_75t_SL g30329 (.A(n_11325),
    .B(n_23018),
    .Y(n_23019));
 XNOR2x1_ASAP7_75t_SL g30330 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_156),
    .Y(n_23018),
    .A(n_12279));
 OAI321xp33_ASAP7_75t_SL g30339 (.A1(n_23031),
    .A2(n_13090),
    .A3(n_7618),
    .B1(n_7619),
    .B2(n_23031),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_281),
    .Y(n_23032));
 NOR2x1_ASAP7_75t_SL g30340 (.A(n_9126),
    .B(n_15353),
    .Y(n_23031));
 XNOR2x1_ASAP7_75t_SL g30341 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_246),
    .Y(n_15353),
    .A(n_10999));
 XNOR2xp5_ASAP7_75t_SL g30342 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_194),
    .B(n_23035),
    .Y(n_23036));
 XOR2xp5_ASAP7_75t_SL g30343 (.A(n_19722),
    .B(n_23033),
    .Y(n_23035));
 NAND2xp5_ASAP7_75t_SL g30345 (.A(n_15192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32),
    .Y(n_23033));
 XNOR2xp5_ASAP7_75t_SL g30349 (.A(n_23076),
    .B(n_23078),
    .Y(n_23079));
 AOI21xp5_ASAP7_75t_SL g30350 (.A1(n_23073),
    .A2(n_23074),
    .B(n_23075),
    .Y(n_23076));
 INVx1_ASAP7_75t_SL g30351 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_135),
    .Y(n_23073));
 INVx1_ASAP7_75t_SL g30352 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_120),
    .Y(n_23074));
 NOR2xp33_ASAP7_75t_SL g30353 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_121),
    .Y(n_23075));
 XNOR2x1_ASAP7_75t_SL g30354 (.B(n_23077),
    .Y(n_23078),
    .A(n_9471));
 INVx1_ASAP7_75t_L g30355 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_91),
    .Y(n_23077));
 NAND2xp5_ASAP7_75t_SL g30357 (.A(n_23079),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_180),
    .Y(n_23083));
 MAJIxp5_ASAP7_75t_SL g30358 (.A(n_23084),
    .B(n_22562),
    .C(n_23085),
    .Y(n_23086));
 INVxp67_ASAP7_75t_SRAM g30359 (.A(n_23078),
    .Y(n_23084));
 XNOR2x1_ASAP7_75t_SL g30360 (.B(n_23091),
    .Y(n_23092),
    .A(n_23087));
 XNOR2xp5_ASAP7_75t_SL g30361 (.A(n_23088),
    .B(n_23090),
    .Y(n_23091));
 MAJx2_ASAP7_75t_SL g30362 (.A(n_18432),
    .B(n_18431),
    .C(n_18430),
    .Y(n_23088));
 XOR2xp5_ASAP7_75t_SL g30363 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_248),
    .Y(n_23090));
 MAJx2_ASAP7_75t_SL g30365 (.A(n_7710),
    .B(n_23093),
    .C(n_23094),
    .Y(n_23095));
 INVxp67_ASAP7_75t_SL g30366 (.A(n_23088),
    .Y(n_23093));
 INVxp67_ASAP7_75t_SRAM g30367 (.A(n_23090),
    .Y(n_23094));
 NAND2xp5_ASAP7_75t_SL g30368 (.A(n_14137),
    .B(n_23101),
    .Y(n_23102));
 XNOR2xp5_ASAP7_75t_SL g30369 (.A(n_23097),
    .B(n_23100),
    .Y(n_23101));
 XNOR2xp5_ASAP7_75t_SL g30370 (.A(n_26035),
    .B(n_26121),
    .Y(n_23097));
 AOI22xp5_ASAP7_75t_SL g30372 (.A1(n_23098),
    .A2(n_9686),
    .B1(n_23099),
    .B2(n_19249),
    .Y(n_23100));
 INVx1_ASAP7_75t_SL g30373 (.A(n_19249),
    .Y(n_23098));
 INVx1_ASAP7_75t_SL g30374 (.A(n_9686),
    .Y(n_23099));
 NOR2xp67_ASAP7_75t_SL g30375 (.A(n_14137),
    .B(n_23101),
    .Y(n_23103));
 MAJx2_ASAP7_75t_SL g30376 (.A(n_23104),
    .B(n_9687),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_224),
    .Y(n_23105));
 INVx1_ASAP7_75t_SL g30377 (.A(n_23097),
    .Y(n_23104));
 XNOR2xp5_ASAP7_75t_SL g30378 (.A(n_13451),
    .B(n_23111),
    .Y(n_23112));
 XNOR2x1_ASAP7_75t_SL g30379 (.B(n_23110),
    .Y(n_23111),
    .A(n_23108));
 OAI22xp5_ASAP7_75t_SL g30380 (.A1(n_23106),
    .A2(n_20888),
    .B1(n_20887),
    .B2(n_20893),
    .Y(n_23108));
 NAND2x1p5_ASAP7_75t_SL g30382 (.A(n_23109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_107),
    .Y(n_23110));
 BUFx2_ASAP7_75t_SL g30383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_96),
    .Y(n_23109));
 MAJIxp5_ASAP7_75t_SL g30384 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_191),
    .B(n_13451),
    .C(n_23111),
    .Y(n_23113));
 OAI21x1_ASAP7_75t_SL g30385 (.A1(n_23114),
    .A2(n_23115),
    .B(n_23116),
    .Y(n_19647));
 INVx1_ASAP7_75t_SL g30386 (.A(n_23110),
    .Y(n_23114));
 NOR2xp33_ASAP7_75t_SL g30387 (.A(n_20887),
    .B(n_20893),
    .Y(n_23115));
 NAND2xp5_ASAP7_75t_SL g30388 (.A(n_20887),
    .B(n_20893),
    .Y(n_23116));
 OAI21xp5_ASAP7_75t_SL g30389 (.A1(n_23121),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_285),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_292),
    .Y(n_23122));
 AO21x1_ASAP7_75t_SL g30390 (.A1(n_11267),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_266),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_264),
    .Y(n_23118));
 NAND2xp5_ASAP7_75t_SL g30391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_248),
    .B(n_4199),
    .Y(n_23119));
 AND2x2_ASAP7_75t_SL g30392 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_275),
    .Y(n_23120));
 OAI22xp33_ASAP7_75t_SL g30393 (.A1(n_23123),
    .A2(n_23126),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_304),
    .B2(n_23121),
    .Y(n_23127));
 INVxp67_ASAP7_75t_SL g30394 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_304),
    .Y(n_23126));
 NAND2xp5_ASAP7_75t_SL g30395 (.A(n_23119),
    .B(n_23129),
    .Y(n_23130));
 INVxp67_ASAP7_75t_SL g30396 (.A(n_23120),
    .Y(n_23129));
 HB1xp67_ASAP7_75t_SL g30397 (.A(n_23118),
    .Y(n_23131));
 XNOR2xp5_ASAP7_75t_SL g304 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_274),
    .B(n_9903),
    .Y(n_7903));
 XNOR2xp5_ASAP7_75t_SL g30400 (.A(n_23133),
    .B(n_23134),
    .Y(n_23135));
 NAND2xp5_ASAP7_75t_SL g30401 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .Y(n_23133));
 OAI22xp5_ASAP7_75t_SL g30402 (.A1(n_18756),
    .A2(n_4044),
    .B1(n_9759),
    .B2(n_9757),
    .Y(n_23134));
 MAJx2_ASAP7_75t_SL g30403 (.A(n_23135),
    .B(n_19821),
    .C(n_3463),
    .Y(n_23138));
 MAJx2_ASAP7_75t_SL g30404 (.A(n_4044),
    .B(n_23133),
    .C(n_9757),
    .Y(n_23139));
 XNOR2xp5_ASAP7_75t_SL g30429 (.A(n_23167),
    .B(n_23168),
    .Y(n_23169));
 XOR2xp5_ASAP7_75t_SL g30430 (.A(n_23165),
    .B(n_23166),
    .Y(n_23167));
 MAJx2_ASAP7_75t_SL g30431 (.A(n_12712),
    .B(n_12708),
    .C(n_22068),
    .Y(n_23165));
 XNOR2xp5_ASAP7_75t_SL g30432 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_151),
    .B(n_11348),
    .Y(n_23166));
 XNOR2xp5_ASAP7_75t_SL g30433 (.A(n_21422),
    .B(n_20248),
    .Y(n_23168));
 XNOR2xp5_ASAP7_75t_SL g30434 (.A(n_23170),
    .B(n_23837),
    .Y(n_23174));
 AOI21xp5_ASAP7_75t_SL g30435 (.A1(n_22536),
    .A2(n_22542),
    .B(n_22543),
    .Y(n_23170));
 INVx2_ASAP7_75t_SL g30437 (.A(n_11819),
    .Y(n_7378));
 MAJIxp5_ASAP7_75t_SL g30439 (.A(n_20720),
    .B(n_8689),
    .C(n_20721),
    .Y(n_23175));
 INVxp67_ASAP7_75t_SL g30440 (.A(n_23170),
    .Y(n_4072));
 INVxp67_ASAP7_75t_SL g30441 (.A(n_23837),
    .Y(n_7370));
 MAJIxp5_ASAP7_75t_SL g30455 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_192),
    .B(n_3459),
    .C(n_23194),
    .Y(n_23195));
 INVxp67_ASAP7_75t_SRAM g30456 (.A(n_23193),
    .Y(n_23194));
 XNOR2x1_ASAP7_75t_SL g30457 (.B(n_23192),
    .Y(n_23193),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_108));
 XNOR2x1_ASAP7_75t_SL g30458 (.B(n_20696),
    .Y(n_23192),
    .A(n_19764));
 XOR2xp5_ASAP7_75t_SL g30459 (.A(n_23193),
    .B(n_23196),
    .Y(n_23197));
 INVx1_ASAP7_75t_SL g30460 (.A(n_8582),
    .Y(n_23196));
 AOI21x1_ASAP7_75t_SL g30479 (.A1(n_23222),
    .A2(n_13623),
    .B(n_23227),
    .Y(n_23228));
 NOR2xp67_ASAP7_75t_SL g30480 (.A(n_23220),
    .B(n_23221),
    .Y(n_23222));
 NAND2xp5_ASAP7_75t_SL g30481 (.A(n_23219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_284),
    .Y(n_23220));
 NAND2xp5_ASAP7_75t_SL g30482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_271),
    .B(n_20853),
    .Y(n_23219));
 NAND2xp5_ASAP7_75t_SL g30483 (.A(n_14024),
    .B(n_14025),
    .Y(n_23221));
 OAI21xp5_ASAP7_75t_SL g30484 (.A1(n_23221),
    .A2(n_23225),
    .B(n_23226),
    .Y(n_23227));
 AOI21xp5_ASAP7_75t_SL g30485 (.A1(n_23223),
    .A2(n_23219),
    .B(n_23224),
    .Y(n_23225));
 NOR2xp33_ASAP7_75t_SL g30486 (.A(n_13530),
    .B(n_7749),
    .Y(n_23223));
 NOR2xp33_ASAP7_75t_SL g30487 (.A(n_20853),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_271),
    .Y(n_23224));
 AOI21xp5_ASAP7_75t_SL g30488 (.A1(n_7531),
    .A2(n_14025),
    .B(n_7540),
    .Y(n_23226));
 AOI21x1_ASAP7_75t_SL g30489 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_309),
    .A2(n_13623),
    .B(n_23229),
    .Y(n_23230));
 INVxp67_ASAP7_75t_SL g30490 (.A(n_23225),
    .Y(n_23229));
 NOR2xp33_ASAP7_75t_L g30491 (.A(n_23231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_285),
    .Y(n_23232));
 NOR2xp33_ASAP7_75t_SL g30492 (.A(n_7749),
    .B(n_13530),
    .Y(n_23231));
 INVxp67_ASAP7_75t_SL g30493 (.A(n_23231),
    .Y(n_23233));
 NOR2xp33_ASAP7_75t_SL g30494 (.A(n_23234),
    .B(n_23235),
    .Y(n_23236));
 NOR2xp33_ASAP7_75t_SRAM g30495 (.A(n_20853),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_271),
    .Y(n_23234));
 INVxp67_ASAP7_75t_SRAM g30496 (.A(n_23219),
    .Y(n_23235));
 MAJIxp5_ASAP7_75t_R g305 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_45),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_29),
    .Y(n_6954));
 OAI22xp5_ASAP7_75t_SL g305_0 (.A1(n_13456),
    .A2(n_10778),
    .B1(n_19830),
    .B2(n_19831),
    .Y(n_19832));
 INVxp67_ASAP7_75t_SL g306 (.A(n_25963),
    .Y(n_19829));
 NOR3xp33_ASAP7_75t_SL g30605 (.A(n_21837),
    .B(n_23367),
    .C(n_21842),
    .Y(n_23368));
 INVx1_ASAP7_75t_SL g30606 (.A(n_23366),
    .Y(n_23367));
 NAND2xp5_ASAP7_75t_SL g30607 (.A(n_21832),
    .B(n_23365),
    .Y(n_23366));
 XNOR2xp5_ASAP7_75t_SL g30608 (.A(n_14059),
    .B(n_9642),
    .Y(n_23365));
 OAI22xp5_ASAP7_75t_SL g30609 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_219),
    .A2(n_23373),
    .B1(n_23374),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_26),
    .Y(n_23375));
 MAJIxp5_ASAP7_75t_SL g30610 (.A(n_23372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_172),
    .C(n_19664),
    .Y(n_23373));
 INVx1_ASAP7_75t_SL g30611 (.A(n_26168),
    .Y(n_23372));
 XNOR2x1_ASAP7_75t_SL g30619 (.B(n_6327),
    .Y(n_23380),
    .A(n_23379));
 XNOR2x1_ASAP7_75t_SL g30620 (.B(n_22437),
    .Y(n_23379),
    .A(n_23378));
 INVx1_ASAP7_75t_SL g30621 (.A(n_9354),
    .Y(n_23378));
 MAJIxp5_ASAP7_75t_SL g30623 (.A(n_14721),
    .B(n_21513),
    .C(n_23386),
    .Y(n_23387));
 XNOR2x1_ASAP7_75t_SL g30624 (.B(n_23385),
    .Y(n_23386),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_126));
 AOI22x1_ASAP7_75t_SL g30625 (.A1(n_21801),
    .A2(n_21800),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_91),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_92),
    .Y(n_23385));
 INVx1_ASAP7_75t_SL g30627 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_92),
    .Y(n_21800));
 HB1xp67_ASAP7_75t_SL g30628 (.A(n_23391),
    .Y(n_23392));
 XNOR2xp5_ASAP7_75t_SL g30629 (.A(n_8053),
    .B(n_23390),
    .Y(n_23391));
 INVxp67_ASAP7_75t_SL g30630 (.A(n_23389),
    .Y(n_23390));
 OA21x2_ASAP7_75t_SL g30631 (.A1(n_10847),
    .A2(n_20938),
    .B(n_23388),
    .Y(n_23389));
 NAND2xp5_ASAP7_75t_SL g30632 (.A(n_10506),
    .B(n_20939),
    .Y(n_23388));
 INVx2_ASAP7_75t_SL g30633 (.A(n_23389),
    .Y(n_23393));
 XNOR2xp5_ASAP7_75t_SL g30634 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_205),
    .B(n_26170),
    .Y(n_23398));
 MAJIxp5_ASAP7_75t_SL g30636 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_36),
    .Y(n_23394));
 XOR2x2_ASAP7_75t_SL g30639 (.A(n_23402),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_44),
    .Y(n_23403));
 OAI22xp5_ASAP7_75t_SL g30640 (.A1(n_23401),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_40),
    .B1(n_23400),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_41),
    .Y(n_23402));
 INVxp67_ASAP7_75t_SL g30641 (.A(n_23400),
    .Y(n_23401));
 AND2x4_ASAP7_75t_SL g30642 (.A(n_23399),
    .B(n_18031),
    .Y(n_23400));
 XNOR2x1_ASAP7_75t_SL g30644 (.B(n_18776),
    .Y(n_23408),
    .A(n_23407));
 XNOR2xp5_ASAP7_75t_SL g30645 (.A(n_26247),
    .B(n_22186),
    .Y(n_23407));
 AND2x2_ASAP7_75t_SL g30647 (.A(n_19682),
    .B(n_26005),
    .Y(n_23404));
 XNOR2xp5_ASAP7_75t_SL g30649 (.A(n_23414),
    .B(n_10465),
    .Y(n_23415));
 XNOR2xp5_ASAP7_75t_SL g30650 (.A(n_23410),
    .B(n_23413),
    .Y(n_23414));
 INVxp67_ASAP7_75t_SL g30651 (.A(n_23409),
    .Y(n_23410));
 INVx1_ASAP7_75t_SL g30652 (.A(n_26053),
    .Y(n_23409));
 OAI22xp5_ASAP7_75t_SL g30653 (.A1(n_23411),
    .A2(n_15384),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_147),
    .B2(n_23412),
    .Y(n_23413));
 INVx1_ASAP7_75t_SL g30654 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_147),
    .Y(n_23411));
 INVx1_ASAP7_75t_SL g30655 (.A(n_15384),
    .Y(n_23412));
 OAI22xp33_ASAP7_75t_SL g30656 (.A1(n_15384),
    .A2(n_26053),
    .B1(n_23412),
    .B2(n_23409),
    .Y(n_23416));
 MAJIxp5_ASAP7_75t_SL g30657 (.A(n_9811),
    .B(n_23422),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_579),
    .Y(n_23423));
 AOI21x1_ASAP7_75t_SL g30658 (.A1(n_23418),
    .A2(n_23420),
    .B(n_23421),
    .Y(n_23422));
 NAND2xp67_ASAP7_75t_SL g30659 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_225),
    .B(n_23417),
    .Y(n_23418));
 INVx1_ASAP7_75t_SL g30660 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_330),
    .Y(n_23417));
 NAND2xp5_ASAP7_75t_SL g30661 (.A(n_23419),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_330),
    .Y(n_23420));
 INVx1_ASAP7_75t_SRAM g30662 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_225),
    .Y(n_23419));
 INVx1_ASAP7_75t_SL g30663 (.A(n_2163),
    .Y(n_23421));
 OAI21x1_ASAP7_75t_SL g30664 (.A1(n_11168),
    .A2(n_23425),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_86),
    .Y(n_23426));
 NOR2xp33_ASAP7_75t_SL g30665 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_651),
    .B(n_23424),
    .Y(n_23425));
 AND2x4_ASAP7_75t_SL g30666 (.A(n_9661),
    .B(n_10538),
    .Y(n_23424));
 MAJIxp5_ASAP7_75t_SL g30667 (.A(n_23430),
    .B(n_8438),
    .C(n_8437),
    .Y(n_23431));
 MAJx2_ASAP7_75t_SL g30668 (.A(n_23427),
    .B(n_23428),
    .C(n_23429),
    .Y(n_23430));
 INVx1_ASAP7_75t_SL g30669 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_1),
    .Y(n_23427));
 INVx1_ASAP7_75t_SL g30670 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_103),
    .Y(n_23428));
 MAJx2_ASAP7_75t_SL g30671 (.A(n_12924),
    .B(n_12926),
    .C(n_12927),
    .Y(n_23429));
 INVx1_ASAP7_75t_SL g30672 (.A(n_23429),
    .Y(n_23432));
 OAI21xp5_ASAP7_75t_SL g30673 (.A1(n_23434),
    .A2(n_23435),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_270),
    .Y(n_23436));
 OA21x2_ASAP7_75t_SL g30674 (.A1(n_11487),
    .A2(n_23433),
    .B(n_21258),
    .Y(n_23434));
 AO21x2_ASAP7_75t_SL g30675 (.A1(n_11475),
    .A2(n_11476),
    .B(n_11477),
    .Y(n_23433));
 HB1xp67_ASAP7_75t_SL g30676 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_272),
    .Y(n_23435));
 NAND2x1_ASAP7_75t_SL g30677 (.A(n_23442),
    .B(n_23444),
    .Y(n_23445));
 OA22x2_ASAP7_75t_SL g30678 (.A1(n_23439),
    .A2(n_21593),
    .B1(n_23441),
    .B2(n_21596),
    .Y(n_23442));
 OR3x1_ASAP7_75t_SL g30679 (.A(n_23437),
    .B(n_12923),
    .C(n_23438),
    .Y(n_23439));
 NOR2xp33_ASAP7_75t_SL g30680 (.A(n_14688),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_268),
    .Y(n_23437));
 INVx1_ASAP7_75t_SL g30681 (.A(n_2182),
    .Y(n_23438));
 NAND2xp5_ASAP7_75t_SL g30682 (.A(n_2182),
    .B(n_23440),
    .Y(n_23441));
 INVxp67_ASAP7_75t_SL g30683 (.A(n_23437),
    .Y(n_23440));
 OAI211xp5_ASAP7_75t_SL g30684 (.A1(n_21593),
    .A2(n_12923),
    .B(n_21596),
    .C(n_23443),
    .Y(n_23444));
 NOR2xp33_ASAP7_75t_SL g30685 (.A(n_23438),
    .B(n_23440),
    .Y(n_23443));
 XNOR2x1_ASAP7_75t_SL g30686 (.B(n_23449),
    .Y(n_23450),
    .A(n_15060));
 XNOR2x1_ASAP7_75t_SL g30687 (.B(n_23448),
    .Y(n_23449),
    .A(n_23447));
 XNOR2x1_ASAP7_75t_SL g30688 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_133),
    .Y(n_23447),
    .A(n_23446));
 INVx1_ASAP7_75t_SL g30689 (.A(n_18771),
    .Y(n_23446));
 XOR2x2_ASAP7_75t_SL g30690 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_4),
    .B(n_9048),
    .Y(n_23448));
 MAJIxp5_ASAP7_75t_SL g30691 (.A(n_11515),
    .B(n_23447),
    .C(n_23448),
    .Y(n_23451));
 OAI21x1_ASAP7_75t_SL g307 (.A1(n_18730),
    .A2(n_4783),
    .B(n_6396),
    .Y(n_6397));
 XNOR2x1_ASAP7_75t_SL g30703 (.B(n_23462),
    .Y(n_23463),
    .A(n_23461));
 XNOR2x1_ASAP7_75t_SL g30704 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_645),
    .Y(n_23462),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_613));
 NAND2xp5_ASAP7_75t_SL g30706 (.A(n_23469),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_61),
    .Y(n_23470));
 INVx1_ASAP7_75t_SL g30707 (.A(n_23468),
    .Y(n_23469));
 NAND2xp5_ASAP7_75t_SL g30708 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(n_23468));
 OAI22xp5_ASAP7_75t_SL g30709 (.A1(n_23468),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_60),
    .B1(n_23469),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_61),
    .Y(n_23471));
 XNOR2xp5_ASAP7_75t_SL g30771 (.A(n_14172),
    .B(n_26172),
    .Y(n_23541));
 MAJIxp5_ASAP7_75t_SL g30779 (.A(n_19950),
    .B(n_23548),
    .C(n_8776),
    .Y(n_23549));
 INVxp67_ASAP7_75t_SL g30780 (.A(n_23547),
    .Y(n_23548));
 XOR2xp5_ASAP7_75t_SL g30781 (.A(n_23546),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_94),
    .Y(n_23547));
 XNOR2x1_ASAP7_75t_SL g30782 (.B(n_5849),
    .Y(n_23546),
    .A(n_19552));
 XNOR2xp5_ASAP7_75t_SL g30783 (.A(n_8777),
    .B(n_23547),
    .Y(n_23550));
 OAI21x1_ASAP7_75t_SL g30784 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_81),
    .A2(n_23546),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_80),
    .Y(n_23551));
 XOR2x2_ASAP7_75t_SL g30785 (.A(n_23554),
    .B(n_19894),
    .Y(n_23555));
 OAI22xp5_ASAP7_75t_SL g30786 (.A1(n_19892),
    .A2(n_23552),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_110),
    .B2(n_23553),
    .Y(n_23554));
 NAND2x1p5_ASAP7_75t_SL g30787 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(n_19645),
    .Y(n_23552));
 INVx1_ASAP7_75t_SL g30788 (.A(n_23552),
    .Y(n_23553));
 OAI21x1_ASAP7_75t_SL g30789 (.A1(n_19893),
    .A2(n_19894),
    .B(n_23557),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_163));
 NAND2xp5_ASAP7_75t_SL g30790 (.A(n_23552),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_110),
    .Y(n_23557));
 NOR2x1_ASAP7_75t_SL g30792 (.A(n_7601),
    .B(n_23563),
    .Y(n_23564));
 AO21x2_ASAP7_75t_SL g30793 (.A1(n_23560),
    .A2(n_9520),
    .B(n_23562),
    .Y(n_23563));
 NOR2xp33_ASAP7_75t_SL g30794 (.A(n_23559),
    .B(n_9518),
    .Y(n_23560));
 INVxp67_ASAP7_75t_SL g30795 (.A(n_2161),
    .Y(n_23559));
 NOR2xp67_ASAP7_75t_SL g30796 (.A(n_23561),
    .B(n_9520),
    .Y(n_23562));
 NAND2xp5_ASAP7_75t_SL g30797 (.A(n_2161),
    .B(n_9518),
    .Y(n_23561));
 NAND2xp5_ASAP7_75t_SL g30798 (.A(n_23563),
    .B(n_23565),
    .Y(n_23566));
 INVx2_ASAP7_75t_SL g30799 (.A(n_7598),
    .Y(n_23565));
 AO21x1_ASAP7_75t_SL g308 (.A1(n_19241),
    .A2(n_24978),
    .B(n_6391),
    .Y(n_6392));
 OAI22xp5_ASAP7_75t_SL g30800 (.A1(n_23565),
    .A2(n_23563),
    .B1(n_23567),
    .B2(n_7598),
    .Y(n_23568));
 INVx1_ASAP7_75t_SL g30801 (.A(n_23563),
    .Y(n_23567));
 NAND2xp5_ASAP7_75t_SL g30803 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(n_23569));
 NOR2x1_ASAP7_75t_SL g30806 (.A(n_23569),
    .B(n_22962),
    .Y(n_23573));
 AO21x2_ASAP7_75t_SL g30811 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .A2(n_23579),
    .B(n_20276),
    .Y(n_23580));
 NOR2xp33_ASAP7_75t_SL g30812 (.A(n_9986),
    .B(n_23578),
    .Y(n_23579));
 NAND2xp5_ASAP7_75t_SL g30813 (.A(n_22786),
    .B(n_10338),
    .Y(n_23578));
 AOI21xp5_ASAP7_75t_SL g30814 (.A1(n_23581),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .B(n_20277),
    .Y(n_23582));
 AND2x2_ASAP7_75t_SL g30890 (.A(n_2985),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .Y(n_23658));
 AND2x4_ASAP7_75t_SL g30891 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(n_16763),
    .Y(n_23659));
 NAND2x1_ASAP7_75t_SL g30892 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B(n_19391),
    .Y(n_23660));
 OAI22xp5_ASAP7_75t_SL g30893 (.A1(n_23663),
    .A2(n_5954),
    .B1(n_5953),
    .B2(n_23662),
    .Y(n_23664));
 INVx1_ASAP7_75t_SL g30894 (.A(n_23662),
    .Y(n_23663));
 XNOR2x1_ASAP7_75t_SL g30895 (.B(n_23661),
    .Y(n_23662),
    .A(n_23658));
 XNOR2x1_ASAP7_75t_SL g30896 (.B(n_23659),
    .Y(n_23661),
    .A(n_23660));
 MAJIxp5_ASAP7_75t_SL g30897 (.A(n_23662),
    .B(n_5954),
    .C(n_5955),
    .Y(n_23665));
 MAJx2_ASAP7_75t_SL g30898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .B(n_23667),
    .C(n_23669),
    .Y(n_23670));
 INVxp67_ASAP7_75t_SL g30899 (.A(n_23666),
    .Y(n_23667));
 AOI21x1_ASAP7_75t_SL g309 (.A1(n_4784),
    .A2(n_6399),
    .B(n_6400),
    .Y(n_6401));
 AND2x2_ASAP7_75t_SL g30900 (.A(n_7595),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_652),
    .Y(n_23666));
 INVxp67_ASAP7_75t_SL g30901 (.A(n_23668),
    .Y(n_23669));
 XNOR2xp5_ASAP7_75t_SL g30913 (.A(n_11142),
    .B(n_18967),
    .Y(n_23682));
 MAJIxp5_ASAP7_75t_SL g30914 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_89),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_80),
    .Y(n_23683));
 OR2x2_ASAP7_75t_SL g30967 (.A(n_24684),
    .B(n_23975),
    .Y(n_23738));
 NAND2x1_ASAP7_75t_SL g31 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(n_2325),
    .Y(n_8781));
 NOR2xp67_ASAP7_75t_SL g310 (.A(n_6394),
    .B(n_6395),
    .Y(n_6396));
 OR2x2_ASAP7_75t_SL g31000 (.A(n_26250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_275),
    .Y(n_23776));
 AND2x2_ASAP7_75t_SL g31003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_185),
    .Y(n_23772));
 NAND2xp5_ASAP7_75t_SL g31044 (.A(n_23818),
    .B(n_23819),
    .Y(n_23820));
 AOI21xp5_ASAP7_75t_SL g31045 (.A1(n_8800),
    .A2(n_8802),
    .B(n_8803),
    .Y(n_23818));
 NAND2xp5_ASAP7_75t_SL g31046 (.A(n_17075),
    .B(n_6730),
    .Y(n_23819));
 INVx1_ASAP7_75t_SL g31050 (.A(n_23824),
    .Y(n_23825));
 NAND2x1_ASAP7_75t_SL g31051 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .B(n_24402),
    .Y(n_23824));
 AOI21xp33_ASAP7_75t_SL g31055 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_319),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_217),
    .B(n_19230),
    .Y(n_23829));
 OAI21x1_ASAP7_75t_SL g31056 (.A1(n_20773),
    .A2(n_22959),
    .B(n_20778),
    .Y(n_23830));
 OAI22xp5_ASAP7_75t_SL g31057 (.A1(n_23833),
    .A2(n_12245),
    .B1(n_19530),
    .B2(n_23834),
    .Y(n_23835));
 AO22x2_ASAP7_75t_SL g31058 (.A1(n_20782),
    .A2(n_23832),
    .B1(n_23829),
    .B2(n_23830),
    .Y(n_23833));
 INVxp67_ASAP7_75t_SL g31060 (.A(n_23829),
    .Y(n_23832));
 AOI22x1_ASAP7_75t_SL g31062 (.A1(n_7378),
    .A2(n_23834),
    .B1(n_11819),
    .B2(n_23833),
    .Y(n_23837));
 INVx2_ASAP7_75t_SL g31063 (.A(n_23833),
    .Y(n_23834));
 OAI22xp33_ASAP7_75t_SL g311 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_266),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_265),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_253),
    .B2(n_10220),
    .Y(n_6395));
 AOI21xp5_ASAP7_75t_SL g31120 (.A1(n_24166),
    .A2(n_23894),
    .B(n_17663),
    .Y(n_23895));
 BUFx3_ASAP7_75t_SL g31121 (.A(n_24167),
    .Y(n_23894));
 NAND2xp5_ASAP7_75t_SL g31157 (.A(n_21881),
    .B(n_21883),
    .Y(n_23931));
 AND2x6_ASAP7_75t_SL g31158 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_pvld[7]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_pvld[7]),
    .Y(n_23932));
 OAI22xp5_ASAP7_75t_SL g31159 (.A1(n_26144),
    .A2(n_23934),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[12]),
    .B2(n_23932),
    .Y(n_23935));
 OAI21xp33_ASAP7_75t_SL g31160 (.A1(n_25833),
    .A2(n_23931),
    .B(n_23932),
    .Y(n_23934));
 INVx1_ASAP7_75t_SL g31163 (.A(n_14998),
    .Y(n_23936));
 XNOR2xp5_ASAP7_75t_SL g31167 (.A(n_23942),
    .B(n_25296),
    .Y(n_9827));
 INVxp67_ASAP7_75t_SL g31168 (.A(n_23941),
    .Y(n_23942));
 MAJIxp5_ASAP7_75t_SL g31169 (.A(n_15719),
    .B(n_15720),
    .C(n_12834),
    .Y(n_23941));
 XNOR2xp5_ASAP7_75t_SL g31196 (.A(n_6045),
    .B(n_8057),
    .Y(n_23972));
 MAJIxp5_ASAP7_75t_SL g31197 (.A(n_12186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_51),
    .C(n_23974),
    .Y(n_23975));
 XOR2xp5_ASAP7_75t_SL g31198 (.A(n_23973),
    .B(n_23972),
    .Y(n_23974));
 XOR2xp5_ASAP7_75t_L g31199 (.A(n_19790),
    .B(n_19865),
    .Y(n_23973));
 MAJIxp5_ASAP7_75t_SL g312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_267),
    .B(n_4068),
    .C(n_21667),
    .Y(n_21668));
 XOR2xp5_ASAP7_75t_SL g31210 (.A(n_23985),
    .B(n_23986),
    .Y(n_23987));
 MAJIxp5_ASAP7_75t_SL g31211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_753),
    .B(n_11904),
    .C(n_22042),
    .Y(n_23985));
 XNOR2xp5_ASAP7_75t_SL g31212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_783),
    .B(n_9726),
    .Y(n_23986));
 INVx1_ASAP7_75t_SL g31213 (.A(n_23986),
    .Y(n_23988));
 AOI22xp5_ASAP7_75t_SL g31247 (.A1(n_24025),
    .A2(n_23936),
    .B1(n_14998),
    .B2(n_24024),
    .Y(n_24027));
 MAJIxp5_ASAP7_75t_SL g31249 (.A(n_12080),
    .B(n_14454),
    .C(n_12077),
    .Y(n_24024));
 MAJIxp5_ASAP7_75t_SL g31251 (.A(n_22321),
    .B(n_24025),
    .C(n_14457),
    .Y(n_24028));
 AOI21xp5_ASAP7_75t_SL g31252 (.A1(n_14457),
    .A2(n_24025),
    .B(n_24022),
    .Y(n_24029));
 MAJIxp5_ASAP7_75t_SL g31255 (.A(n_24033),
    .B(n_8248),
    .C(n_19404),
    .Y(n_24034));
 AOI21xp5_ASAP7_75t_SL g31256 (.A1(n_7170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_241),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_236),
    .Y(n_24033));
 INVx1_ASAP7_75t_SL g31257 (.A(n_24033),
    .Y(n_24035));
 NOR2xp33_ASAP7_75t_SL g313 (.A(n_24979),
    .B(n_18667),
    .Y(n_6404));
 OAI22x1_ASAP7_75t_SL g31320 (.A1(n_24104),
    .A2(n_24105),
    .B1(n_14799),
    .B2(n_24106),
    .Y(n_24107));
 NAND2xp5_ASAP7_75t_SL g31321 (.A(n_24102),
    .B(n_24103),
    .Y(n_24104));
 AND3x2_ASAP7_75t_SL g31322 (.A(n_23932),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .C(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[1]),
    .Y(n_24102));
 INVxp67_ASAP7_75t_SL g31323 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_305),
    .Y(n_24103));
 INVx1_ASAP7_75t_SL g31324 (.A(n_14799),
    .Y(n_24105));
 A2O1A1Ixp33_ASAP7_75t_SL g3133 (.A1(n_15173),
    .A2(n_15181),
    .B(n_15186),
    .C(n_15187),
    .Y(n_15188));
 OAI22xp5_ASAP7_75t_SL g3134 (.A1(n_15169),
    .A2(n_15172),
    .B1(n_19201),
    .B2(n_15185),
    .Y(n_15186));
 NAND2x1_ASAP7_75t_SL g3135 (.A(n_15169),
    .B(n_15172),
    .Y(n_15173));
 NAND2xp5_ASAP7_75t_SL g3136 (.A(n_19201),
    .B(n_15185),
    .Y(n_15187));
 NAND2x1p5_ASAP7_75t_SL g31362 (.A(n_9832),
    .B(n_24152),
    .Y(n_24153));
 BUFx2_ASAP7_75t_SL g31363 (.A(n_9831),
    .Y(n_9832));
 XOR2x2_ASAP7_75t_SL g31364 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_34),
    .B(n_9833),
    .Y(n_24152));
 NAND2xp5_ASAP7_75t_SL g31376 (.A(n_20873),
    .B(n_17661),
    .Y(n_24166));
 OAI21x1_ASAP7_75t_SL g31377 (.A1(n_21434),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .B(n_24153),
    .Y(n_24167));
 AOI21xp5_ASAP7_75t_SL g31378 (.A1(n_24168),
    .A2(n_22087),
    .B(n_16676),
    .Y(n_24169));
 NAND2xp5_ASAP7_75t_SL g31379 (.A(n_24167),
    .B(n_24166),
    .Y(n_24168));
 OAI21xp33_ASAP7_75t_SL g31381 (.A1(n_24172),
    .A2(n_24173),
    .B(n_24175),
    .Y(n_24176));
 NAND2xp5_ASAP7_75t_SL g31382 (.A(n_23580),
    .B(n_24171),
    .Y(n_24172));
 NAND2xp5_ASAP7_75t_SL g31383 (.A(n_5351),
    .B(n_5349),
    .Y(n_24171));
 INVxp67_ASAP7_75t_SL g31384 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_466),
    .Y(n_24173));
 OAI21xp5_ASAP7_75t_SL g31385 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_473),
    .A2(n_24174),
    .B(n_24171),
    .Y(n_24175));
 NAND2xp5_ASAP7_75t_SL g31386 (.A(n_5349),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_24174));
 AOI21xp33_ASAP7_75t_SL g31387 (.A1(n_24178),
    .A2(n_24179),
    .B(n_26037),
    .Y(n_24181));
 NOR2xp33_ASAP7_75t_SL g31388 (.A(n_24177),
    .B(n_11320),
    .Y(n_24178));
 NAND2xp5_ASAP7_75t_SL g31389 (.A(n_5322),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_437),
    .Y(n_24177));
 MAJIxp5_ASAP7_75t_SL g3139 (.A(n_15176),
    .B(n_15178),
    .C(n_15180),
    .Y(n_15181));
 NAND2xp5_ASAP7_75t_SL g31390 (.A(n_22439),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_466),
    .Y(n_24179));
 HB1xp67_ASAP7_75t_SL g314 (.A(n_6394),
    .Y(n_6400));
 XOR2xp5_ASAP7_75t_SL g31407 (.A(n_24200),
    .B(n_24201),
    .Y(n_24202));
 OAI22xp5_ASAP7_75t_SL g31408 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .A2(n_23834),
    .B1(n_23833),
    .B2(n_17414),
    .Y(n_24201));
 AOI21x1_ASAP7_75t_SL g31409 (.A1(n_24203),
    .A2(n_24204),
    .B(n_25450),
    .Y(n_24206));
 MAJIxp5_ASAP7_75t_SL g3141 (.A(n_15164),
    .B(n_15166),
    .C(n_15168),
    .Y(n_15169));
 AO21x2_ASAP7_75t_SL g31410 (.A1(n_22379),
    .A2(n_20623),
    .B(n_21692),
    .Y(n_24203));
 NOR2xp67_ASAP7_75t_SL g31411 (.A(n_20629),
    .B(n_20630),
    .Y(n_24204));
 XNOR2x1_ASAP7_75t_SL g31413 (.B(n_24212),
    .Y(n_24213),
    .A(n_24207));
 INVxp67_ASAP7_75t_SL g31414 (.A(n_26249),
    .Y(n_24212));
 HB1xp67_ASAP7_75t_SL g31417 (.A(n_7379),
    .Y(n_24208));
 OR2x2_ASAP7_75t_SL g31418 (.A(n_2591),
    .B(n_24208),
    .Y(n_24210));
 NOR2xp67_ASAP7_75t_SL g3142 (.A(n_15177),
    .B(n_15179),
    .Y(n_15191));
 XNOR2x1_ASAP7_75t_SL g3143 (.B(n_15171),
    .Y(n_15172),
    .A(n_18094));
 NAND2xp5_ASAP7_75t_SL g31435 (.A(n_2168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_586),
    .Y(n_24230));
 NAND2xp5_ASAP7_75t_SL g3145 (.A(n_15174),
    .B(n_15175),
    .Y(n_15176));
 INVxp67_ASAP7_75t_SL g3147 (.A(n_15179),
    .Y(n_15180));
 XNOR2xp5_ASAP7_75t_SL g3148 (.A(n_15164),
    .B(n_18883),
    .Y(n_15179));
 MAJIxp5_ASAP7_75t_SL g3149 (.A(n_7859),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_9),
    .C(n_4805),
    .Y(n_15174));
 OAI21xp5_ASAP7_75t_SL g315 (.A1(n_10744),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_285),
    .B(n_10741),
    .Y(n_6394));
 HB1xp67_ASAP7_75t_SL g3150 (.A(n_15167),
    .Y(n_15168));
 MAJIxp5_ASAP7_75t_SL g3151 (.A(n_14741),
    .B(n_7297),
    .C(n_7296),
    .Y(n_15167));
 MAJIxp5_ASAP7_75t_SL g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_178),
    .B(n_19571),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_18),
    .Y(n_15171));
 INVx1_ASAP7_75t_SL g3153 (.A(n_15177),
    .Y(n_15178));
 MAJx2_ASAP7_75t_SL g3154 (.A(n_12308),
    .B(n_18699),
    .C(n_5564),
    .Y(n_15177));
 XOR2xp5_ASAP7_75t_SL g3156 (.A(n_7128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_10),
    .Y(n_15164));
 XNOR2xp5_ASAP7_75t_SL g3159 (.A(n_8006),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_216),
    .Y(n_15185));
 INVxp67_ASAP7_75t_SL g316 (.A(n_18667),
    .Y(n_6406));
 XOR2xp5_ASAP7_75t_SL g3160 (.A(n_12308),
    .B(n_12304),
    .Y(n_15175));
 OAI21xp5_ASAP7_75t_SL g31795 (.A1(n_24669),
    .A2(n_24670),
    .B(n_12975),
    .Y(n_24671));
 NOR2xp67_ASAP7_75t_SL g31796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_17),
    .Y(n_24669));
 AOI21x1_ASAP7_75t_SL g31797 (.A1(n_21830),
    .A2(n_23368),
    .B(n_21853),
    .Y(n_24670));
 INVx2_ASAP7_75t_SL g318 (.A(n_21664),
    .Y(n_21665));
 MAJIxp5_ASAP7_75t_SL g31804 (.A(n_22617),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_54),
    .Y(n_24679));
 XNOR2xp5_ASAP7_75t_SL g31805 (.A(n_24682),
    .B(n_24683),
    .Y(n_24684));
 HB1xp67_ASAP7_75t_SL g31806 (.A(n_24681),
    .Y(n_24682));
 OAI22xp5_ASAP7_75t_L g31807 (.A1(n_6323),
    .A2(n_19866),
    .B1(n_23972),
    .B2(n_21939),
    .Y(n_24681));
 OAI22xp5_ASAP7_75t_SL g31808 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .A2(n_6076),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .B2(n_18856),
    .Y(n_24683));
 AO21x2_ASAP7_75t_SL g31834 (.A1(n_24710),
    .A2(n_20236),
    .B(n_24711),
    .Y(n_24712));
 NOR2xp33_ASAP7_75t_SL g31835 (.A(n_19193),
    .B(n_7516),
    .Y(n_24710));
 XNOR2x1_ASAP7_75t_SL g31887 (.B(n_22500),
    .Y(n_24766),
    .A(n_21913));
 MAJx2_ASAP7_75t_SL g31888 (.A(n_9214),
    .B(n_11249),
    .C(n_24768),
    .Y(n_24769));
 XNOR2x2_ASAP7_75t_SL g31889 (.A(n_24767),
    .B(n_24766),
    .Y(n_24768));
 XNOR2xp5_ASAP7_75t_SL g31890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_647),
    .B(n_22097),
    .Y(n_24767));
 XNOR2x1_ASAP7_75t_SL g31891 (.B(n_9447),
    .Y(n_24770),
    .A(n_24768));
 NOR2xp33_ASAP7_75t_SL g319 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_266),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_265),
    .Y(n_6391));
 HB1xp67_ASAP7_75t_SL g32 (.A(n_21793),
    .Y(n_25596));
 AO22x1_ASAP7_75t_SL g320 (.A1(n_20950),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_131),
    .B1(n_20951),
    .B2(n_20953),
    .Y(n_20954));
 NOR2x1_ASAP7_75t_SL g32030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_230),
    .B(n_14344),
    .Y(n_24912));
 NAND2xp5_ASAP7_75t_SL g32031 (.A(n_6353),
    .B(n_6352),
    .Y(n_24913));
 AO21x1_ASAP7_75t_SL g32032 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_268),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_273),
    .B(n_24915),
    .Y(n_24916));
 OAI21xp5_ASAP7_75t_SL g32033 (.A1(n_24912),
    .A2(n_24913),
    .B(n_24914),
    .Y(n_24915));
 NAND2xp5_ASAP7_75t_L g32034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_230),
    .B(n_14344),
    .Y(n_24914));
 AOI321xp33_ASAP7_75t_SL g32035 (.A1(n_6975),
    .A2(n_24915),
    .A3(n_6974),
    .B1(n_6978),
    .B2(n_6974),
    .C(n_6979),
    .Y(n_24917));
 XNOR2xp5_ASAP7_75t_SL g32094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_146),
    .Y(n_24976));
 INVx2_ASAP7_75t_SL g32095 (.A(n_24976),
    .Y(n_24977));
 NAND2xp5_ASAP7_75t_L g32096 (.A(n_10220),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_253),
    .Y(n_24978));
 INVxp67_ASAP7_75t_SL g32097 (.A(n_24978),
    .Y(n_24979));
 INVx1_ASAP7_75t_SL g321 (.A(n_25292),
    .Y(n_25294));
 A2O1A1Ixp33_ASAP7_75t_SL g3218 (.A1(n_19495),
    .A2(n_19496),
    .B(n_19501),
    .C(n_19502),
    .Y(n_19503));
 NAND2xp5_ASAP7_75t_SL g3219 (.A(n_19497),
    .B(n_19500),
    .Y(n_19501));
 OAI21x1_ASAP7_75t_SL g3220 (.A1(n_12503),
    .A2(n_22498),
    .B(n_12504),
    .Y(n_19496));
 OAI21x1_ASAP7_75t_SL g3221 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_283),
    .A2(n_4286),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_282),
    .Y(n_19495));
 NOR2xp33_ASAP7_75t_SL g32218 (.A(n_25128),
    .B(n_25882),
    .Y(n_25130));
 NOR2x1p5_ASAP7_75t_SL g32219 (.A(n_21246),
    .B(n_10933),
    .Y(n_25128));
 INVxp67_ASAP7_75t_SL g3222 (.A(n_19497),
    .Y(n_19504));
 NAND3xp33_ASAP7_75t_SL g3223 (.A(n_22496),
    .B(n_12508),
    .C(n_22497),
    .Y(n_19497));
 NAND2xp5_ASAP7_75t_SL g3224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266),
    .Y(n_19502));
 NAND2xp5_ASAP7_75t_SL g3225 (.A(n_19498),
    .B(n_19499),
    .Y(n_19500));
 NOR2xp33_ASAP7_75t_SRAM g3226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266),
    .Y(n_19505));
 INVxp67_ASAP7_75t_SL g3227 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265),
    .Y(n_19498));
 INVxp67_ASAP7_75t_SL g3228 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266),
    .Y(n_19499));
 INVx1_ASAP7_75t_SL g323 (.A(n_18730),
    .Y(n_6399));
 XOR2xp5_ASAP7_75t_SL g32379 (.A(n_26051),
    .B(n_25295),
    .Y(n_25296));
 AOI22xp5_ASAP7_75t_SL g32380 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .A2(n_25292),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_148),
    .B2(n_25294),
    .Y(n_25295));
 MAJx2_ASAP7_75t_SL g32381 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_627),
    .B(n_18800),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_659),
    .Y(n_25292));
 INVx1_ASAP7_75t_SL g32382 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_148));
 XOR2xp5_ASAP7_75t_SL g32383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_148),
    .B(n_26051),
    .Y(n_25298));
 MAJIxp5_ASAP7_75t_SL g32384 (.A(n_22129),
    .B(n_25301),
    .C(n_21097),
    .Y(n_25302));
 XNOR2x1_ASAP7_75t_SL g32385 (.B(n_25300),
    .Y(n_25301),
    .A(n_25299));
 XNOR2x1_ASAP7_75t_SL g32388 (.B(n_22129),
    .Y(n_25303),
    .A(n_25301));
 XOR2xp5_ASAP7_75t_SL g32396 (.A(n_25311),
    .B(n_25312),
    .Y(n_25313));
 XNOR2xp5_ASAP7_75t_SL g32397 (.A(n_20857),
    .B(n_21394),
    .Y(n_25311));
 OAI22xp5_ASAP7_75t_SL g32398 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_85),
    .A2(n_20285),
    .B1(n_20283),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_86),
    .Y(n_25312));
 NOR2xp33_ASAP7_75t_SL g324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_137),
    .B(n_20949),
    .Y(n_20950));
 XOR2xp5_ASAP7_75t_SL g32418 (.A(n_25335),
    .B(n_25336),
    .Y(n_25337));
 AND2x2_ASAP7_75t_SL g32419 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .Y(n_25335));
 NAND2x1_ASAP7_75t_SL g32420 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(n_4275),
    .Y(n_25336));
 NAND2xp5_ASAP7_75t_SL g32421 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(n_4275),
    .Y(n_20514));
 AND2x2_ASAP7_75t_SL g325 (.A(n_3309),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .Y(n_6569));
 XNOR2xp5_ASAP7_75t_SL g32508 (.A(n_25425),
    .B(n_25428),
    .Y(n_25429));
 XNOR2xp5_ASAP7_75t_SL g32510 (.A(n_25429),
    .B(n_20994),
    .Y(n_25431));
 OR2x2_ASAP7_75t_SL g32524 (.A(n_25981),
    .B(n_25445),
    .Y(n_25446));
 XNOR2xp5_ASAP7_75t_SL g32526 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_343),
    .B(n_16060),
    .Y(n_25445));
 NAND3xp33_ASAP7_75t_SL g32527 (.A(n_25446),
    .B(n_5943),
    .C(n_5944),
    .Y(n_25448));
 NAND2xp5_ASAP7_75t_SL g32528 (.A(n_5383),
    .B(n_25446),
    .Y(n_25449));
 OAI21xp5_ASAP7_75t_SL g32529 (.A1(n_25446),
    .A2(n_20630),
    .B(n_20633),
    .Y(n_25450));
 MAJx2_ASAP7_75t_SL g32581 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_25),
    .B(n_25502),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_156),
    .Y(n_25503));
 MAJx2_ASAP7_75t_SL g32653 (.A(n_8773),
    .B(n_25596),
    .C(n_25597),
    .Y(n_25598));
 BUFx2_ASAP7_75t_L g32654 (.A(n_12250),
    .Y(n_25597));
 INVx1_ASAP7_75t_SL g32655 (.A(n_21793),
    .Y(n_25599));
 MAJIxp5_ASAP7_75t_SL g32658 (.A(n_22989),
    .B(n_7318),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_174),
    .Y(n_25602));
 AOI21x1_ASAP7_75t_SL g32660 (.A1(n_13599),
    .A2(n_25604),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273),
    .Y(n_25605));
 OAI21xp5_ASAP7_75t_SL g3269 (.A1(n_12033),
    .A2(n_12026),
    .B(n_12035),
    .Y(n_12036));
 XOR2xp5_ASAP7_75t_SL g327 (.A(n_8022),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_8),
    .Y(n_8862));
 AOI21xp5_ASAP7_75t_SL g3271 (.A1(n_15559),
    .A2(n_12013),
    .B(n_17559),
    .Y(n_12033));
 OAI21xp5_ASAP7_75t_SL g3273 (.A1(n_12025),
    .A2(n_12026),
    .B(n_12027),
    .Y(n_12028));
 NOR2x1p5_ASAP7_75t_SL g3275 (.A(n_12016),
    .B(n_12017),
    .Y(n_12018));
 NOR2xp33_ASAP7_75t_SL g3276 (.A(n_12017),
    .B(n_12026),
    .Y(n_12038));
 OAI211xp5_ASAP7_75t_SL g3279 (.A1(n_11000),
    .A2(n_10902),
    .B(n_9503),
    .C(n_11872),
    .Y(n_12013));
 AND2x2_ASAP7_75t_SL g3282 (.A(n_7927),
    .B(n_15645),
    .Y(n_12017));
 NOR2x1_ASAP7_75t_SL g3284 (.A(n_7927),
    .B(n_15645),
    .Y(n_12026));
 NOR2xp33_ASAP7_75t_SL g3285 (.A(n_14864),
    .B(n_11220),
    .Y(n_12025));
 INVxp67_ASAP7_75t_SL g3286 (.A(n_12016),
    .Y(n_12027));
 AND2x2_ASAP7_75t_SL g3287 (.A(n_14864),
    .B(n_11220),
    .Y(n_12016));
 AO21x2_ASAP7_75t_SL g32876 (.A1(n_23820),
    .A2(n_21875),
    .B(n_21876),
    .Y(n_25833));
 MAJIxp5_ASAP7_75t_SL g329 (.A(n_10612),
    .B(n_7805),
    .C(n_3358),
    .Y(n_14059));
 INVxp67_ASAP7_75t_SL g32925 (.A(n_25881),
    .Y(n_25882));
 NAND2x1_ASAP7_75t_SL g32926 (.A(n_21246),
    .B(n_10933),
    .Y(n_25881));
 NOR2xp67_ASAP7_75t_SL g32974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_62),
    .Y(n_25963));
 OAI21x1_ASAP7_75t_SL g32982 (.A1(n_22147),
    .A2(n_26237),
    .B(n_21789),
    .Y(n_25971));
 OR2x2_ASAP7_75t_SL g32987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_87),
    .Y(n_25976));
 MAJx2_ASAP7_75t_SL g32988 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_132),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_152),
    .Y(n_25977));
 AND2x2_ASAP7_75t_SL g32989 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(n_2307),
    .Y(n_25978));
 OR2x2_ASAP7_75t_SL g32990 (.A(n_17244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_139),
    .Y(n_25979));
 MAJx2_ASAP7_75t_SL g32991 (.A(n_19878),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_27),
    .C(n_3445),
    .Y(n_25980));
 MAJx2_ASAP7_75t_SL g32992 (.A(n_2578),
    .B(n_15067),
    .C(n_15226),
    .Y(n_25981));
 OR2x2_ASAP7_75t_SL g32993 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_47),
    .Y(n_25982));
 AND2x2_ASAP7_75t_SL g32994 (.A(n_6589),
    .B(n_19808),
    .Y(n_25983));
 AND2x2_ASAP7_75t_SL g32995 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(n_2359),
    .Y(n_25984));
 AND2x2_ASAP7_75t_SL g32998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_282),
    .Y(n_25987));
 AND2x2_ASAP7_75t_SL g32999 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_25988));
 NAND2x1_ASAP7_75t_SL g33 (.A(n_16763),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .Y(n_14671));
 XNOR2xp5_ASAP7_75t_SL g330 (.A(n_14017),
    .B(n_14021),
    .Y(n_14022));
 AND2x2_ASAP7_75t_SL g33000 (.A(n_7508),
    .B(n_7506),
    .Y(n_25989));
 AND2x2_ASAP7_75t_SL g33001 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(n_2307),
    .Y(n_25990));
 MAJx2_ASAP7_75t_SL g33003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_67),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_35),
    .Y(n_25992));
 XOR2xp5_ASAP7_75t_SL g33007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_751),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_12),
    .Y(n_25996));
 AND2x2_ASAP7_75t_SL g33010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_59),
    .Y(n_25999));
 XOR2x2_ASAP7_75t_SL g33011 (.A(n_10613),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_142),
    .Y(n_26000));
 AND2x2_ASAP7_75t_SL g33014 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[63]),
    .Y(n_26003));
 OAI22xp5_ASAP7_75t_SL g33015 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_n_737),
    .A2(n_18964),
    .B1(n_6082),
    .B2(n_6669),
    .Y(n_26004));
 AND2x4_ASAP7_75t_SL g33016 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(n_19391),
    .Y(n_26005));
 NAND2xp5_ASAP7_75t_SL g33019 (.A(n_16769),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .Y(n_26008));
 XOR2x2_ASAP7_75t_SL g33020 (.A(n_19480),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_135),
    .Y(n_26009));
 AND2x2_ASAP7_75t_SL g33021 (.A(n_6209),
    .B(n_6211),
    .Y(n_26010));
 XOR2xp5_ASAP7_75t_SL g33022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_165),
    .B(n_19024),
    .Y(n_26011));
 AND2x2_ASAP7_75t_SL g33023 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .B(n_3868),
    .Y(n_26012));
 AND2x2_ASAP7_75t_SL g33026 (.A(n_5324),
    .B(n_5994),
    .Y(n_26015));
 MAJx2_ASAP7_75t_SL g33027 (.A(n_4038),
    .B(n_13725),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_111),
    .Y(n_26016));
 OA21x2_ASAP7_75t_SL g33028 (.A1(n_10895),
    .A2(n_22983),
    .B(n_26245),
    .Y(n_26017));
 AND2x2_ASAP7_75t_SL g33032 (.A(n_21861),
    .B(n_4826),
    .Y(n_26021));
 MAJx2_ASAP7_75t_SL g33035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_565),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_725),
    .Y(n_26024));
 XOR2xp5_ASAP7_75t_SL g33037 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_35),
    .B(n_8035),
    .Y(n_26026));
 XNOR2xp5_ASAP7_75t_SL g33039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_252),
    .B(n_10742),
    .Y(n_26028));
 AND2x2_ASAP7_75t_SL g33040 (.A(n_19838),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_269),
    .Y(n_26029));
 OR2x2_ASAP7_75t_SL g33041 (.A(n_19840),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_269),
    .Y(n_26030));
 AND2x2_ASAP7_75t_SL g33042 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270),
    .B(n_14177),
    .Y(n_26031));
 XNOR2xp5_ASAP7_75t_SL g33043 (.A(n_22719),
    .B(n_22720),
    .Y(n_26032));
 MAJx2_ASAP7_75t_SL g33044 (.A(n_22725),
    .B(n_22726),
    .C(n_22727),
    .Y(n_26033));
 MAJx2_ASAP7_75t_SL g33046 (.A(n_4231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_149),
    .C(n_26266),
    .Y(n_26035));
 AND2x2_ASAP7_75t_SL g33048 (.A(n_5322),
    .B(n_5324),
    .Y(n_26037));
 OR2x2_ASAP7_75t_SL g33049 (.A(n_21651),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_243),
    .Y(n_26038));
 XNOR2x1_ASAP7_75t_SL g33050 (.B(n_18711),
    .Y(n_26039),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_83));
 XOR2xp5_ASAP7_75t_SL g33051 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_29),
    .B(n_10686),
    .Y(n_26040));
 XNOR2xp5_ASAP7_75t_SL g33052 (.A(n_13097),
    .B(n_23463),
    .Y(n_26041));
 XNOR2xp5_ASAP7_75t_SL g33055 (.A(n_11270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_100),
    .Y(n_26044));
 NOR2xp33_ASAP7_75t_SL g33056 (.A(n_21851),
    .B(n_21842),
    .Y(n_26045));
 XOR2x2_ASAP7_75t_SL g33057 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_147),
    .Y(n_26046));
 XOR2x1_ASAP7_75t_SL g33060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_643),
    .Y(n_26049),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_739));
 XNOR2x2_ASAP7_75t_SL g33062 (.A(n_5806),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_625),
    .Y(n_26051));
 XOR2xp5_ASAP7_75t_SL g33063 (.A(n_20945),
    .B(n_10408),
    .Y(n_26052));
 XNOR2xp5_ASAP7_75t_SL g33064 (.A(n_13769),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_101),
    .Y(n_26053));
 XOR2xp5_ASAP7_75t_SL g33065 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_36),
    .Y(n_26054));
 XOR2xp5_ASAP7_75t_SL g33066 (.A(n_19453),
    .B(n_19454),
    .Y(n_26055));
 XOR2xp5_ASAP7_75t_SL g33068 (.A(n_7025),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_279),
    .Y(n_26057));
 XNOR2xp5_ASAP7_75t_SL g33069 (.A(n_7665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_25),
    .Y(n_26058));
 XNOR2xp5_ASAP7_75t_SL g33070 (.A(n_19146),
    .B(n_7675),
    .Y(n_26059));
 XOR2xp5_ASAP7_75t_SL g33071 (.A(n_7753),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_83),
    .Y(n_26060));
 XOR2xp5_ASAP7_75t_SL g33073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_217),
    .B(n_7854),
    .Y(n_26062));
 XNOR2xp5_ASAP7_75t_SL g33074 (.A(n_7894),
    .B(n_7893),
    .Y(n_26063));
 XOR2xp5_ASAP7_75t_SL g33077 (.A(n_19915),
    .B(n_8732),
    .Y(n_26066));
 XOR2xp5_ASAP7_75t_SL g33079 (.A(n_2437),
    .B(n_14111),
    .Y(n_26068));
 XNOR2xp5_ASAP7_75t_SL g33082 (.A(n_10236),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_205),
    .Y(n_26071));
 XOR2xp5_ASAP7_75t_SL g33084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_174),
    .B(n_10092),
    .Y(n_26073));
 XOR2xp5_ASAP7_75t_SL g33085 (.A(n_18430),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_275),
    .Y(n_26074));
 XNOR2x1_ASAP7_75t_SL g33087 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_649),
    .Y(n_26076),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_617));
 XOR2xp5_ASAP7_75t_SL g33088 (.A(n_11333),
    .B(n_26068),
    .Y(n_26077));
 XOR2x1_ASAP7_75t_SL g33089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_220),
    .Y(n_26078),
    .B(n_22000));
 XOR2xp5_ASAP7_75t_SL g33090 (.A(n_22043),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_753),
    .Y(n_26079));
 XNOR2xp5_ASAP7_75t_SL g33091 (.A(n_26212),
    .B(n_12402),
    .Y(n_26080));
 XOR2xp5_ASAP7_75t_SL g33092 (.A(n_23426),
    .B(n_21489),
    .Y(n_26081));
 XOR2xp5_ASAP7_75t_SL g33094 (.A(n_22477),
    .B(n_13387),
    .Y(n_26083));
 OAI21xp5_ASAP7_75t_SL g331 (.A1(n_14018),
    .A2(n_14019),
    .B(n_14020),
    .Y(n_14021));
 XOR2xp5_ASAP7_75t_SL g33100 (.A(n_18799),
    .B(n_7162),
    .Y(n_26089));
 XOR2xp5_ASAP7_75t_SL g33102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_589),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_685),
    .Y(n_26091));
 XNOR2x1_ASAP7_75t_SL g33104 (.B(n_19310),
    .Y(n_26093),
    .A(n_19306));
 XOR2xp5_ASAP7_75t_SL g33108 (.A(n_19400),
    .B(n_21469),
    .Y(n_26097));
 XNOR2x1_ASAP7_75t_SL g33109 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_79),
    .Y(n_26098),
    .A(n_13245));
 OR2x2_ASAP7_75t_SL g33110 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_87),
    .Y(n_26099));
 XNOR2xp5_ASAP7_75t_SL g33111 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_10),
    .B(n_12414),
    .Y(n_26100));
 XNOR2xp5_ASAP7_75t_SL g33112 (.A(n_19478),
    .B(n_26009),
    .Y(n_26101));
 XNOR2xp5_ASAP7_75t_SL g33113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_111),
    .Y(n_26102));
 XNOR2xp5_ASAP7_75t_SL g33114 (.A(n_22154),
    .B(n_24712),
    .Y(n_26103));
 XNOR2xp5_ASAP7_75t_SL g33116 (.A(n_19647),
    .B(n_18939),
    .Y(n_26105));
 OR2x2_ASAP7_75t_SL g33118 (.A(n_6209),
    .B(n_6211),
    .Y(n_26107));
 OR2x2_ASAP7_75t_SL g33119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_47),
    .Y(n_26108));
 XOR2xp5_ASAP7_75t_SL g33120 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_20),
    .B(n_10073),
    .Y(n_26109));
 XNOR2xp5_ASAP7_75t_SL g33121 (.A(n_19736),
    .B(n_19737),
    .Y(n_26110));
 XOR2xp5_ASAP7_75t_SL g33122 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_137),
    .Y(n_26111));
 XOR2xp5_ASAP7_75t_SL g33123 (.A(n_23036),
    .B(n_8841),
    .Y(n_26112));
 XOR2xp5_ASAP7_75t_SL g33124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_177),
    .B(n_8150),
    .Y(n_26113));
 XOR2xp5_ASAP7_75t_SL g33125 (.A(n_22172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_27),
    .Y(n_26114));
 XNOR2xp5_ASAP7_75t_SL g33128 (.A(n_20096),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_185),
    .Y(n_26117));
 OR2x2_ASAP7_75t_SL g33129 (.A(n_10888),
    .B(n_12576),
    .Y(n_26118));
 XOR2xp5_ASAP7_75t_SL g33130 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_150),
    .B(n_20103),
    .Y(n_26119));
 XNOR2x1_ASAP7_75t_SL g33131 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_79),
    .Y(n_26120),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_72));
 XOR2xp5_ASAP7_75t_SL g33132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_21),
    .Y(n_26121));
 XOR2xp5_ASAP7_75t_SL g33133 (.A(n_20294),
    .B(n_13712),
    .Y(n_26122));
 AND2x2_ASAP7_75t_SL g33134 (.A(n_20365),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_288),
    .Y(n_26123));
 XOR2xp5_ASAP7_75t_SL g33135 (.A(n_5781),
    .B(n_20380),
    .Y(n_26124));
 XOR2xp5_ASAP7_75t_SL g33136 (.A(n_20675),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_18),
    .Y(n_26125));
 XNOR2xp5_ASAP7_75t_SL g33137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .B(n_20789),
    .Y(n_26126));
 XOR2xp5_ASAP7_75t_SL g33138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_90),
    .Y(n_26127));
 OR2x2_ASAP7_75t_SL g33139 (.A(n_20927),
    .B(n_20926),
    .Y(n_26128));
 XNOR2x1_ASAP7_75t_SL g33140 (.B(n_21007),
    .Y(n_26129),
    .A(n_21004));
 XOR2x2_ASAP7_75t_SL g33141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_128),
    .Y(n_26130));
 XOR2xp5_ASAP7_75t_SL g33142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_164),
    .B(n_12948),
    .Y(n_26131));
 XOR2xp5_ASAP7_75t_SL g33143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .B(n_21131),
    .Y(n_26132));
 XNOR2x1_ASAP7_75t_SL g33144 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_627),
    .Y(n_26133),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_659));
 XNOR2xp5_ASAP7_75t_SL g33145 (.A(n_26000),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_9),
    .Y(n_26134));
 XOR2xp5_ASAP7_75t_SL g33146 (.A(n_8115),
    .B(n_8107),
    .Y(n_26135));
 XOR2xp5_ASAP7_75t_SL g33148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_113),
    .B(n_21454),
    .Y(n_26137));
 XNOR2xp5_ASAP7_75t_SL g33149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_118),
    .B(n_21467),
    .Y(n_26138));
 XOR2xp5_ASAP7_75t_SL g33150 (.A(n_9156),
    .B(n_9155),
    .Y(n_26139));
 XNOR2x1_ASAP7_75t_SL g33151 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_35),
    .Y(n_26140),
    .A(n_21606));
 XOR2xp5_ASAP7_75t_SL g33152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_89),
    .Y(n_26141));
 XOR2xp5_ASAP7_75t_SL g33153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_587),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_683),
    .Y(n_26142));
 XOR2xp5_ASAP7_75t_SL g33154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_36),
    .Y(n_26143));
 AND2x2_ASAP7_75t_SL g33155 (.A(n_25833),
    .B(n_23931),
    .Y(n_26144));
 XNOR2xp5_ASAP7_75t_SL g33156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_40),
    .Y(n_26145));
 XOR2xp5_ASAP7_75t_SL g33157 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_13),
    .Y(n_26146));
 XNOR2xp5_ASAP7_75t_SL g33158 (.A(n_7239),
    .B(n_17978),
    .Y(n_26147));
 XNOR2xp5_ASAP7_75t_SL g33159 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_79),
    .Y(n_26148));
 XOR2xp5_ASAP7_75t_SL g33160 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_183),
    .B(n_11194),
    .Y(n_26149));
 XNOR2xp5_ASAP7_75t_SL g33161 (.A(n_11289),
    .B(n_22167),
    .Y(n_26150));
 XNOR2xp5_ASAP7_75t_SL g33162 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_31),
    .Y(n_26151));
 XNOR2xp5_ASAP7_75t_SL g33163 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_111),
    .Y(n_26152));
 XOR2xp5_ASAP7_75t_SL g33164 (.A(n_13418),
    .B(n_9079),
    .Y(n_26153));
 XOR2xp5_ASAP7_75t_SL g33170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_153),
    .Y(n_26159));
 OR2x2_ASAP7_75t_SL g33175 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_75),
    .Y(n_26164));
 OR2x2_ASAP7_75t_SL g33177 (.A(n_23079),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_180),
    .Y(n_26166));
 XOR2xp5_ASAP7_75t_SL g33178 (.A(n_19945),
    .B(n_23135),
    .Y(n_26167));
 XNOR2xp5_ASAP7_75t_SL g33179 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_150),
    .Y(n_26168));
 XOR2xp5_ASAP7_75t_SL g33180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_212),
    .B(n_23380),
    .Y(n_26169));
 XNOR2xp5_ASAP7_75t_SL g33181 (.A(n_23394),
    .B(n_10648),
    .Y(n_26170));
 XOR2xp5_ASAP7_75t_SL g33183 (.A(n_18720),
    .B(n_3806),
    .Y(n_26172));
 XNOR2xp5_ASAP7_75t_SL g33184 (.A(n_23569),
    .B(n_22962),
    .Y(n_26173));
 XNOR2x1_ASAP7_75t_SL g33185 (.B(n_11533),
    .Y(n_26174),
    .A(n_19719));
 XNOR2x2_ASAP7_75t_SL g33186 (.A(n_19607),
    .B(n_20210),
    .Y(n_26175));
 FAx1_ASAP7_75t_SL g33188 (.SN(n_26177),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_38),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_87),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_159),
    .CON(UNCONNECTED20));
 AO21x1_ASAP7_75t_SL g33189 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_142),
    .A2(n_13248),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_167),
    .Y(n_26178));
 FAx1_ASAP7_75t_SL g33190 (.SN(n_26179),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .CON(UNCONNECTED21));
 FAx1_ASAP7_75t_SL g33191 (.SN(n_26180),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_573),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_n_701),
    .CON(UNCONNECTED22));
 FAx1_ASAP7_75t_SL g33192 (.SN(n_26181),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_767),
    .B(n_19057),
    .CI(n_19058),
    .CON(UNCONNECTED23));
 FAx1_ASAP7_75t_SL g33194 (.SN(n_26183),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_38),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_87),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_159),
    .CON(UNCONNECTED24));
 FAx1_ASAP7_75t_SL g33195 (.SN(n_26184),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_96),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_159),
    .CON(UNCONNECTED25));
 FAx1_ASAP7_75t_SL g33197 (.SN(n_26186),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_573),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_n_701),
    .CON(UNCONNECTED26));
 FAx1_ASAP7_75t_SL g33198 (.SN(n_26187),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_43),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_145),
    .CON(UNCONNECTED27));
 AOI21xp33_ASAP7_75t_SL g332 (.A1(n_11812),
    .A2(n_13521),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_276),
    .Y(n_14020));
 MAJIxp5_ASAP7_75t_SL g33200 (.A(n_2592),
    .B(n_8773),
    .C(n_25597),
    .Y(n_26189));
 FAx1_ASAP7_75t_SL g33201 (.SN(n_26190),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_573),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_n_701),
    .CON(UNCONNECTED28));
 FAx1_ASAP7_75t_SL g33202 (.SN(n_26191),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_43),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_145),
    .CON(UNCONNECTED29));
 OAI21xp33_ASAP7_75t_SL g33204 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_209),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_175),
    .B(n_19542),
    .Y(n_26193));
 FAx1_ASAP7_75t_SL g33205 (.SN(n_26194),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_38),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_87),
    .CI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_159),
    .CON(UNCONNECTED30));
 AOI22xp5_ASAP7_75t_SL g33207 (.A1(n_22162),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_76),
    .B1(n_22157),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_75),
    .Y(n_26196));
 MAJIxp5_ASAP7_75t_SL g33211 (.A(n_19913),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_17),
    .Y(n_26200));
 MAJIxp5_ASAP7_75t_SL g33213 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_673),
    .B(n_12550),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_737),
    .Y(n_26202));
 XNOR2xp5_ASAP7_75t_SL g33218 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_123),
    .Y(n_26207));
 MAJIxp5_ASAP7_75t_SL g33219 (.A(n_22841),
    .B(n_9709),
    .C(n_9711),
    .Y(n_26208));
 AOI31xp33_ASAP7_75t_SL g33221 (.A1(n_10677),
    .A2(n_10676),
    .A3(n_19194),
    .B(n_19279),
    .Y(n_26210));
 MAJIxp5_ASAP7_75t_SL g33223 (.A(n_12414),
    .B(n_12412),
    .C(n_12411),
    .Y(n_26212));
 XNOR2xp5_ASAP7_75t_SL g33224 (.A(n_11070),
    .B(n_25980),
    .Y(n_26213));
 MAJIxp5_ASAP7_75t_SL g33225 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_42),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_88),
    .Y(n_26214));
 AOI22xp5_ASAP7_75t_SL g33226 (.A1(n_21858),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_52),
    .B1(n_21857),
    .B2(n_21856),
    .Y(n_26215));
 MAJIxp5_ASAP7_75t_SL g33227 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_119),
    .Y(n_26216));
 XNOR2xp5_ASAP7_75t_SL g33229 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_51),
    .B(n_25988),
    .Y(n_26218));
 XNOR2xp5_ASAP7_75t_SL g33232 (.A(n_25989),
    .B(n_20236),
    .Y(n_26221));
 MAJx2_ASAP7_75t_SL g33233 (.A(n_23168),
    .B(n_23165),
    .C(n_20405),
    .Y(n_26222));
 MAJx2_ASAP7_75t_SL g33235 (.A(n_20379),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_100),
    .C(n_11270),
    .Y(n_26224));
 OAI21xp5_ASAP7_75t_SL g33237 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_65),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_167),
    .B(n_20825),
    .Y(n_26226));
 MAJIxp5_ASAP7_75t_SL g33238 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_22),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_113),
    .C(n_19796),
    .Y(n_26227));
 A2O1A1Ixp33_ASAP7_75t_SL g33239 (.A1(n_22634),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_71),
    .B(n_6614),
    .C(n_21023),
    .Y(n_26228));
 MAJx2_ASAP7_75t_SL g33242 (.A(n_21598),
    .B(n_21600),
    .C(n_13435),
    .Y(n_26231));
 MAJIxp5_ASAP7_75t_SL g33246 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_238),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_26),
    .C(n_4956),
    .Y(n_26235));
 INVx1_ASAP7_75t_SL g33247 (.A(n_26236),
    .Y(n_26237));
 A2O1A1Ixp33_ASAP7_75t_SL g33248 (.A1(n_22141),
    .A2(n_22142),
    .B(n_22143),
    .C(n_18767),
    .Y(n_26236));
 XNOR2xp5_ASAP7_75t_SL g33249 (.A(n_25987),
    .B(n_23228),
    .Y(n_26238));
 A2O1A1Ixp33_ASAP7_75t_SL g33250 (.A1(n_19531),
    .A2(n_20682),
    .B(n_20684),
    .C(n_12748),
    .Y(n_26239));
 XNOR2xp5_ASAP7_75t_SL g33252 (.A(n_20083),
    .B(n_25977),
    .Y(n_26241));
 OAI21xp5_ASAP7_75t_SL g33253 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_83),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_23),
    .B(n_22460),
    .Y(n_26242));
 XNOR2xp5_ASAP7_75t_SL g33254 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_133),
    .B(n_25992),
    .Y(n_26243));
 OAI211xp5_ASAP7_75t_SL g33255 (.A1(n_15561),
    .A2(n_13629),
    .B(n_9866),
    .C(n_22787),
    .Y(n_26244));
 NAND3xp33_ASAP7_75t_SL g33256 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_225),
    .B(n_24102),
    .C(n_22983),
    .Y(n_26245));
 OA22x2_ASAP7_75t_SL g33258 (.A1(n_23404),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_113),
    .B1(n_19682),
    .B2(n_26005),
    .Y(n_26247));
 A2O1A1Ixp33_ASAP7_75t_SL g33260 (.A1(n_2591),
    .A2(n_24208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_298),
    .C(n_24210),
    .Y(n_26249));
 OA22x2_ASAP7_75t_SL g33261 (.A1(n_23772),
    .A2(n_7577),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_174),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_185),
    .Y(n_26250));
 AOI21xp5_ASAP7_75t_SL g33262 (.A1(n_8178),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_217),
    .B(n_26251),
    .Y(n_26252));
 OAI21xp5_ASAP7_75t_SL g33263 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_193),
    .B(n_7595),
    .Y(n_26251));
 XOR2xp5_ASAP7_75t_SL g33266 (.A(n_26255),
    .B(n_17078),
    .Y(n_26256));
 AO21x1_ASAP7_75t_SL g33267 (.A1(n_8800),
    .A2(n_8802),
    .B(n_17443),
    .Y(n_26255));
 NAND2xp5_ASAP7_75t_SL g33268 (.A(n_26257),
    .B(n_2180),
    .Y(n_26258));
 XOR2xp5_ASAP7_75t_SL g33269 (.A(n_22081),
    .B(n_5724),
    .Y(n_26257));
 NAND2xp5_ASAP7_75t_SL g333 (.A(n_11812),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_310),
    .Y(n_14019));
 NAND2xp5_ASAP7_75t_SL g334 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_265),
    .Y(n_14017));
 INVx1_ASAP7_75t_SL g336 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_131),
    .Y(n_20951));
 AOI22xp5_ASAP7_75t_SL g337 (.A1(n_8105),
    .A2(n_8109),
    .B1(n_8108),
    .B2(n_22604),
    .Y(n_8115));
 MAJx2_ASAP7_75t_SL g338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_89),
    .C(n_17245),
    .Y(n_8107));
 INVx1_ASAP7_75t_SL g339 (.A(n_8108),
    .Y(n_8109));
 XNOR2xp5_ASAP7_75t_SL g34 (.A(n_20214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_31),
    .Y(n_20215));
 XNOR2xp5_ASAP7_75t_SL g340 (.A(n_17250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_128),
    .Y(n_8108));
 XNOR2xp5_ASAP7_75t_SL g342 (.A(n_19273),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_247),
    .Y(n_21840));
 XNOR2xp5_ASAP7_75t_SL g343 (.A(n_8104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_141),
    .Y(n_8105));
 INVx1_ASAP7_75t_SL g344 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_0),
    .Y(n_8104));
 AND2x2_ASAP7_75t_SL g345 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_249),
    .Y(n_21828));
 XNOR2xp5_ASAP7_75t_SL g346 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_272),
    .B(n_11032),
    .Y(n_11033));
 MAJx2_ASAP7_75t_SL g347 (.A(n_9525),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_210),
    .C(n_11169),
    .Y(n_12652));
 AND2x2_ASAP7_75t_SL g348 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_236),
    .B(n_11388),
    .Y(n_9776));
 NOR2xp33_ASAP7_75t_SL g349 (.A(n_14061),
    .B(n_14059),
    .Y(n_21850));
 NOR2x1_ASAP7_75t_SL g350 (.A(n_11521),
    .B(n_19912),
    .Y(n_7618));
 NAND2xp5_ASAP7_75t_SL g351 (.A(n_19912),
    .B(n_11521),
    .Y(n_7619));
 MAJIxp5_ASAP7_75t_SL g354 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_267),
    .B(n_7370),
    .C(n_4072),
    .Y(n_7371));
 OAI21xp5_ASAP7_75t_SL g355 (.A1(n_7378),
    .A2(n_20783),
    .B(n_20784),
    .Y(n_7379));
 OAI22xp5_ASAP7_75t_SL g358 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_49),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_40),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_48),
    .B2(n_13498),
    .Y(n_13499));
 XOR2xp5_ASAP7_75t_SL g359 (.A(n_20931),
    .B(n_20935),
    .Y(n_20936));
 NAND2xp5_ASAP7_75t_SL g360 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(n_16753),
    .Y(n_13495));
 MAJx2_ASAP7_75t_SL g362 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_92),
    .B(n_13797),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_78),
    .Y(n_20934));
 XNOR2xp5_ASAP7_75t_SL g363 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_61),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_1),
    .Y(n_20931));
 NAND2xp5_ASAP7_75t_SL g364 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(n_20932),
    .Y(n_20933));
 XOR2xp5_ASAP7_75t_SL g365 (.A(n_19769),
    .B(n_26214),
    .Y(n_19773));
 INVx1_ASAP7_75t_SL g366 (.A(n_19768),
    .Y(n_19769));
 MAJIxp5_ASAP7_75t_SL g367 (.A(n_19563),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_93),
    .C(n_15163),
    .Y(n_19768));
 XNOR2xp5_ASAP7_75t_SL g371 (.A(n_7222),
    .B(n_7212),
    .Y(n_7223));
 OAI21xp33_ASAP7_75t_SL g372 (.A1(n_5323),
    .A2(n_20066),
    .B(n_24181),
    .Y(n_20071));
 OAI22xp5_ASAP7_75t_SL g373 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .A2(n_6251),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .B2(n_15626),
    .Y(n_24207));
 XNOR2x1_ASAP7_75t_SL g374 (.B(n_6452),
    .Y(n_6453),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_26));
 XOR2xp5_ASAP7_75t_SL g375 (.A(n_23174),
    .B(n_23175),
    .Y(n_2588));
 MAJx2_ASAP7_75t_SL g376 (.A(n_23988),
    .B(n_23985),
    .C(n_18862),
    .Y(n_6452));
 OAI21xp5_ASAP7_75t_SL g377 (.A1(n_20783),
    .A2(n_19530),
    .B(n_20784),
    .Y(n_24200));
 AOI21x1_ASAP7_75t_SL g378 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_309),
    .A2(n_23123),
    .B(n_20393),
    .Y(n_23124));
 AOI21x1_ASAP7_75t_SL g379 (.A1(n_23123),
    .A2(n_21471),
    .B(n_20650),
    .Y(n_23125));
 AOI221xp5_ASAP7_75t_SL g38 (.A1(n_19697),
    .A2(n_19698),
    .B1(n_21045),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_115),
    .C(n_19699),
    .Y(n_19700));
 AOI321xp33_ASAP7_75t_SL g380 (.A1(n_20649),
    .A2(n_23123),
    .A3(n_20646),
    .B1(n_20650),
    .B2(n_20651),
    .C(n_20654),
    .Y(n_23128));
 INVx1_ASAP7_75t_SL g381 (.A(n_18862),
    .Y(n_6456));
 INVx2_ASAP7_75t_SL g382 (.A(n_23121),
    .Y(n_23123));
 AOI21x1_ASAP7_75t_SL g383 (.A1(n_23118),
    .A2(n_23119),
    .B(n_23120),
    .Y(n_23121));
 XNOR2xp5_ASAP7_75t_SL g384 (.A(n_23130),
    .B(n_23131),
    .Y(n_23132));
 XNOR2xp5_ASAP7_75t_SL g385 (.A(n_8581),
    .B(n_7537),
    .Y(n_7542));
 MAJIxp5_ASAP7_75t_SL g386 (.A(n_20139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_29),
    .C(n_3364),
    .Y(n_7534));
 INVxp67_ASAP7_75t_SL g387 (.A(n_8581),
    .Y(n_7536));
 NOR2xp33_ASAP7_75t_SL g388 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_247),
    .Y(n_8166));
 INVxp67_ASAP7_75t_SL g389 (.A(n_7537),
    .Y(n_7538));
 AOI221xp5_ASAP7_75t_SL g39 (.A1(n_13483),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_212),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_221),
    .B2(n_20114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_230),
    .Y(n_13487));
 XNOR2xp5_ASAP7_75t_SL g390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_192),
    .B(n_23197),
    .Y(n_7537));
 XOR2x2_ASAP7_75t_SL g391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_135),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_114),
    .Y(n_9632));
 OAI21xp5_ASAP7_75t_SL g392 (.A1(n_20902),
    .A2(n_20903),
    .B(n_20904),
    .Y(n_20905));
 A2O1A1Ixp33_ASAP7_75t_SL g393 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .B(n_12698),
    .C(n_12700),
    .Y(n_12701));
 MAJIxp5_ASAP7_75t_SL g394 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_325),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(n_12700));
 OAI21xp5_ASAP7_75t_SL g395 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(n_12707));
 NAND2xp5_ASAP7_75t_SL g396 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .Y(n_12696));
 NOR2xp33_ASAP7_75t_SL g397 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .Y(n_12698));
 NAND2xp5_ASAP7_75t_SL g398 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .Y(n_12697));
 INVx1_ASAP7_75t_SL g399 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .Y(n_12702));
 AOI21xp33_ASAP7_75t_SL g40 (.A1(n_13687),
    .A2(n_5456),
    .B(n_16458),
    .Y(n_5457));
 INVx1_ASAP7_75t_SL g400 (.A(n_5994),
    .Y(n_5996));
 NAND2xp5_ASAP7_75t_SL g401 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[17]),
    .B(n_17870),
    .Y(n_5994));
 MAJIxp5_ASAP7_75t_SL g403 (.A(n_23682),
    .B(n_23683),
    .C(n_23684),
    .Y(n_23685));
 XNOR2xp5_ASAP7_75t_SL g405 (.A(n_10745),
    .B(n_13054),
    .Y(n_23684));
 INVx1_ASAP7_75t_SL g406 (.A(n_18933),
    .Y(n_6295));
 AOI21xp5_ASAP7_75t_SL g407 (.A1(n_22790),
    .A2(n_22791),
    .B(n_22792),
    .Y(n_22793));
 XNOR2xp5_ASAP7_75t_SL g409 (.A(n_13644),
    .B(n_13650),
    .Y(n_13651));
 XNOR2x1_ASAP7_75t_SL g41 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_221),
    .Y(n_13480),
    .A(n_20114));
 NAND2xp5_ASAP7_75t_SL g410 (.A(n_13652),
    .B(n_13649),
    .Y(n_13654));
 INVxp67_ASAP7_75t_SRAM g412 (.A(n_6979),
    .Y(n_6989));
 NOR2xp33_ASAP7_75t_SL g413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_238),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_241),
    .Y(n_6979));
 NAND2xp5_ASAP7_75t_SL g414 (.A(n_7099),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_310),
    .Y(n_7100));
 NAND2xp5_ASAP7_75t_SL g415 (.A(n_6985),
    .B(n_6986),
    .Y(n_6987));
 NOR2xp33_ASAP7_75t_SL g416 (.A(n_6368),
    .B(n_9404),
    .Y(n_6978));
 OAI21xp5_ASAP7_75t_SL g418 (.A1(n_20160),
    .A2(n_5371),
    .B(n_5873),
    .Y(n_5874));
 NAND2xp5_ASAP7_75t_SL g419 (.A(n_20158),
    .B(n_5872),
    .Y(n_5873));
 OAI21xp5_ASAP7_75t_SL g42 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_65),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_189),
    .Y(n_19523));
 A2O1A1Ixp33_ASAP7_75t_SL g4226 (.A1(n_23059),
    .A2(n_23060),
    .B(n_23064),
    .C(n_23065),
    .Y(n_23066));
 OAI21xp5_ASAP7_75t_SL g4227 (.A1(n_23067),
    .A2(n_23069),
    .B(n_23296),
    .Y(n_23070));
 AOI21xp5_ASAP7_75t_SL g4228 (.A1(n_14689),
    .A2(n_23054),
    .B(n_23057),
    .Y(n_23058));
 OAI21xp5_ASAP7_75t_SL g4229 (.A1(n_23041),
    .A2(n_23047),
    .B(n_23051),
    .Y(n_23052));
 OAI31xp33_ASAP7_75t_SL g4230 (.A1(n_23046),
    .A2(n_23043),
    .A3(n_23053),
    .B(n_23056),
    .Y(n_23057));
 NOR2xp33_ASAP7_75t_SL g4231 (.A(n_23043),
    .B(n_23046),
    .Y(n_23047));
 NAND2xp5_ASAP7_75t_SL g4232 (.A(n_23039),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_295),
    .Y(n_23041));
 NAND3x1_ASAP7_75t_L g4233 (.A(n_23296),
    .B(n_23062),
    .C(n_23063),
    .Y(n_23064));
 AOI21xp33_ASAP7_75t_SL g4234 (.A1(n_23037),
    .A2(n_23049),
    .B(n_23038),
    .Y(n_23056));
 AO21x1_ASAP7_75t_SL g4235 (.A1(n_23049),
    .A2(n_10181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_274),
    .Y(n_23065));
 AOI22xp5_ASAP7_75t_SL g4236 (.A1(n_23068),
    .A2(n_23042),
    .B1(n_9392),
    .B2(n_22956),
    .Y(n_23069));
 AOI21xp5_ASAP7_75t_SL g4237 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_295),
    .B(n_23050),
    .Y(n_23051));
 OR2x2_ASAP7_75t_SL g4239 (.A(n_25983),
    .B(n_23045),
    .Y(n_23046));
 OAI21xp5_ASAP7_75t_SL g424 (.A1(n_5369),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_468),
    .B(n_5372),
    .Y(n_5872));
 NOR2xp33_ASAP7_75t_SL g4240 (.A(n_23049),
    .B(n_20324),
    .Y(n_23050));
 NOR2xp33_ASAP7_75t_SL g4241 (.A(n_23037),
    .B(n_23038),
    .Y(n_23039));
 NOR2xp33_ASAP7_75t_SL g4242 (.A(n_23053),
    .B(n_23045),
    .Y(n_23054));
 NOR2xp33_ASAP7_75t_SL g4243 (.A(n_23038),
    .B(n_23053),
    .Y(n_23072));
 NOR2xp33_ASAP7_75t_SRAM g4244 (.A(n_23045),
    .B(n_23037),
    .Y(n_23071));
 INVxp67_ASAP7_75t_SL g4245 (.A(n_23038),
    .Y(n_23063));
 AND2x2_ASAP7_75t_SL g4246 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_270),
    .Y(n_23038));
 INVx2_ASAP7_75t_SL g4247 (.A(n_23042),
    .Y(n_23043));
 INVxp67_ASAP7_75t_SL g4248 (.A(n_23043),
    .Y(n_23059));
 OR2x2_ASAP7_75t_SL g4250 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_289),
    .Y(n_23042));
 HB1xp67_ASAP7_75t_SL g4251 (.A(n_23045),
    .Y(n_23067));
 NOR2x1_ASAP7_75t_SL g4252 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_266),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_284),
    .Y(n_23045));
 NOR2x1_ASAP7_75t_SL g4253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_268),
    .Y(n_23053));
 OR2x2_ASAP7_75t_SL g4254 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_268),
    .Y(n_23049));
 AND2x2_ASAP7_75t_SL g4256 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_284),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_266),
    .Y(n_23037));
 NOR2xp67_ASAP7_75t_L g426 (.A(n_5869),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_447),
    .Y(n_5870));
 INVx1_ASAP7_75t_SL g4260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_274),
    .Y(n_23062));
 INVxp33_ASAP7_75t_SRAM g427 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_447),
    .Y(n_5867));
 INVx1_ASAP7_75t_SL g428 (.A(n_5372),
    .Y(n_5869));
 INVx2_ASAP7_75t_SL g431 (.A(n_5953),
    .Y(n_5954));
 XNOR2x1_ASAP7_75t_SL g433 (.B(n_26125),
    .Y(n_5953),
    .A(n_5951));
 INVxp67_ASAP7_75t_SL g434 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_63),
    .Y(n_5951));
 MAJIxp5_ASAP7_75t_SL g436 (.A(n_19670),
    .B(n_19674),
    .C(n_19676),
    .Y(n_19677));
 NAND2x1_ASAP7_75t_SL g437 (.A(n_7777),
    .B(n_13361),
    .Y(n_7778));
 OR2x2_ASAP7_75t_SL g438 (.A(n_6830),
    .B(n_13361),
    .Y(n_7780));
 NOR2xp67_ASAP7_75t_L g439 (.A(n_6830),
    .B(n_13361),
    .Y(n_7784));
 NAND2xp5_ASAP7_75t_L g44 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_290),
    .B(n_11858),
    .Y(n_19732));
 XNOR2xp5_ASAP7_75t_SL g440 (.A(n_14116),
    .B(n_19014),
    .Y(n_14117));
 MAJIxp5_ASAP7_75t_SL g441 (.A(n_13416),
    .B(n_8241),
    .C(n_14115),
    .Y(n_14118));
 INVxp67_ASAP7_75t_SL g442 (.A(n_14115),
    .Y(n_14116));
 XNOR2xp5_ASAP7_75t_SL g443 (.A(n_9065),
    .B(n_18875),
    .Y(n_14115));
 INVx1_ASAP7_75t_SL g446 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_80),
    .Y(n_19673));
 AOI22x1_ASAP7_75t_SL g448 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_n_709),
    .A2(n_6325),
    .B1(n_6326),
    .B2(n_19555),
    .Y(n_6327));
 INVxp67_ASAP7_75t_SL g449 (.A(n_22437),
    .Y(n_6331));
 AND2x2_ASAP7_75t_SL g45 (.A(n_2161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_620),
    .Y(n_23668));
 HB1xp67_ASAP7_75t_SL g451 (.A(n_9354),
    .Y(n_6329));
 OR2x2_ASAP7_75t_SL g453 (.A(n_19554),
    .B(n_19555),
    .Y(n_6325));
 HB1xp67_ASAP7_75t_SL g455 (.A(n_20945),
    .Y(n_6324));
 XNOR2x1_ASAP7_75t_SL g46 (.B(n_12754),
    .Y(n_8689),
    .A(n_8688));
 XNOR2xp5_ASAP7_75t_SL g460 (.A(n_6348),
    .B(n_6350),
    .Y(n_6351));
 OA21x2_ASAP7_75t_SL g461 (.A1(n_19380),
    .A2(n_25605),
    .B(n_12680),
    .Y(n_13605));
 OAI22xp5_ASAP7_75t_SL g463 (.A1(n_6342),
    .A2(n_6339),
    .B1(n_6341),
    .B2(n_6349),
    .Y(n_6350));
 OAI21x1_ASAP7_75t_SL g465 (.A1(n_13600),
    .A2(n_25606),
    .B(n_13602),
    .Y(n_13603));
 INVx1_ASAP7_75t_SL g466 (.A(n_6341),
    .Y(n_6342));
 MAJIxp5_ASAP7_75t_SL g467 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_751),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_687),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_591),
    .Y(n_6341));
 INVx1_ASAP7_75t_SL g468 (.A(n_6339),
    .Y(n_6349));
 XNOR2x1_ASAP7_75t_SL g469 (.B(n_16000),
    .Y(n_6339),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_717));
 XNOR2xp5_ASAP7_75t_SL g47 (.A(n_13413),
    .B(n_13415),
    .Y(n_13416));
 INVxp67_ASAP7_75t_SL g470 (.A(n_6343),
    .Y(n_6348));
 XNOR2xp5_ASAP7_75t_SL g471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_17),
    .B(n_17553),
    .Y(n_6343));
 INVx1_ASAP7_75t_SL g472 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_57),
    .Y(n_8324));
 INVxp67_ASAP7_75t_SL g473 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_62),
    .Y(n_8325));
 INVxp67_ASAP7_75t_SL g474 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273),
    .Y(n_13602));
 AOI21xp5_ASAP7_75t_SL g479 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_217),
    .A2(n_20326),
    .B(n_19232),
    .Y(n_20327));
 XOR2xp5_ASAP7_75t_SL g48 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_779),
    .B(n_21697),
    .Y(n_13415));
 XNOR2xp5_ASAP7_75t_SL g480 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_223),
    .B(n_20326),
    .Y(n_20328));
 OAI21xp5_ASAP7_75t_SL g481 (.A1(n_20322),
    .A2(n_10180),
    .B(n_23052),
    .Y(n_20326));
 NAND2xp5_ASAP7_75t_SL g482 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_26),
    .Y(n_8323));
 NAND2xp5_ASAP7_75t_SL g483 (.A(n_23054),
    .B(n_20321),
    .Y(n_20322));
 INVx1_ASAP7_75t_SL g484 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_286),
    .Y(n_20321));
 INVx1_ASAP7_75t_SL g485 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_295),
    .Y(n_20324));
 INVx1_ASAP7_75t_SL g49 (.A(n_21697),
    .Y(n_13417));
 AOI21x1_ASAP7_75t_SL g50 (.A1(n_22013),
    .A2(n_25833),
    .B(n_5420),
    .Y(n_5421));
 MAJIxp5_ASAP7_75t_SL g505 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_115),
    .B(n_14820),
    .C(n_26089),
    .Y(n_3611));
 NAND2xp5_ASAP7_75t_SL g509 (.A(n_18799),
    .B(n_7162),
    .Y(n_7166));
 INVxp67_ASAP7_75t_SL g51 (.A(n_20624),
    .Y(n_5420));
 AND2x2_ASAP7_75t_SL g512 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .Y(n_7162));
 NAND2xp5_ASAP7_75t_SL g513 (.A(n_21659),
    .B(n_21661),
    .Y(n_21662));
 AOI21xp33_ASAP7_75t_SL g514 (.A1(n_21656),
    .A2(n_21657),
    .B(n_21658),
    .Y(n_21659));
 XNOR2xp5_ASAP7_75t_SL g515 (.A(n_18712),
    .B(n_21655),
    .Y(n_21663));
 OAI21xp33_ASAP7_75t_SL g516 (.A1(n_21655),
    .A2(n_21222),
    .B(n_21660),
    .Y(n_21661));
 INVx1_ASAP7_75t_SL g517 (.A(n_21655),
    .Y(n_21656));
 AOI21x1_ASAP7_75t_SL g518 (.A1(n_9037),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_319),
    .B(n_11077),
    .Y(n_21655));
 NOR2xp33_ASAP7_75t_SL g519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_280),
    .B(n_21222),
    .Y(n_21657));
 INVxp33_ASAP7_75t_SL g52 (.A(n_23578),
    .Y(n_23581));
 AND2x2_ASAP7_75t_SL g520 (.A(n_21224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_280),
    .Y(n_21660));
 NOR2xp33_ASAP7_75t_SL g521 (.A(n_21224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_280),
    .Y(n_21658));
 XNOR2xp5_ASAP7_75t_SL g524 (.A(n_12386),
    .B(n_12390),
    .Y(n_12391));
 OAI211xp5_ASAP7_75t_SL g525 (.A1(n_12380),
    .A2(n_12376),
    .B(n_12381),
    .C(n_12385),
    .Y(n_12386));
 OAI21xp5_ASAP7_75t_SL g526 (.A1(n_12387),
    .A2(n_12388),
    .B(n_12389),
    .Y(n_12390));
 NAND2xp5_ASAP7_75t_SL g527 (.A(n_12387),
    .B(n_12388),
    .Y(n_12389));
 NAND3xp33_ASAP7_75t_SL g528 (.A(n_18753),
    .B(n_12379),
    .C(n_9384),
    .Y(n_12381));
 AOI21xp5_ASAP7_75t_SL g529 (.A1(n_12379),
    .A2(n_9385),
    .B(n_12384),
    .Y(n_12385));
 AND2x2_ASAP7_75t_SL g53 (.A(n_19370),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_708),
    .Y(n_21052));
 OAI21x1_ASAP7_75t_SL g530 (.A1(n_12392),
    .A2(n_12376),
    .B(n_12393),
    .Y(n_12394));
 NAND2xp33_ASAP7_75t_SL g531 (.A(n_10427),
    .B(n_12379),
    .Y(n_12380));
 OAI22xp5_ASAP7_75t_SL g532 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_3),
    .A2(n_6794),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_140),
    .B2(n_6795),
    .Y(n_6796));
 XNOR2xp5_ASAP7_75t_SL g533 (.A(n_6797),
    .B(n_6798),
    .Y(n_6799));
 INVx1_ASAP7_75t_SL g534 (.A(n_6794),
    .Y(n_6795));
 MAJIxp5_ASAP7_75t_SL g535 (.A(n_6789),
    .B(n_6791),
    .C(n_6793),
    .Y(n_6794));
 XOR2xp5_ASAP7_75t_SL g536 (.A(n_13726),
    .B(n_6792),
    .Y(n_6798));
 NOR2xp33_ASAP7_75t_SL g537 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_46),
    .B(n_12120),
    .Y(n_6789));
 NOR2xp33_ASAP7_75t_SL g538 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_46),
    .B(n_12120),
    .Y(n_6797));
 INVx1_ASAP7_75t_SL g539 (.A(n_6792),
    .Y(n_6793));
 AOI22xp5_ASAP7_75t_SL g54 (.A1(n_13788),
    .A2(n_22069),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_101),
    .B2(n_9341),
    .Y(n_22071));
 NAND2xp5_ASAP7_75t_SL g540 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .Y(n_6792));
 INVx1_ASAP7_75t_SL g541 (.A(n_13726),
    .Y(n_6791));
 NAND2xp5_ASAP7_75t_SL g543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_174),
    .Y(n_12383));
 NAND2x1_ASAP7_75t_SL g545 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_224),
    .Y(n_12382));
 XNOR2x1_ASAP7_75t_SL g55 (.B(n_9141),
    .Y(n_9142),
    .A(n_18925));
 OAI22xp5_ASAP7_75t_SL g551 (.A1(n_19785),
    .A2(n_23393),
    .B1(n_20943),
    .B2(n_23389),
    .Y(n_20945));
 INVx1_ASAP7_75t_SL g554 (.A(n_20943),
    .Y(n_19785));
 XNOR2x2_ASAP7_75t_SL g555 (.A(n_11630),
    .B(n_16367),
    .Y(n_11638));
 MAJIxp5_ASAP7_75t_SL g556 (.A(n_11630),
    .B(n_16365),
    .C(n_13181),
    .Y(n_11644));
 NAND2xp5_ASAP7_75t_SL g557 (.A(n_2176),
    .B(n_18774),
    .Y(n_20938));
 MAJIxp5_ASAP7_75t_SL g559 (.A(n_21351),
    .B(n_7754),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_180),
    .Y(n_11630));
 XNOR2x2_ASAP7_75t_SL g56 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_65),
    .B(n_18832),
    .Y(n_5398));
 XOR2xp5_ASAP7_75t_SL g560 (.A(n_14742),
    .B(n_19033),
    .Y(n_14746));
 INVxp67_ASAP7_75t_SRAM g561 (.A(n_10506),
    .Y(n_20946));
 INVx1_ASAP7_75t_SL g563 (.A(n_18774),
    .Y(n_20939));
 INVx1_ASAP7_75t_SL g564 (.A(n_14902),
    .Y(n_14910));
 XNOR2x1_ASAP7_75t_SL g565 (.B(n_14748),
    .Y(n_14749),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_3));
 AND2x2_ASAP7_75t_SL g566 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_0),
    .Y(n_14742));
 OA21x2_ASAP7_75t_SL g567 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_229),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_228),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_231),
    .Y(n_14929));
 INVxp67_ASAP7_75t_SL g568 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_141),
    .Y(n_14739));
 NAND2xp5_ASAP7_75t_SL g57 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .B(n_19645),
    .Y(n_19446));
 INVxp67_ASAP7_75t_SL g571 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_73),
    .Y(n_14748));
 XOR2xp5_ASAP7_75t_SL g572 (.A(n_11121),
    .B(n_22260),
    .Y(n_22261));
 A2O1A1Ixp33_ASAP7_75t_SL g573 (.A1(n_12379),
    .A2(n_12394),
    .B(n_10320),
    .C(n_10321),
    .Y(n_10322));
 MAJx2_ASAP7_75t_SL g574 (.A(n_26128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_80),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_89),
    .Y(n_22257));
 OAI22xp33_ASAP7_75t_SL g575 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_264),
    .A2(n_12394),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_265),
    .B2(n_10318),
    .Y(n_10319));
 INVx1_ASAP7_75t_SL g576 (.A(n_22258),
    .Y(n_22259));
 XNOR2xp5_ASAP7_75t_SL g577 (.A(n_10905),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_128),
    .Y(n_22258));
 OR2x2_ASAP7_75t_SL g578 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_191),
    .B(n_12384),
    .Y(n_10320));
 OR2x2_ASAP7_75t_SL g579 (.A(n_12389),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_191),
    .Y(n_10321));
 INVxp67_ASAP7_75t_SL g58 (.A(n_19447),
    .Y(n_19448));
 NAND2x1_ASAP7_75t_SL g59 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_14987),
    .Y(n_19447));
 NAND2xp5_ASAP7_75t_SL g6 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .Y(n_9350));
 MAJIxp5_ASAP7_75t_SL g61 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_98),
    .B(n_19557),
    .C(n_19558),
    .Y(n_5536));
 OAI22xp5_ASAP7_75t_SL g62 (.A1(n_19567),
    .A2(n_19568),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_49),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_40),
    .Y(n_19570));
 AOI321xp33_ASAP7_75t_SL g633 (.A1(n_6727),
    .A2(n_11454),
    .A3(n_6733),
    .B1(n_16706),
    .B2(n_16705),
    .C(n_10177),
    .Y(n_8803));
 INVxp67_ASAP7_75t_SL g634 (.A(n_8801),
    .Y(n_8802));
 MAJIxp5_ASAP7_75t_SL g635 (.A(n_11453),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_320),
    .C(n_16705),
    .Y(n_8801));
 XNOR2xp5_ASAP7_75t_SL g637 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_349),
    .Y(n_8799));
 OAI22xp5_ASAP7_75t_SL g639 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_158),
    .A2(n_9123),
    .B1(n_9120),
    .B2(n_12252),
    .Y(n_11108));
 NAND2xp5_ASAP7_75t_SL g64 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .Y(n_19567));
 MAJx2_ASAP7_75t_SL g640 (.A(n_19826),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_17),
    .C(n_20770),
    .Y(n_14881));
 XOR2xp5_ASAP7_75t_SL g641 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_175),
    .B(n_5744),
    .Y(n_14880));
 OAI22xp5_ASAP7_75t_SL g644 (.A1(n_14439),
    .A2(n_3522),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_226),
    .B2(n_14442),
    .Y(n_14443));
 MAJIxp5_ASAP7_75t_SL g645 (.A(n_13359),
    .B(n_3521),
    .C(n_14444),
    .Y(n_14445));
 HB1xp67_ASAP7_75t_SL g646 (.A(n_14442),
    .Y(n_14444));
 MAJIxp5_ASAP7_75t_SL g647 (.A(n_14440),
    .B(n_14441),
    .C(n_14437),
    .Y(n_14442));
 MAJIxp5_ASAP7_75t_SL g648 (.A(n_14438),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_171),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_10),
    .Y(n_14439));
 MAJIxp5_ASAP7_75t_SL g65 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_95),
    .B(n_5548),
    .C(n_14704),
    .Y(n_5549));
 INVx1_ASAP7_75t_SL g652 (.A(n_6156),
    .Y(n_6157));
 AOI211x1_ASAP7_75t_SL g653 (.A1(n_6149),
    .A2(n_6150),
    .B(n_6153),
    .C(n_19128),
    .Y(n_6156));
 OAI21xp5_ASAP7_75t_SL g654 (.A1(n_6145),
    .A2(n_6147),
    .B(n_6152),
    .Y(n_6153));
 NAND2xp5_ASAP7_75t_SL g655 (.A(n_6147),
    .B(n_6151),
    .Y(n_6152));
 NOR2xp33_ASAP7_75t_SL g658 (.A(n_6144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_37),
    .Y(n_6151));
 NAND2xp5_ASAP7_75t_SL g66 (.A(n_24102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_305),
    .Y(n_24106));
 NOR2xp67_ASAP7_75t_SL g660 (.A(n_6144),
    .B(n_6148),
    .Y(n_6149));
 INVx1_ASAP7_75t_SL g663 (.A(n_6144),
    .Y(n_6145));
 AND2x2_ASAP7_75t_SL g664 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .B(n_3275),
    .Y(n_6144));
 INVx1_ASAP7_75t_SL g665 (.A(n_6147),
    .Y(n_6148));
 NAND2xp5_ASAP7_75t_SL g666 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_36),
    .Y(n_6147));
 INVxp67_ASAP7_75t_SL g667 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_84),
    .Y(n_6150));
 OAI22xp5_ASAP7_75t_SL g669 (.A1(n_8919),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_n_757),
    .B2(n_8926),
    .Y(n_8929));
 NOR2xp67_ASAP7_75t_SL g67 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_117),
    .Y(n_9375));
 INVx1_ASAP7_75t_SL g674 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .Y(n_8926));
 INVxp67_ASAP7_75t_SL g675 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_757),
    .Y(n_8919));
 XNOR2xp5_ASAP7_75t_SL g68 (.A(n_19601),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_36),
    .Y(n_19602));
 INVxp67_ASAP7_75t_SL g686 (.A(n_9501),
    .Y(n_9507));
 NOR2xp67_ASAP7_75t_SL g687 (.A(n_5793),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_243),
    .Y(n_9501));
 INVx1_ASAP7_75t_SL g688 (.A(n_9498),
    .Y(n_9506));
 MAJIxp5_ASAP7_75t_SL g69 (.A(n_5411),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_152),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_203),
    .Y(n_5412));
 AOI21xp5_ASAP7_75t_SL g690 (.A1(n_8623),
    .A2(n_8625),
    .B(n_8628),
    .Y(n_8629));
 NAND2xp5_ASAP7_75t_SL g691 (.A(n_8623),
    .B(n_8621),
    .Y(n_8624));
 NOR2xp67_ASAP7_75t_SL g693 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_241),
    .B(n_22819),
    .Y(n_8628));
 NAND2xp5_ASAP7_75t_SL g694 (.A(n_22819),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_241),
    .Y(n_8623));
 NOR2xp33_ASAP7_75t_SL g695 (.A(n_8626),
    .B(n_8637),
    .Y(n_8638));
 INVxp67_ASAP7_75t_SL g696 (.A(n_8626),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_241));
 MAJIxp5_ASAP7_75t_SL g697 (.A(n_7223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_167),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_7),
    .Y(n_8626));
 MAJx2_ASAP7_75t_SL g698 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_141),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_66),
    .Y(n_8660));
 INVx1_ASAP7_75t_SL g7 (.A(n_24230),
    .Y(n_24231));
 OAI22xp5_ASAP7_75t_SL g70 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_154),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_151),
    .B1(n_5409),
    .B2(n_5410),
    .Y(n_5411));
 AND2x2_ASAP7_75t_SL g700 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_179),
    .Y(n_8658));
 INVx1_ASAP7_75t_SL g702 (.A(n_8621),
    .Y(n_8639));
 NAND2xp5_ASAP7_75t_SL g703 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_243),
    .Y(n_8621));
 INVxp67_ASAP7_75t_SL g704 (.A(n_8625),
    .Y(n_8640));
 NOR2xp33_ASAP7_75t_SL g705 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_243),
    .Y(n_8625));
 HB1xp67_ASAP7_75t_SL g708 (.A(n_8069),
    .Y(n_8631));
 INVx1_ASAP7_75t_SL g71 (.A(n_13794),
    .Y(n_20217));
 OAI22x1_ASAP7_75t_SL g715 (.A1(n_12980),
    .A2(n_12985),
    .B1(n_12986),
    .B2(n_12987),
    .Y(n_12988));
 NOR2x1_ASAP7_75t_SL g716 (.A(n_12982),
    .B(n_12984),
    .Y(n_12985));
 AND3x1_ASAP7_75t_SL g717 (.A(n_12511),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_680),
    .C(n_12979),
    .Y(n_12980));
 INVxp67_ASAP7_75t_SL g718 (.A(n_6879),
    .Y(n_12982));
 AND3x1_ASAP7_75t_SL g719 (.A(n_9301),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .C(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[0]),
    .Y(n_12981));
 INVx1_ASAP7_75t_SL g72 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_154),
    .Y(n_5409));
 XNOR2xp5_ASAP7_75t_SL g720 (.A(n_18787),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_298),
    .Y(n_12984));
 AND2x2_ASAP7_75t_SL g723 (.A(n_2160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_680),
    .Y(n_12987));
 INVxp67_ASAP7_75t_SL g724 (.A(n_5986),
    .Y(n_5988));
 AOI21xp5_ASAP7_75t_SL g725 (.A1(n_5983),
    .A2(n_21644),
    .B(n_5985),
    .Y(n_5986));
 XNOR2x1_ASAP7_75t_SL g726 (.B(n_5980),
    .Y(n_5990),
    .A(n_5981));
 NOR2xp33_ASAP7_75t_SL g727 (.A(n_5980),
    .B(n_5982),
    .Y(n_5985));
 NAND2xp5_ASAP7_75t_SL g728 (.A(n_5980),
    .B(n_5982),
    .Y(n_5983));
 INVx2_ASAP7_75t_SL g729 (.A(n_21644),
    .Y(n_5991));
 XOR2xp5_ASAP7_75t_SL g73 (.A(n_21164),
    .B(n_21159),
    .Y(n_21160));
 OAI21x1_ASAP7_75t_SL g731 (.A1(n_18582),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_86),
    .Y(n_5980));
 XOR2x2_ASAP7_75t_SL g733 (.A(n_22002),
    .B(n_9794),
    .Y(n_5981));
 OAI22x1_ASAP7_75t_SL g74 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_101),
    .A2(n_11826),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_102),
    .B2(n_11827),
    .Y(n_11828));
 NOR3xp33_ASAP7_75t_SL g756 (.A(n_14894),
    .B(n_14896),
    .C(n_17870),
    .Y(n_14897));
 NOR2xp33_ASAP7_75t_SL g758 (.A(n_17870),
    .B(n_2850),
    .Y(n_14893));
 AOI21xp5_ASAP7_75t_SL g759 (.A1(n_16162),
    .A2(n_12778),
    .B(n_12779),
    .Y(n_12780));
 NOR2x1_ASAP7_75t_SL g761 (.A(n_12775),
    .B(n_12774),
    .Y(n_12779));
 MAJx2_ASAP7_75t_SL g762 (.A(n_2791),
    .B(n_18069),
    .C(n_8588),
    .Y(n_12775));
 XOR2x2_ASAP7_75t_SL g764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_349),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .Y(n_12774));
 NAND2xp5_ASAP7_75t_SL g765 (.A(n_11384),
    .B(n_10205),
    .Y(n_12778));
 HB1xp67_ASAP7_75t_SL g77 (.A(n_20103),
    .Y(n_20107));
 AOI21xp33_ASAP7_75t_SL g78 (.A1(n_14177),
    .A2(n_22307),
    .B(n_22308),
    .Y(n_22309));
 NAND2xp5_ASAP7_75t_L g8 (.A(n_3528),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .Y(n_21157));
 INVx1_ASAP7_75t_SL g80 (.A(n_13723),
    .Y(n_5602));
 NOR2xp33_ASAP7_75t_SL g82 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_246),
    .Y(n_20977));
 AOI21xp33_ASAP7_75t_SL g833 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_304),
    .A2(n_19281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_308),
    .Y(n_19282));
 INVxp67_ASAP7_75t_SL g836 (.A(n_19281),
    .Y(n_19283));
 OAI21x1_ASAP7_75t_SL g837 (.A1(n_19278),
    .A2(n_19279),
    .B(n_19280),
    .Y(n_19281));
 AOI21x1_ASAP7_75t_SL g838 (.A1(n_19275),
    .A2(n_19276),
    .B(n_19277),
    .Y(n_19278));
 NOR2xp33_ASAP7_75t_SL g839 (.A(n_19290),
    .B(n_19277),
    .Y(n_19291));
 XNOR2x1_ASAP7_75t_SL g84 (.B(n_5640),
    .Y(n_5641),
    .A(n_5639));
 INVxp67_ASAP7_75t_SL g841 (.A(n_19275),
    .Y(n_19290));
 OAI21xp5_ASAP7_75t_SL g842 (.A1(n_10588),
    .A2(n_11746),
    .B(n_19169),
    .Y(n_19275));
 INVxp33_ASAP7_75t_SRAM g843 (.A(n_19276),
    .Y(n_19288));
 AO21x1_ASAP7_75t_SL g844 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_250),
    .A2(n_13389),
    .B(n_13390),
    .Y(n_19276));
 AOI21xp5_ASAP7_75t_SL g845 (.A1(n_10677),
    .A2(n_10676),
    .B(n_19194),
    .Y(n_19279));
 NAND3xp33_ASAP7_75t_SL g846 (.A(n_10677),
    .B(n_10676),
    .C(n_19194),
    .Y(n_19280));
 NOR3xp33_ASAP7_75t_SL g848 (.A(n_10588),
    .B(n_19169),
    .C(n_11746),
    .Y(n_19277));
 XNOR2x1_ASAP7_75t_SL g85 (.B(n_5800),
    .Y(n_5640),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_779));
 AOI21xp5_ASAP7_75t_SL g852 (.A1(n_6190),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_290),
    .B(n_5544),
    .Y(n_8787));
 XOR2xp5_ASAP7_75t_SL g855 (.A(n_19188),
    .B(n_12813),
    .Y(n_12814));
 INVxp67_ASAP7_75t_SL g856 (.A(n_19188),
    .Y(n_12818));
 INVx1_ASAP7_75t_SL g86 (.A(n_22001),
    .Y(n_5639));
 OAI22xp5_ASAP7_75t_SL g860 (.A1(n_12813),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_n_757),
    .B2(n_12819),
    .Y(n_12820));
 INVxp67_ASAP7_75t_SL g865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .Y(n_12819));
 INVx1_ASAP7_75t_SL g866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_757),
    .Y(n_12813));
 MAJIxp5_ASAP7_75t_SL g87 (.A(n_12258),
    .B(n_3511),
    .C(n_3917),
    .Y(n_9614));
 XOR2xp5_ASAP7_75t_SL g88 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_74),
    .B(n_26099),
    .Y(n_19461));
 OAI21xp5_ASAP7_75t_SL g889 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_297),
    .A2(n_11481),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_295),
    .Y(n_11483));
 OAI21xp5_ASAP7_75t_SL g892 (.A1(n_10187),
    .A2(n_23433),
    .B(n_20500),
    .Y(n_11489));
 INVx1_ASAP7_75t_SL g893 (.A(n_11480),
    .Y(n_11481));
 OAI21x1_ASAP7_75t_SL g894 (.A1(n_11472),
    .A2(n_23433),
    .B(n_11479),
    .Y(n_11480));
 XNOR2xp5_ASAP7_75t_SL g898 (.A(n_11490),
    .B(n_11495),
    .Y(n_11496));
 NAND3xp33_ASAP7_75t_SL g899 (.A(n_11471),
    .B(n_19242),
    .C(n_9206),
    .Y(n_11487));
 INVx1_ASAP7_75t_SL g9 (.A(n_12643),
    .Y(n_12644));
 OAI21x1_ASAP7_75t_SL g90 (.A1(n_5376),
    .A2(n_15798),
    .B(n_5377),
    .Y(n_5378));
 AOI21xp5_ASAP7_75t_SL g900 (.A1(n_11473),
    .A2(n_11474),
    .B(n_22061),
    .Y(n_11475));
 AOI21xp33_ASAP7_75t_SRAM g901 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_32),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_262),
    .B(n_22061),
    .Y(n_11490));
 AOI22xp5_ASAP7_75t_SL g902 (.A1(n_11474),
    .A2(n_11493),
    .B1(n_17979),
    .B2(n_11492),
    .Y(n_11495));
 OA21x2_ASAP7_75t_SL g903 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_285),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_282),
    .Y(n_11479));
 NAND2xp5_ASAP7_75t_SL g904 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_262),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_32),
    .Y(n_11476));
 INVxp67_ASAP7_75t_SL g905 (.A(n_11471),
    .Y(n_11472));
 NOR2x1_ASAP7_75t_SL g906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283),
    .B(n_10187),
    .Y(n_11471));
 AND2x2_ASAP7_75t_SL g907 (.A(n_21503),
    .B(n_17979),
    .Y(n_11477));
 OR2x2_ASAP7_75t_SL g91 (.A(n_5375),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_93),
    .Y(n_5377));
 AND2x2_ASAP7_75t_SL g92 (.A(n_5375),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_93),
    .Y(n_5376));
 NAND2xp5_ASAP7_75t_SL g93 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .Y(n_5375));
 INVx1_ASAP7_75t_L g94 (.A(n_5422),
    .Y(n_5423));
 NAND2x1_ASAP7_75t_SL g95 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .Y(n_5422));
 AOI21xp5_ASAP7_75t_SL g951 (.A1(n_6219),
    .A2(n_6222),
    .B(n_6224),
    .Y(n_6230));
 XNOR2xp5_ASAP7_75t_SL g954 (.A(n_6219),
    .B(n_6232),
    .Y(n_6233));
 AOI22xp5_ASAP7_75t_SL g955 (.A1(n_6221),
    .A2(n_6224),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_240),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_255),
    .Y(n_6225));
 NAND2xp5_ASAP7_75t_SL g956 (.A(n_6221),
    .B(n_6222),
    .Y(n_6223));
 AOI21xp5_ASAP7_75t_SL g957 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_255),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_240),
    .B(n_6234),
    .Y(n_6235));
 AOI321xp33_ASAP7_75t_SL g9571__5477 (.A1(n_2100),
    .A2(n_333),
    .A3(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .B1(n_2115),
    .B2(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .C(n_2118),
    .Y(n_2121));
 AOI322xp5_ASAP7_75t_SL g9574__2398 (.A1(n_2102),
    .A2(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .A3(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .B1(u_NV_NVDLA_cmac_u_reg_n_1258),
    .B2(cmac_a2csb_resp_pd[12]),
    .C1(n_2115),
    .C2(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .Y(n_2120));
 AOI322xp5_ASAP7_75t_SL g9575__5107 (.A1(n_2102),
    .A2(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .A3(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .B1(u_NV_NVDLA_cmac_u_reg_n_1258),
    .B2(cmac_a2csb_resp_pd[13]),
    .C1(n_2115),
    .C2(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .Y(n_2119));
 NAND2xp5_ASAP7_75t_SL g958 (.A(n_6222),
    .B(n_6231),
    .Y(n_6232));
 INVx1_ASAP7_75t_SL g9582 (.A(n_2116),
    .Y(n_2118));
 AOI21xp5_ASAP7_75t_SL g9583__6260 (.A1(cmac_a2csb_resp_pd[16]),
    .A2(u_NV_NVDLA_cmac_u_reg_n_1258),
    .B(n_2110),
    .Y(n_2117));
 AOI322xp5_ASAP7_75t_SL g9584__4319 (.A1(n_2097),
    .A2(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .A3(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .B1(n_2098),
    .B2(n_2032),
    .C1(cmac_a2csb_resp_pd[0]),
    .C2(u_NV_NVDLA_cmac_u_reg_n_1258),
    .Y(n_2116));
 AOI22xp5_ASAP7_75t_SL g9589__8428 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[34]),
    .A2(n_2094),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .B2(n_2095),
    .Y(n_2114));
 INVx1_ASAP7_75t_SL g959 (.A(n_6219),
    .Y(n_6220));
 AOI22xp5_ASAP7_75t_SL g9590__5526 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .A2(n_2094),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .B2(n_2095),
    .Y(n_2113));
 AOI32xp33_ASAP7_75t_SL g9591__6783 (.A1(n_576),
    .A2(n_2098),
    .A3(n_333),
    .B1(cmac_a2csb_resp_pd[17]),
    .B2(u_NV_NVDLA_cmac_u_reg_n_1258),
    .Y(n_2112));
 AOI22xp5_ASAP7_75t_SL g9592__3680 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[35]),
    .A2(n_2094),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .B2(n_2095),
    .Y(n_2111));
 NOR2xp33_ASAP7_75t_SL g9593__1617 (.A(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .B(n_2101),
    .Y(n_2115));
 INVx1_ASAP7_75t_SL g9595 (.A(n_2106),
    .Y(n_2110));
 AOI32xp33_ASAP7_75t_SL g9596__2802 (.A1(n_2098),
    .A2(u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en),
    .A3(n_662),
    .B1(cmac_a2csb_resp_pd[1]),
    .B2(u_NV_NVDLA_cmac_u_reg_n_1258),
    .Y(n_2109));
 AOI22xp5_ASAP7_75t_SL g9597__1705 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[34]),
    .A2(n_2092),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .B2(n_2093),
    .Y(n_2108));
 AOI22xp5_ASAP7_75t_SL g9598__5122 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[35]),
    .A2(n_2092),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .B2(n_2093),
    .Y(n_2107));
 A2O1A1Ixp33_ASAP7_75t_SL g9599__8246 (.A1(n_2091),
    .A2(u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en),
    .B(n_2097),
    .C(n_662),
    .Y(n_2106));
 INVx1_ASAP7_75t_SL g96 (.A(n_13502),
    .Y(n_5570));
 AO21x2_ASAP7_75t_SL g960 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_248),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_251),
    .Y(n_6219));
 AOI22xp33_ASAP7_75t_SL g9600__7098 (.A1(n_2096),
    .A2(n_670),
    .B1(n_733),
    .B2(u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en),
    .Y(n_2105));
 AOI22xp33_ASAP7_75t_SL g9601__6131 (.A1(n_2096),
    .A2(n_669),
    .B1(n_19237),
    .B2(u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en),
    .Y(n_2104));
 AOI22xp5_ASAP7_75t_SL g9602__1881 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .A2(n_2092),
    .B1(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .B2(n_2093),
    .Y(n_2103));
 INVxp67_ASAP7_75t_SL g9603 (.A(n_2101),
    .Y(n_2102));
 NAND2xp5_ASAP7_75t_SL g9604__5115 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .B(n_2097),
    .Y(n_2101));
 AO21x1_ASAP7_75t_SL g9605__7482 (.A1(n_2091),
    .A2(n_573),
    .B(n_2097),
    .Y(n_2100));
 AOI22xp5_ASAP7_75t_SL g9606__4733 (.A1(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .A2(n_2089),
    .B1(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .B2(n_2088),
    .Y(n_2099));
 NOR2xp33_ASAP7_75t_SL g9607__6161 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .B(n_2090),
    .Y(n_2098));
 AND2x2_ASAP7_75t_SL g9608__9315 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .B(n_2091),
    .Y(n_2097));
 INVx1_ASAP7_75t_SL g9609 (.A(n_2095),
    .Y(n_2094));
 INVxp67_ASAP7_75t_SL g961 (.A(n_6221),
    .Y(n_6234));
 INVx1_ASAP7_75t_SL g9610 (.A(n_2093),
    .Y(n_2092));
 NOR3xp33_ASAP7_75t_SL g9611__9945 (.A(n_2086),
    .B(n_337),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .Y(n_2096));
 NAND3xp33_ASAP7_75t_SL g9612__2883 (.A(n_669),
    .B(n_2087),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .Y(n_2095));
 NAND3xp33_ASAP7_75t_SL g9613__2346 (.A(n_670),
    .B(n_2087),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .Y(n_2093));
 INVxp67_ASAP7_75t_SL g9614 (.A(n_2091),
    .Y(n_2090));
 NOR2xp33_ASAP7_75t_SL g9615__1666 (.A(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .B(n_2084),
    .Y(n_2091));
 INVx1_ASAP7_75t_SL g9616 (.A(n_2088),
    .Y(n_2089));
 INVxp67_ASAP7_75t_SL g9617 (.A(n_2086),
    .Y(n_2087));
 NAND4xp25_ASAP7_75t_SL g9618__7410 (.A(n_2085),
    .B(n_333),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .D(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .Y(n_2088));
 NAND3xp33_ASAP7_75t_SL g9619__6417 (.A(n_2085),
    .B(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .C(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .Y(n_2086));
 NAND2xp5_ASAP7_75t_SL g962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_241),
    .Y(n_6221));
 NAND2xp5_ASAP7_75t_SL g963 (.A(n_19141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_243),
    .Y(n_6222));
 INVx1_ASAP7_75t_SL g964 (.A(n_6224),
    .Y(n_6231));
 NOR2xp67_ASAP7_75t_SL g965 (.A(n_19141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_243),
    .Y(n_6224));
 INVx1_ASAP7_75t_SL g966 (.A(n_9392),
    .Y(n_6218));
 NAND2xp67_ASAP7_75t_SL g970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_17),
    .Y(n_12975));
 INVx1_ASAP7_75t_SL g972 (.A(n_24669),
    .Y(n_12978));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_904),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_903),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_892),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_889),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_902),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_897),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_888),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_891),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_890),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1391),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1388),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1385),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1376),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1372),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1365),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1364),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1451),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_in_dat_pd_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1363),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pd_d2[8]));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1_reg (.CLK(nvdla_core_clk),
    .D(n_3),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d1));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2_reg (.CLK(nvdla_core_clk),
    .D(n_27),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pvld_d2));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_391),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .SE(n_661),
    .SI(n_4462));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_443),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .SE(n_833),
    .SI(n_2718));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_432),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .SE(n_833),
    .SI(n_22836));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_382),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[12]),
    .SE(n_833),
    .SI(n_4268));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_411),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .SE(n_833),
    .SI(n_3873));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_374),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .SE(n_833),
    .SI(n_3113));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_433),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .SE(n_833),
    .SI(n_15046));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_418),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .SE(n_621),
    .SI(n_2524));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_55),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .SE(n_621),
    .SI(n_4315));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_360),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .SE(n_621),
    .SI(n_2465));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_48),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[19]),
    .SE(n_621),
    .SI(n_4385));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_50),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .SE(n_661),
    .SI(n_3759));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_368),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[20]),
    .SE(n_621),
    .SI(n_16751));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_49),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .SE(n_621),
    .SI(n_2841));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_446),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .SE(n_621),
    .SI(n_15013));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_402),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .SE(n_621),
    .SI(n_2552));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_429),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .SE(n_626),
    .SI(n_2943));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_414),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .SE(n_626),
    .SI(n_3332));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_370),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .SE(n_626),
    .SI(n_14181));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_381),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[27]),
    .SE(n_626),
    .SI(n_3433));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_400),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[28]),
    .SE(n_626),
    .SI(n_14977));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_444),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .SE(n_626),
    .SI(n_3493));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_460),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[2]),
    .SE(n_661),
    .SI(n_2865));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_406),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .SE(n_626),
    .SI(n_2384));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_405),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .SE(n_626),
    .SI(n_2298));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_372),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .SE(n_838),
    .SI(n_3170));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_54),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .SE(n_838),
    .SI(n_3398));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_422),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[34]),
    .SE(n_838),
    .SI(n_3224));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_395),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[35]),
    .SE(n_838),
    .SI(n_18034));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_346),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[36]),
    .SE(n_838),
    .SI(n_22742));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_348),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .SE(n_838),
    .SI(n_15200));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_353),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .SE(n_838),
    .SI(n_4124));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_373),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[39]),
    .SE(n_838),
    .SI(n_428));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_47),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[3]),
    .SE(n_661),
    .SI(n_2766));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_359),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .SE(n_849),
    .SI(n_18050));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_431),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .SE(n_849),
    .SI(n_23277));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_453),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[42]),
    .SE(n_849),
    .SI(n_3314));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_385),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[43]),
    .SE(n_849),
    .SI(n_22638));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_366),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[44]),
    .SE(n_849),
    .SI(n_16764));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_425),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .SE(n_849),
    .SI(n_3714));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_354),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[46]),
    .SE(n_849),
    .SI(n_407));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_423),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[47]),
    .SE(n_849),
    .SI(n_434));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_341),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .SE(n_22863),
    .SI(n_20463));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_344),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .SE(n_22863),
    .SI(n_3409));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_416),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[4]),
    .SE(n_661),
    .SI(n_2331));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_22864),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .SE(n_22863),
    .SI(n_22866));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_457),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[51]),
    .SE(n_22863),
    .SI(n_3469));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_343),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[52]),
    .SE(n_22863),
    .SI(n_2934));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_347),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .SE(n_22863),
    .SI(n_3593));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_413),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .SE(n_22863),
    .SI(n_2700));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_449),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .SE(n_22863),
    .SI(n_2366));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_355),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .SE(n_828),
    .SI(n_2747));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_376),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[57]),
    .SE(n_828),
    .SI(n_13230));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_388),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .SE(n_828),
    .SI(n_12134));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_398),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .SE(n_828),
    .SI(n_3527));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_452),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .SE(n_661),
    .SI(n_2673));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_351),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[60]),
    .SE(n_828),
    .SI(n_2821));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_365),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .SE(n_828),
    .SI(n_3376));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_403),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .SE(n_828),
    .SI(n_4555));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_417),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[63]),
    .SE(n_828),
    .SI(n_3633));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_364),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .SE(n_661),
    .SI(n_3265));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_339),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .SE(n_661),
    .SI(n_3149));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_358),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .SE(n_833),
    .SI(n_4528));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_data_reg0_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_397),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .SE(n_833),
    .SI(n_2507));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1314),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1313),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1312),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1311),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1310),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1309),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1308),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_nz_reg0_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1307),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_actv_pvld_reg0_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_26),
    .QN(u_NV_NVDLA_cmac_u_core_dat0_actv_pvld[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_dat_actv_stripe_end_reg (.CLK(nvdla_core_clk),
    .D(n_2144),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_actv_stripe_end),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1681),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1669),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1663),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1668),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1667),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1666),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1665),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1664),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1660),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1662),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1661),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1678),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1659),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1658),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1657),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1656),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1655),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1654),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1653),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1652),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1651),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1650),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1677),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1649),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1648),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1647),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1646),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1645),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1644),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1643),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1642),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1641),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1640),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1676),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1639),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1638),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1637),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1635),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1636),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1634),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1633),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1632),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1631),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1629),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1675),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1630),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1628),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1627),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1626),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1625),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1624),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1623),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1622),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1621),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1620),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1672),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1619),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1618),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1617),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1616),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1674),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1673),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1671),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1670),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_901),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_900),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_899),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_898),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_896),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_895),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_894),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_893),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_3),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_pvld_3521),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_end_reg (.CLK(nvdla_core_clk),
    .D(n_2137),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_end_3520),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_st_reg (.CLK(nvdla_core_clk),
    .D(n_2139),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_dat_pre_stripe_st_3519),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_677),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .SE(n_820),
    .SI(n_261));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_574),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_796),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_765),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .SE(n_820),
    .SI(n_306));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_771),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .SE(n_820),
    .SI(n_196));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_785),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_510),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .SE(n_820),
    .SI(n_4048));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_531),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .SE(n_820),
    .SI(n_68));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_810),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .SE(n_820),
    .SI(n_103));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_511),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .SE(n_820),
    .SI(n_220));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_528),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .SE(n_820),
    .SI(n_57));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_549),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .SE(n_820),
    .SI(n_56));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_564),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .SE(n_820),
    .SI(n_229));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_466),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .SE(n_820),
    .SI(n_67));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_472),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .SE(n_820),
    .SI(n_266));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_520),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .SE(n_820),
    .SI(n_288));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_483),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .SE(n_820),
    .SI(n_157));
 SDFHx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[25]  (.CLK(nvdla_core_clk),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[25]),
    .D(n_519),
    .SE(n_820),
    .SI(n_214));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_516),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .SE(n_820),
    .SI(n_209));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_504),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .SE(n_820),
    .SI(n_153));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_508),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .SE(n_820),
    .SI(n_245));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_538),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .SE(n_820),
    .SI(n_267));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_721),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .SE(n_820),
    .SI(n_94));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_569),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .SE(n_820),
    .SI(n_218));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_774),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .SE(n_820),
    .SI(n_309));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_577),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .SE(n_820),
    .SI(n_251));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_794),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .SE(n_820),
    .SI(n_126));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_719),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .SE(n_820),
    .SI(n_98));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_499),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .SE(n_820),
    .SI(n_142));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_561),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .SE(n_820),
    .SI(n_254));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_521),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .SE(n_820),
    .SI(n_292));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_801),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .SE(n_820),
    .SI(n_88));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_769),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .SE(n_820),
    .SI(n_311));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_548),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .SE(n_820),
    .SI(n_257));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_575),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .SE(n_820),
    .SI(n_58));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_775),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .SE(n_820),
    .SI(n_207));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_735),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .SE(n_820),
    .SI(n_289));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_673),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .SE(n_820),
    .SI(n_262));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_578),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .SE(n_820),
    .SI(n_4354));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_702),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .SE(n_820),
    .SI(n_236));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_704),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .SE(n_820),
    .SI(n_95));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_490),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .SE(n_820),
    .SI(n_166));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_766),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .SE(n_820),
    .SI(n_71));
 SDFHx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[49]  (.CLK(nvdla_core_clk),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[49]),
    .D(n_802),
    .SE(n_820),
    .SI(n_59));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_547),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .SE(n_820),
    .SI(n_187));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_486),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .SE(n_820),
    .SI(n_158));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_684),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .SE(n_820),
    .SI(n_256));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_479),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .SE(n_820),
    .SI(n_221));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_463),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .SE(n_820),
    .SI(n_250));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_485),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .SE(n_820),
    .SI(n_78));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_725),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .SE(n_820),
    .SI(n_198));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_565),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_517),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .SE(n_820),
    .SI(n_92));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_470),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_570),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_763),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .SE(n_820),
    .SI(n_84));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_777),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .SE(n_820),
    .SI(n_170));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_568),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .SE(n_820),
    .SI(n_143));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_473),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_779),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .SE(n_820),
    .SI(n_4140));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_542),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .SE(n_820),
    .SI(n_301));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_493),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .SE(n_820),
    .SI(n_199));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_502),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .SE(n_820),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_539),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .SE(n_820),
    .SI(n_217));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2007),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2006),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2005),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2004),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2003),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2002),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2001),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2000),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_actv_pvld_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2080),
    .QN(u_NV_NVDLA_cmac_u_core_wt0_actv_pvld[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1749),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1995),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1994),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1993),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1991),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1992),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1990),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1989),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1988),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1987),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1985),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1748),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1986),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1984),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1983),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1982),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1979),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1972),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1971),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1968),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1964),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1960),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1747),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1956),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1953),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1952),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1945),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1943),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1939),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1936),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1932),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1930),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1923),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1746),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1922),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1917),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1913),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1910),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1909),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1902),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1901),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1898),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1894),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1892),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1745),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1891),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1889),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1890),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1888),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1887),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1885),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1886),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1884),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1883),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1882),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1744),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1881),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1880),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1879),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1878),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1999),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1998),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1997),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1996),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_879),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_878),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_877),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_876),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_875),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_874),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_873),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_872),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_4413),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt0_sd_pvld_3195),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_740),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .SE(n_17240),
    .SI(n_294));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_718),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_716),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_713),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .SE(n_17240),
    .SI(n_191));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_710),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .SE(n_17240),
    .SI(n_279));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_709),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_708),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .SE(n_17240),
    .SI(n_3957));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_784),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .SE(n_17240),
    .SI(n_194));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_706),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .SE(n_17240),
    .SI(n_295));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_787),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .SE(n_17240),
    .SI(n_300));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_791),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .SE(n_17240),
    .SI(n_297));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_739),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .SE(n_17240),
    .SI(n_179));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_813),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .SE(n_17240),
    .SI(n_308));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_729),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .SE(n_17240),
    .SI(n_172));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_497),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .SE(n_17240),
    .SI(n_228));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_701),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .SE(n_17240),
    .SI(n_296));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_700),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .SE(n_17240),
    .SI(n_73));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_699),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .SE(n_17240),
    .SI(n_145));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_698),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .SE(n_17240),
    .SI(n_223));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_465),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .SE(n_17240),
    .SI(n_125));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_694),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .SE(n_17240),
    .SI(n_150));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_692),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .SE(n_17240),
    .SI(n_211));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_738),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .SE(n_17240),
    .SI(n_131));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_691),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .SE(n_17240),
    .SI(n_152));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_481),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .SE(n_17240),
    .SI(n_146));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_690),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .SE(n_17240),
    .SI(n_238));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_689),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .SE(n_17240),
    .SI(n_240));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_696),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .SE(n_17240),
    .SI(n_242));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_688),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .SE(n_17240),
    .SI(n_210));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_494),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .SE(n_17240),
    .SI(n_246));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_686),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .SE(n_17240),
    .SI(n_138));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_685),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .SE(n_17240),
    .SI(n_181));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_683),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .SE(n_17240),
    .SI(n_230));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_816),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .SE(n_17240),
    .SI(n_164));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_682),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .SE(n_17240),
    .SI(n_83));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_506),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .SE(n_17240),
    .SI(n_93));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_679),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .SE(n_17240),
    .SI(n_161));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_678),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .SE(n_17240),
    .SI(n_124));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_676),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .SE(n_17240),
    .SI(n_185));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_675),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .SE(n_17240),
    .SI(n_183));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_715),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .SE(n_17240),
    .SI(n_105));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_529),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .SE(n_17240),
    .SI(n_237));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_680),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .SE(n_17240),
    .SI(n_286));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_17241),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .SE(n_17240),
    .SI(n_17242));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_507),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .SE(n_17240),
    .SI(n_277));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_703),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .SE(n_17240),
    .SI(n_252));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_711),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .SE(n_17240),
    .SI(n_189));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_724),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .SE(n_17240),
    .SI(n_117));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_551),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .SE(n_17240),
    .SI(n_307));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_728),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .SE(n_17240),
    .SI(n_62));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_742),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .SE(n_17240),
    .SI(n_107));
 SDFHx4_ASAP7_75t_L \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_730),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_741),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .SE(n_17240),
    .SI(n_177));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_749),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_754),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_46));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_732),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .SE(n_17240),
    .SI(n_184));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_755),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .SE(n_17240),
    .SI(n_291));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_752),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .SE(n_17240),
    .SI(n_182));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_759),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_761),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .SE(n_17240),
    .SI(n_4239));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_731),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .SE(n_17240),
    .SI(n_91));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_727),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .SE(n_17240),
    .SI(n_129));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_726),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .SE(n_17240),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_720),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .SE(n_17240),
    .SI(n_160));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2023),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2022),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2021),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2020),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2019),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2018),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2017),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2016),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_actv_pvld_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2082),
    .QN(u_NV_NVDLA_cmac_u_core_wt1_actv_pvld[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1877),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1867),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1866),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1865),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1864),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1863),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1862),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1861),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1860),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1859),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1858),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1876),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1857),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1856),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1855),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1854),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1853),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1852),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1851),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1850),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1849),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1848),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1875),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1847),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1846),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1845),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1844),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1843),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1842),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1841),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1840),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1839),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1838),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1874),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1837),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1836),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1835),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1834),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1833),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1832),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1831),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1830),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1829),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1828),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1873),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1827),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1826),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1825),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1824),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1823),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1822),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1821),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1820),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1819),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1818),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1872),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1817),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1816),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1815),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1814),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1871),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1870),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1869),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1868),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_871),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_870),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_869),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_868),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_867),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_866),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_865),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_864),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_4414),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt1_sd_pvld_3196),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_558),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .SE(n_580),
    .SI(n_120));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_553),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_758),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_550),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .SE(n_580),
    .SI(n_168));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_717),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .SE(n_580),
    .SI(n_260));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_722),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_734),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .SE(n_580),
    .SI(n_3965));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_744),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .SE(n_580),
    .SI(n_77));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_747),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .SE(n_580),
    .SI(n_114));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_753),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .SE(n_580),
    .SI(n_280));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_545),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .SE(n_580),
    .SI(n_72));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_707),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .SE(n_580),
    .SI(n_154));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_544),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .SE(n_580),
    .SI(n_64));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_543),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .SE(n_580),
    .SI(n_102));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_556),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .SE(n_580),
    .SI(n_162));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_541),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .SE(n_580),
    .SI(n_132));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_540),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .SE(n_580),
    .SI(n_155));
 SDFHx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[25]  (.CLK(nvdla_core_clk),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[25]),
    .D(n_500),
    .SE(n_580),
    .SI(n_253));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_503),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .SE(n_580),
    .SI(n_275));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_505),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .SE(n_580),
    .SI(n_80));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_562),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .SE(n_580),
    .SI(n_134));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_571),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .SE(n_580),
    .SI(n_305));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_557),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .SE(n_580),
    .SI(n_173));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_572),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .SE(n_580),
    .SI(n_116));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_757),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .SE(n_580),
    .SI(n_174));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_712),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .SE(n_580),
    .SI(n_259));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_756),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .SE(n_580),
    .SI(n_82));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_764),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .SE(n_580),
    .SI(n_192));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_767),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .SE(n_580),
    .SI(n_135));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_768),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[36]),
    .SE(n_580),
    .SI(n_165));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_772),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .SE(n_580),
    .SI(n_293));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_778),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .SE(n_580),
    .SI(n_208));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_781),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .SE(n_580),
    .SI(n_287));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_809),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .SE(n_580),
    .SI(n_215));
 SDFHx4_ASAP7_75t_L \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_789),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .SE(n_580),
    .SI(n_188));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_533),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .SE(n_580),
    .SI(n_203));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_530),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .SE(n_580),
    .SI(n_193));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_527),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .SE(n_580),
    .SI(n_255));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_773),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .SE(n_580),
    .SI(n_70));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_513),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .SE(n_580),
    .SI(n_272));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_811),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .SE(n_580),
    .SI(n_232));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_792),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .SE(n_580),
    .SI(n_76));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_492),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .SE(n_580),
    .SI(n_87));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_526),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .SE(n_580),
    .SI(n_20503));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_555),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .SE(n_580),
    .SI(n_176));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_705),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .SE(n_580),
    .SI(n_159));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_477),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .SE(n_580),
    .SI(n_263));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_467),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .SE(n_580),
    .SI(n_139));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_524),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .SE(n_580),
    .SI(n_285));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_522),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .SE(n_580),
    .SI(n_213));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_474),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .SE(n_580),
    .SI(n_106));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_478),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_480),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .SE(n_580),
    .SI(n_104));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_482),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_523),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_537),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .SE(n_580),
    .SI(n_265));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_487),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .SE(n_580),
    .SI(n_243));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_489),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .SE(n_580),
    .SI(n_283));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_498),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_560),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .SE(n_580),
    .SI(n_4253));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_697),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .SE(n_580),
    .SI(n_205));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_554),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .SE(n_580),
    .SI(n_156));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_512),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .SE(n_580),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_814),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .SE(n_580),
    .SI(n_231));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2015),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2014),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2013),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2012),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2011),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2010),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2009),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2008),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_actv_pvld_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2081),
    .QN(u_NV_NVDLA_cmac_u_core_wt2_actv_pvld[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1813),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1803),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1802),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1801),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1800),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1799),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1798),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1797),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1796),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1795),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1794),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1812),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1793),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1792),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1791),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1790),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1789),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1788),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1787),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1786),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1785),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1784),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1811),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1783),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1782),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1781),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1780),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1779),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1778),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1777),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1776),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1775),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1774),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1810),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1773),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1772),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1771),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1770),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1769),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1768),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1767),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1766),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1765),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1764),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1809),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1763),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1762),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1761),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1760),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1759),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1758),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1757),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1756),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1755),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1754),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1808),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1753),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1752),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1751),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1750),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1807),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1806),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1805),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1804),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_856),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_857),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_858),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_863),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_859),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_861),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_862),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_860),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_4415),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt2_sd_pvld_3197),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_681),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .SE(n_582),
    .SI(n_90));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_736),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_546),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_46));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_552),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .SE(n_582),
    .SI(n_310));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_476),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .SE(n_582),
    .SI(n_299));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_518),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .SE(n_582),
    .SI(n_202));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_566),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .SE(n_582),
    .SI(n_3975));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_790),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .SE(n_582),
    .SI(n_269));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_762),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .SE(n_582),
    .SI(n_281));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_745),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .SE(n_582),
    .SI(n_118));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_495),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .SE(n_582),
    .SI(n_200));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_484),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .SE(n_582),
    .SI(n_186));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_746),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .SE(n_582),
    .SI(n_130));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_782),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .SE(n_582),
    .SI(n_144));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_471),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .SE(n_582),
    .SI(n_99));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_693),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .SE(n_582),
    .SI(n_112));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_468),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .SE(n_582),
    .SI(n_226));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_695),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .SE(n_582),
    .SI(n_101));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_751),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .SE(n_582),
    .SI(n_273));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_770),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .SE(n_582),
    .SI(n_140));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_723),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .SE(n_582),
    .SI(n_111));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_750),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .SE(n_582),
    .SI(n_244));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_567),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .SE(n_582),
    .SI(n_61));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_464),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .SE(n_582),
    .SI(n_79));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_743),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .SE(n_582),
    .SI(n_222));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_748),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .SE(n_582),
    .SI(n_284));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_475),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .SE(n_582),
    .SI(n_147));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_496),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .SE(n_582),
    .SI(n_190));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_532),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .SE(n_582),
    .SI(n_298));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_534),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .SE(n_582),
    .SI(n_268));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_535),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .SE(n_582),
    .SI(n_151));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_559),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .SE(n_582),
    .SI(n_206));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_776),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .SE(n_582),
    .SI(n_74));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_525),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .SE(n_582),
    .SI(n_195));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_815),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .SE(n_582),
    .SI(n_63));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_780),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .SE(n_582),
    .SI(n_225));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_783),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .SE(n_582),
    .SI(n_85));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_788),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .SE(n_582),
    .SI(n_123));
 SDFHx4_ASAP7_75t_L \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_793),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .SE(n_582),
    .SI(n_276));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_795),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .SE(n_582),
    .SI(n_122));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_812),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .SE(n_582),
    .SI(n_119));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_501),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .SE(n_582),
    .SI(n_60));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_714),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .SE(n_582),
    .SI(n_163));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_674),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .SE(n_582),
    .SI(n_304));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_509),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .SE(n_582),
    .SI(n_219));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_808),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .SE(n_582),
    .SI(n_96));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_806),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .SE(n_582),
    .SI(n_258));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_805),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .SE(n_582),
    .SI(n_216));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_804),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .SE(n_582),
    .SI(n_178));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_563),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .SE(n_582),
    .SI(n_113));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_515),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .SE(n_582),
    .SI(n_169));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_803),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_799),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .SE(n_582),
    .SI(n_175));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_786),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_43));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_800),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_46));
 SDFHx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_491),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .SE(n_582),
    .SI(n_148));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_798),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .SE(n_582),
    .SI(n_290));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_807),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .SE(n_582),
    .SI(n_201));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_737),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_47));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_797),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .SE(n_582),
    .SI(n_4262));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_488),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .SE(n_582),
    .SI(n_224));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_469),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .SE(n_582),
    .SI(n_89));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_760),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .SE(n_582),
    .SI(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_40));
 SDFHx4_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_536),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .SE(n_582),
    .SI(n_149));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2031),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2030),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2029),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2028),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2027),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2026),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2025),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2024),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_actv_pvld_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1599),
    .QN(u_NV_NVDLA_cmac_u_core_wt3_actv_pvld[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1981),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1967),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1966),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1965),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1963),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1962),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1961),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1959),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1958),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1957),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1955),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1980),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1954),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1951),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1950),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1949),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1948),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1947),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1946),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1944),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1942),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1941),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1978),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1940),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1938),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1937),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1935),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1934),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1933),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1931),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1929),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1928),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1927),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1977),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1926),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1925),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1924),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1921),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1920),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1919),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1918),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1916),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1915),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1914),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1976),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1912),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1911),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1908),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1907),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1906),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1905),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1904),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1903),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1900),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1899),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1975),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1897),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1896),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1895),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1893),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1974),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1973),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1970),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1969),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_887),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_886),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_885),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_884),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_883),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_882),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_881),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_880),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_4412),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt3_sd_pvld_3198),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1743),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1733),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1732),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1731),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1730),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1729),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1728),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1727),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1726),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1725),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[19]  (.CLK(nvdla_core_clk),
    .D(n_1724),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[19]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1742),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[20]  (.CLK(nvdla_core_clk),
    .D(n_1723),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[20]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[21]  (.CLK(nvdla_core_clk),
    .D(n_1722),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[21]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1721),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[22]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[23]  (.CLK(nvdla_core_clk),
    .D(n_1720),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[23]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[24]  (.CLK(nvdla_core_clk),
    .D(n_1719),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[24]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[25]  (.CLK(nvdla_core_clk),
    .D(n_1718),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[25]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[26]  (.CLK(nvdla_core_clk),
    .D(n_1717),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[26]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[27]  (.CLK(nvdla_core_clk),
    .D(n_1716),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[27]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[28]  (.CLK(nvdla_core_clk),
    .D(n_1715),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[28]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[29]  (.CLK(nvdla_core_clk),
    .D(n_1714),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[29]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1741),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[30]  (.CLK(nvdla_core_clk),
    .D(n_1713),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[30]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[31]  (.CLK(nvdla_core_clk),
    .D(n_1712),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[31]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[32]  (.CLK(nvdla_core_clk),
    .D(n_1711),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[32]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_1710),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[33]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1709),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[34]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1708),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[35]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[36]  (.CLK(nvdla_core_clk),
    .D(n_1707),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[36]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[37]  (.CLK(nvdla_core_clk),
    .D(n_1706),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[37]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[38]  (.CLK(nvdla_core_clk),
    .D(n_1705),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[38]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[39]  (.CLK(nvdla_core_clk),
    .D(n_1704),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[39]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1740),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[40]  (.CLK(nvdla_core_clk),
    .D(n_1703),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[40]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[41]  (.CLK(nvdla_core_clk),
    .D(n_1702),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[41]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[42]  (.CLK(nvdla_core_clk),
    .D(n_1701),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[42]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[43]  (.CLK(nvdla_core_clk),
    .D(n_1700),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[43]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[44]  (.CLK(nvdla_core_clk),
    .D(n_1699),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[44]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[45]  (.CLK(nvdla_core_clk),
    .D(n_1698),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[45]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[46]  (.CLK(nvdla_core_clk),
    .D(n_1697),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[46]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[47]  (.CLK(nvdla_core_clk),
    .D(n_1696),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[47]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[48]  (.CLK(nvdla_core_clk),
    .D(n_1695),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[48]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[49]  (.CLK(nvdla_core_clk),
    .D(n_1694),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[49]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1739),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[50]  (.CLK(nvdla_core_clk),
    .D(n_1693),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[50]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[51]  (.CLK(nvdla_core_clk),
    .D(n_1692),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[51]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[52]  (.CLK(nvdla_core_clk),
    .D(n_1691),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[52]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[53]  (.CLK(nvdla_core_clk),
    .D(n_1690),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[53]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1689),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[54]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1688),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[55]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[56]  (.CLK(nvdla_core_clk),
    .D(n_1687),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[56]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[57]  (.CLK(nvdla_core_clk),
    .D(n_1686),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[57]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[58]  (.CLK(nvdla_core_clk),
    .D(n_1685),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[58]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[59]  (.CLK(nvdla_core_clk),
    .D(n_1684),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[59]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1738),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[60]  (.CLK(nvdla_core_clk),
    .D(n_1683),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[60]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[61]  (.CLK(nvdla_core_clk),
    .D(n_1682),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[61]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[62]  (.CLK(nvdla_core_clk),
    .D(n_1680),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[62]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[63]  (.CLK(nvdla_core_clk),
    .D(n_1679),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[63]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1737),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1736),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1735),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1734),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_data[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1306),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1305),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1304),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1303),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1302),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1301),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1300),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1299),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_nz[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2140),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2136),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2135),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2138),
    .QN(u_NV_NVDLA_cmac_u_core_u_active_wt_pre_sel[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_448),
    .B(n_3938),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_180));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g20733 (.A(n_23976),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_366),
    .Y(n_12190));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g20737 (.A(n_23976),
    .Y(n_12191));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g24095 (.A1(n_10205),
    .A2(n_3560),
    .B(n_18084),
    .Y(n_16160));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g24249 (.A(n_19445),
    .B(n_10841),
    .Y(n_16316));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g26367 (.A1(n_5683),
    .A2(n_18579),
    .B1(n_5681),
    .B2(n_18580),
    .Y(n_18581));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g26370 (.A(n_18579),
    .Y(n_18580));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g29958 (.A(n_22608),
    .B(n_22609),
    .Y(n_22610));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g29959 (.A1(n_9513),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .B(n_22610),
    .Y(n_22612));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g29960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_430),
    .B(n_23495),
    .Y(n_22614));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g30160 (.A1(n_10290),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_421),
    .B(n_22850),
    .Y(n_22851));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g31200 (.A(n_23974),
    .B(n_12188),
    .Y(n_23976));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6011 (.A1(n_3668),
    .A2(n_10455),
    .B(n_3736),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_500));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6024 (.A1(n_12780),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_440),
    .B(n_22851),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_489));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6029 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_439),
    .B(n_3560),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_178));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6033 (.A(n_11385),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_481),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_177));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_481));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6035 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_480));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6036 (.A(n_3208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_450),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_176));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_472),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_64));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6039 (.A1(n_22611),
    .A2(n_9367),
    .B(n_22612),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_478));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_472),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_175));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6042 (.A(n_9367),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_475));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6045 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_386),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_383),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_472));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6051 (.A(n_12190),
    .B(n_21266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_466));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6052 (.A(n_12190),
    .B(n_4087),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_465));
 INVxp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6055 (.A(n_21480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_462));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6057 (.A(n_21266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_455));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_453));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6062 (.A(n_3737),
    .B(n_3669),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_451));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6063 (.A(n_2850),
    .B(n_16316),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_458));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_432),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_450));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6071 (.A(n_12190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_445));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_173));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6074 (.A(n_3988),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_421),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_440));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6075 (.A(n_10205),
    .B(n_18085),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_439));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6077 (.A(n_10290),
    .B(n_3987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_448));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_379),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_387),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_437));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_408),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_404),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_436));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6080 (.A(n_12191),
    .B(n_6601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_446));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6082 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_443));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_432));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_430));
 INVxp33_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6087 (.A(n_16316),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_425));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6089 (.A(n_10290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_424));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_433));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6095 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_431));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6096 (.A(n_22608),
    .B(n_22609),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_429));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6101 (.A(n_10419),
    .B(n_22037),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_62));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6102 (.A(n_22848),
    .B(n_22849),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_421));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6109 (.A(n_12779),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_408));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_380),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_172));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6113 (.A(n_12774),
    .B(n_12775),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_404));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6125 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_397));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_386),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_384),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_396));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_401));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6130 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_356),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_398));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_347),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_395));
 MAJIxp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6139 (.A(n_24681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .C(n_6078),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_387));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_383),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_384));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_345),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_171));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_353),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_360),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_386));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_385));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_381));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6145 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_380));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_353),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_360),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_383));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_308),
    .B(n_10512),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_379));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6149 (.A(n_22035),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_303),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_377));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6154 (.A(n_6601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_366));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6157 (.A(n_12817),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_372));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .C(n_13175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_363));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_356));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6169 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .A2(n_12817),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_354));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_361));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_360));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_359));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_358));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_325),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_353));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6177 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_304),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_305),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_349));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6180 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .A2(n_13176),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_347));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_352));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6183 (.A1(n_19068),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_345));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_344));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6196 (.A(n_12817),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_330));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_337));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_328));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6201 (.A(n_19068),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_327));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_326));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6203 (.A(n_19068),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_336));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6208 (.A(n_22320),
    .B(n_26052),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_58));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6210 (.A(n_22972),
    .B(n_17401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_332));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6213 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_325));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_322));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6219 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_314));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_308));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_324));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_321));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_318));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6233 (.A(n_10505),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_315));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6234 (.A(n_19186),
    .B(n_12818),
    .C(n_12820),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_312));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6239 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_305));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6242 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_300));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6243 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_307));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6246 (.A(n_11295),
    .B(n_10143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_304));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6248 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_24),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_303));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6257 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_52));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_290));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6266 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_289));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6267 (.A(n_6045),
    .B(n_8053),
    .C(n_18154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_288));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6272 (.A1(n_19865),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_281));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6274 (.A(n_8476),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_279));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6279 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .B2(n_2741),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_277));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6282 (.A(n_18064),
    .B(n_18067),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_275));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_283));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6286 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_51));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6289 (.A(n_22320),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_267));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6290 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_265));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6293 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_254));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6301 (.A(n_11433),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_264));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_263));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6304 (.A(n_19069),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .C(n_19071),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_261));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6305 (.A(n_19070),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_260));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6306 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_259));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6307 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_216),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_258));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6309 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_250));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_251));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6324 (.A(n_23551),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_243));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_240));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6328 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_137),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_164),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_138),
    .B2(n_11377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_239));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_237));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6337 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_233));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_231));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_229));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6351 (.A(n_18155),
    .B(n_19867),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_232));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6352 (.A(n_19867),
    .B(n_9246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_230));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6353 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_697),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_228));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6354 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_227));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6356 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6362 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_221));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6363 (.A(n_18582),
    .B(n_9234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_220));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6365 (.A(n_21998),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_218));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_216));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6374 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6376 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_204));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6377 (.A1(n_19866),
    .A2(n_8053),
    .B1(n_19865),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_203));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6379 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6380 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_215));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_75),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_212));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6389 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_209));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6390 (.A(n_18803),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_657),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_207));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_152),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_655),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_623),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_206));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6394 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_195));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6405 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_200));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6409 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_721),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6412 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_663),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_699),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_190));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_633),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_185));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6423 (.A(n_11433),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_170));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6424 (.A(n_11377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6430 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_797),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_181));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6434 (.B(n_19556),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_176),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_709));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6436 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_174));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6439 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_745),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6441 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_168));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6442 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_167));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6444 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_729),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6448 (.A(n_19428),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_156));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6450 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_152));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6451 (.A(n_22002),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_601),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_88),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_161));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6459 (.A(n_19065),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_767),
    .C(n_19064),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6463 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_785),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_721),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6466 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_733),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_637),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_797),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6467 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_691),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_145));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_553),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_713),
    .C(n_22441),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_639),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_671),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_143));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_745),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_585),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_681),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_141));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6472 (.A(n_13474),
    .B(n_5929),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_583),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6473 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6474 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_135));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_131));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6477 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_129));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6492 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_757),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_693),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_597),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_137));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6493 (.A(n_12785),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_611),
    .C(n_9874),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6494 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_701),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_793),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_729),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_130));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6497 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_599),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_727),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_567),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_128));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6499 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_591),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_751),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_126));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6500 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_695),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_663),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_125));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_761),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_665),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_633),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_123));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_763),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_635),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_667),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_122));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_603),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_731),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_n_699),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_121));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6505 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_747),
    .B(n_21638),
    .C(n_21639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_120));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_597),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_693),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_111));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6514 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_761),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_109));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_791),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_695),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_108));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_667),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_763),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_107));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_106));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6524 (.A(n_13544),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_547),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_104));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6525 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_623),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_655),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_103));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6530 (.A(n_19054),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_575),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_115));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_625),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_100));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_565),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_98));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6544 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_629),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_661),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_97));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6545 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_731),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_96));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6548 (.A(n_8482),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_615),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_94));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6551 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_567),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_599),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_92));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_637),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_733),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_91));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6553 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_90));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_691),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_89));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6556 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_571),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_102));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_795),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6559 (.A(n_9235),
    .B(n_5733),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_575),
    .B(n_19054),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_85));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6562 (.A(n_5733),
    .B(n_9235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_82));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6564 (.A(n_8482),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_615),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6565 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_615),
    .B(n_8482),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_80));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6581 (.A(n_9795),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_74));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6586 (.A(n_9793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_72));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6621 (.A(n_22973),
    .B(n_10501),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_34));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6622 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .A(n_6119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6629 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_26));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6630 (.A(n_19070),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_25));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6631 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_24));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6633 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(n_22076),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_22));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6637 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_621),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_653),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_18));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6641 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_581),
    .B(n_22312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_14));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6643 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_591),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_12));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6645 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_769),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_10),
    .A(n_21519));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6647 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_785),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_561),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6650 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_585),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_5));
 XNOR2x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_g6652 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_n_689),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_csa_tree_ADD_TC_OP_6_groupi_n_3),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_n_593));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g20834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_36),
    .Y(n_12290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g29208 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_6965),
    .Y(n_21798));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2959 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_268),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_270),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_197),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_736));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_271),
    .B(n_10056),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_744));
 OAI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2966 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_264),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_265),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_742));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_748));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2969 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_263),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_287),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_294));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_293));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2972 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_287),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_24));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2975 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_274),
    .A2(n_21401),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_273),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_287),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_750));
 OA211x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_283),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_280),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_282),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_289));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2978 (.A(n_21401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_287));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2980 (.A(n_21400),
    .B(n_21397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_752));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_277),
    .B(n_4085),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_285));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_284));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_283));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_282));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2985 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_281));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2986 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_258),
    .A2(n_21654),
    .B(n_26038),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2989 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_23));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_278));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_277));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2992 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_245),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_276));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2993 (.A(n_21654),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_275));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2994 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_274));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_273));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_271));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g2998 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_239),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_270));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3000 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_241),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_22));
 XNOR2x2_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_754));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_265));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3003 (.A(n_26038),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_262));
 NOR2xp33_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_268));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_264));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_248),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_263));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_260));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_256));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_259));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_258));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3018 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_252));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_240),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_222),
    .B(n_17057),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_255));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_254));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3023 (.A1(n_19850),
    .A2(n_8991),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_21));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_253));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3029 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_249));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3030 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_221),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_248),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3032 (.A(n_22034),
    .B(n_18843),
    .C(n_4541),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_212),
    .B(n_10965),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3034 (.A(n_15217),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_201),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_242));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_225),
    .B(n_10789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_240));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3037 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_239));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_238));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_237));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3040 (.A(n_10789),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_236));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3041 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_235));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3042 (.A(n_8989),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_758));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3043 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_200),
    .A2(n_15218),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_201),
    .B2(n_19783),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_233));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3044 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_173),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_232));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3045 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_170),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_231));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3046 (.A(n_17057),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_185),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3047 (.A(n_26216),
    .B(n_19851),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_229));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3048 (.A(n_19850),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_228));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_224));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3055 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_222));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3056 (.A(n_10964),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3059 (.A(n_8980),
    .B(n_8993),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_218));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_760));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_211),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_212));
 XNOR2x2_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3067 (.A(n_18806),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3068 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_13),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_210));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3069 (.A(n_26111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_136),
    .C(n_19777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_209));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3072 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_197),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_204));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_206));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3075 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_205));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_200));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_199));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_166),
    .B(n_13193),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_19));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_35),
    .C(n_10973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_99),
    .C(n_5643),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_201));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3085 (.A(n_12625),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_18));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_147),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_198));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3088 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106),
    .B(n_19072),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_762));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_180),
    .B(n_18695),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_192));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3091 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3092 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_190));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_197));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3095 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_150),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_133),
    .B(n_12623),
    .C(n_4665),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_186));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_149),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_185));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_35),
    .B(n_10973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_177));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_175));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3114 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_174));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_1),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_139),
    .C(n_3090),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_17));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3116 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_31),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_173));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3123 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3125 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_162));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_170));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_169));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3129 (.B(n_12289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_16),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_66));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3130 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_166),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_101));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_158));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_150));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3138 (.A(n_3090),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_74),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_159));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_44),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_157));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_156));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_155));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_34),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_151));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_146));
 MAJIxp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_63),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_48),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_145));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_81),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_140));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3162 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_12),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3164 (.A(n_12290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_137));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_58),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3168 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_10),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_13));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_764));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_59),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_73),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_126));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3177 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_76),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_10),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3179 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_31),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_122));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_131));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3183 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_117));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_116));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_115));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3186 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_39),
    .A2(n_21798),
    .B1(n_21797),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_114));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3187 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_113));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_121));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3190 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_43),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_110));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3192 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_120));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3193 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_118));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_109));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3196 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_108));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3197 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_107));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3198 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_105));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_104));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_103));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3203 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_101));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3204 (.A(n_12622),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_99));
 AOI22xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3206 (.A1(n_4463),
    .A2(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B1(n_3760),
    .B2(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_98));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_766));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3210 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_89));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_77));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_10));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_73));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3221 (.A(n_3150),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3222 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_94));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_12));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3227 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(n_3760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3228 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_90));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3229 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_88));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3231 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3232 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3239 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_11));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3242 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_68));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3247 (.A(n_2325),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .B(n_3275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(n_6972),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_63));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_59));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3255 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_51));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_42));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_39));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_33));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_62));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_58));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3266 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_57));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3269 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3270 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3271 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3272 (.A(n_21183),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_48));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3274 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_47));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3275 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[7]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3279 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .B(n_3275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3280 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3281 (.A(n_2325),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_36));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3283 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_6973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_34));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_32));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[3]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_31));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3287 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_30));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3288 (.A(n_6973),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_29));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3289 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[5]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_28));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_27));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[2]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[1]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_25));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3296 (.A(n_8992),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_756));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_2));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[4]),
    .B(n_2337),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_122_55_n_0));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1740 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_324),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_298),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_301),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_211),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_768));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1743 (.A(n_15090),
    .B(n_14430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_776));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1744 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_283),
    .A2(n_11739),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_332));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1746 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_298),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_324),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_301),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_330));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1747 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_324),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_293),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_294),
    .B2(n_11739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_774));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1748 (.A(n_14431),
    .B(n_6265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_778));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1751 (.A(n_11739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_324));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_304),
    .B(n_7781),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_782));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1767 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_308),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_309));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_290),
    .B(n_6189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_308));
 NOR2xp33_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1771 (.A(n_5544),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_305));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1772 (.A(n_5048),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_304));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1775 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_281),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_263),
    .B(n_12261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_301));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_786));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_294));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_291));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_298));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1786 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_293));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1788 (.A(n_11418),
    .B(n_6191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_290));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1791 (.A(n_6189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_285));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1794 (.A(n_11423),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_288));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1798 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_282));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_17),
    .B(n_11137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_283));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1800 (.A(n_11137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_281));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1803 (.A(n_13655),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_278));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_265));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1817 (.A(n_7228),
    .B(n_13658),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_266));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1818 (.A(n_13658),
    .B(n_7228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_264));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_263));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1825 (.A1(n_15456),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_215),
    .B1(n_4107),
    .B2(n_15457),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_256));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1833 (.A(n_7227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_249));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1838 (.A(n_11138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_250));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1840 (.A(n_12616),
    .B(n_15097),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_243));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1841 (.A(n_15097),
    .B(n_12616),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_242));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_792));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1843 (.A(n_15213),
    .B(n_13295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_240));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1844 (.A(n_15213),
    .B(n_13295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_226));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1873 (.A(n_19002),
    .B(n_2663),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_224));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1879 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_187),
    .B(n_2744),
    .C(n_2431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_215));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_182),
    .B(n_5890),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_214));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_794));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_11),
    .B(n_5045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_204));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_201));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_199));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_27),
    .B(n_21511),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_197));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1902 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_166),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_85),
    .B2(n_21932),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_195));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1905 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_161),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_30),
    .B1(n_4518),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_190));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_183));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_182));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1920 (.A(n_11729),
    .B(n_5126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_187));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_184));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_66),
    .C(n_22838),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_180));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_168));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1942 (.A(n_21932),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_166));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1943 (.A(n_21932),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_165));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_169));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1951 (.A(n_14237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_112),
    .C(n_14238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_163));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1952 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_33));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1953 (.A(n_15589),
    .B(n_13291),
    .C(n_13289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_32));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1954 (.A(n_15215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_161));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_158));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1959 (.A(n_11821),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1966 (.A(n_15093),
    .B(n_15094),
    .C(n_15092),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_30));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_118),
    .C(n_5894),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_154));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_152));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_796));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_143));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1984 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_23),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_27),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_151));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_66),
    .B(n_22838),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1997 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_115),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_138));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2002 (.A(n_13537),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_128));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_126));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_23),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_27));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_119),
    .B(n_2718),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_123));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_115));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_110));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(n_6576),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_98));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_92));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_43),
    .B(n_3107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2064 (.A(n_14373),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_77),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_78));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_22));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g20805 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_193),
    .Y(n_12261));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_67));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g20830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_96),
    .Y(n_12286));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_56));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_40),
    .B(n_4528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_798));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2094 (.A(n_6576),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2096 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(n_14373),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_48));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2098 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2102 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_77));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2107 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_66));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2111 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_64));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_46),
    .B(n_14372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_47),
    .B(n_3113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_58));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2120 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[15]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_53));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2123 (.A(n_14523),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2124 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_50));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_208),
    .B(n_11138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_17));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_185),
    .B(n_7553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2143 (.A(n_14724),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_11));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g2151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_3));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g21592 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .Y(n_13289));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g21594 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_13291));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g21597 (.A(n_13291),
    .B(n_13289),
    .Y(n_13292));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g22440 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(n_14237));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g22441 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .Y(n_14238));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_n_224),
    .B(n_11133),
    .Y(n_15085));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23145 (.A(n_15086),
    .Y(n_15088));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23149 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[10]),
    .Y(n_15092));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23150 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_15093));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23151 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(n_15094));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23153 (.A(n_15095),
    .B(n_15092),
    .Y(n_15096));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23154 (.A(n_15094),
    .B(n_15093),
    .Y(n_15095));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23155 (.A(n_15096),
    .B(n_14718),
    .Y(n_15098));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g23557 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[11]),
    .B(n_24402),
    .Y(n_15589));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_124_55_g30148 (.A(n_22834),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[8]),
    .Y(n_22838));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1686 (.A1(n_14730),
    .A2(n_4377),
    .B(n_14733),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_189),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_704));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1688 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_708));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1689 (.A(n_19147),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_287),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_712));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1690 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_246),
    .A2(n_14732),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_288));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1691 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_269),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_279),
    .B(n_18698),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_287));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1694 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_271),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_714));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1695 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_716));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1696 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_249),
    .A2(n_16663),
    .B(n_3619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_282));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1699 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_279));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1700 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_268),
    .A2(n_16664),
    .B(n_15181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_278));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_264),
    .B(n_16664),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_718));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1706 (.A(n_26062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_720));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1707 (.A(n_18698),
    .B(n_15173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_271));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1709 (.A(n_15173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_269));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1712 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_249),
    .B(n_15191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_268));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1715 (.A1(n_15179),
    .A2(n_15177),
    .B(n_15191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_265));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1716 (.A(n_3619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_264));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1721 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_234),
    .A2(n_7588),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_28));
 XOR2xp5_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_242),
    .B(n_7589),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_722));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1726 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_257));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1732 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1738 (.A(n_15174),
    .B(n_15175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_245));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_246));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_244));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_243));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_242));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_237));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1752 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_235));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_236));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1754 (.A(n_13641),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_231));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_224),
    .B(n_21630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_234));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1756 (.A(n_21630),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_233));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_232));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1761 (.A(n_8006),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_228));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1764 (.A(n_13640),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_222));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1766 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_184),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_204),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_224));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_216));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_130),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_218));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1776 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_7),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_150),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_217));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_728));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_204));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_169),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_199));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_196));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1804 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_1),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_129),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_194));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1809 (.A(n_5739),
    .B(n_19073),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_730));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_7),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_150),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_184));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1812 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_183));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_182));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_181));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1818 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_180));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1819 (.A(n_16466),
    .B(n_19566),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_177));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1824 (.A(n_19183),
    .B(n_26214),
    .C(n_19768),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_178));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_173));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_172));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1829 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_132),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_81),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_169));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_168));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1831 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_171));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1832 (.A1(one_),
    .A2(n_5739),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_170));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_72),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_167));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1837 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_78),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_164));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1843 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_103),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_128),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_102),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_155));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1844 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_154));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1848 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_160));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_159));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1853 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_153));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1857 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_69),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_150));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_147));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1869 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_141));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1871 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_30),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_49),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_140));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_137));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_19));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_54),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_135));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1885 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_55),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_20));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_98),
    .C(n_15799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1888 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_94),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_131));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1889 (.A(n_14742),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_15),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_34),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_18));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_130));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1891 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_128));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1893 (.A1(n_5738),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_64),
    .B(n_5739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_732));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_124));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1895 (.A1(n_15799),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_83),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_38),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_84),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_122));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_121));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1901 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_129));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_114));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_112));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_118));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_110));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1915 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_90),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_91),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_117));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1916 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_57),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_107));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_106));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_104));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_103));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_17));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_91));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1936 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_81));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1945 (.A(n_16749),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_98));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1947 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(n_16749),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_94));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1951 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_93));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_92));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1953 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1954 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1955 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1957 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_87));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(n_2831),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_78));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1969 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_69));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1974 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_68));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_58));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1981 (.A(n_19567),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_49));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1984 (.A(n_15799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_66));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1987 (.A(n_2544),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_64));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_63));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_59));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_55));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .B(n_16749),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_54));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_50));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_45));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2007 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2012 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_35));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_34));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_33));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[23]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_32));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[21]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_30));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2023 (.A(n_19571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_10));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_7));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2028 (.B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_5),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_0));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2031 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_43),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g2033 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_n_0));
 NAND2x1p5_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_126_55_g23756 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[22]),
    .B(n_16749),
    .Y(n_15799));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g14545 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_32),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_258),
    .Y(n_4771));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g14546 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_16),
    .B(n_10278),
    .Y(n_4772));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g14547 (.A(n_10278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_16),
    .Y(n_4773));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g14551 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_277),
    .A2(n_4777),
    .B(n_4233),
    .Y(n_4778));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g14552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_293),
    .B(n_4777),
    .Y(n_4779));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_288),
    .A2(n_22307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_672));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_226),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_674));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_680));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1709 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_288),
    .A2(n_22307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_315));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1711 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_297),
    .A2(n_12561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_300),
    .B(n_12561),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_682));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1714 (.A(n_22847),
    .B(n_4778),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_684));
 AOI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1720 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_299),
    .A2(n_9008),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_33),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_305));
 NAND3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1721 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_296),
    .B(n_9008),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_304));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1724_dup (.A1(n_4771),
    .A2(n_4772),
    .B(n_4773),
    .Y(n_4777));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_275),
    .B(n_4771),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_688));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1726 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_300));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1727 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_285),
    .A2(n_22846),
    .B(n_22844),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_299));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1728 (.A(n_9008),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_297));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1730 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_277),
    .B(n_22846),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_296));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1731 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_295));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1733 (.A(n_26208),
    .B(n_10416),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_33));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1735 (.A(n_4234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_293));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1736 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_292));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_291));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_268),
    .B(n_3823),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_690));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1745 (.A(n_6373),
    .B(n_12063),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_285));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1747 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_280));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1748 (.A(n_2694),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_692));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_274),
    .B(n_4772),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_275));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_265),
    .B(n_20143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_279));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1752 (.A(n_20143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_278));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1753 (.A(n_12063),
    .B(n_6373),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_277));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1754 (.A(n_4773),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_274));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_269));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_268));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_14),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_270));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_265));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1767 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_247),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_261));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1770 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_694));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_260));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1773 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_190),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_254));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1782 (.A(n_13125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1784 (.A(n_13125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_247));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1786 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_227),
    .A2(n_18904),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_31));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1787 (.A(n_10280),
    .B(n_18144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1792 (.A(n_11095),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_243));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1794 (.A(n_8265),
    .B(n_18904),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_241));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1795 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_240));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_696));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_216),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_154),
    .C(n_2891),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_231));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1807 (.A(n_8265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_230));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_226));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1814 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_196),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_227));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1815 (.A(n_11097),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_30));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_224));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_197),
    .B(n_6444),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_223));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_123),
    .B(n_19075),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_698));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_211));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1840 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_210));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_215));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1848 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_173),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_186),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_172),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_202));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1849 (.A(n_6444),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_201));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_166),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_122),
    .B(n_10009),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1856 (.A(n_10009),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_198));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_145),
    .B(n_11446),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_197));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1860 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_196));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1864 (.A1(n_9577),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_165),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_162),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1868 (.A(n_11446),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_190));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_186));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_184));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_138),
    .B(n_10005),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_180));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_177));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_99),
    .B(n_11098),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1896 (.A(n_19559),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_172));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_166));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1902 (.A(n_9577),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_163));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1903 (.A(n_9577),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_162));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_165));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1924 (.A(n_19446),
    .B(n_19447),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_154));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_149));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_700));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_144));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_150));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1937 (.A1(n_9576),
    .A2(n_9573),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_110),
    .B2(n_9574),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_141));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_148));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_135));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_133));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_130));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_128));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_127));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_46),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_132));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_119));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_118));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_116));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_114),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1971 (.A(n_9576),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_94));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_79));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(n_14981),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .B(n_2944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(n_14984),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_14183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(n_14981),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(n_14186),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_2392),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(n_14987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_78));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2014 (.A(n_2381),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[31]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .B(n_14987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_50));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[30]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_45));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[24]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_39));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[29]),
    .B(n_3504),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2063 (.A(n_14183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[27]),
    .B(n_14183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_35));
 BUFx2_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2069 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_34));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2071 (.A(n_19129),
    .B(n_12069),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_16));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_211),
    .B(n_11095),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2075 (.A(n_3990),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_115),
    .B(n_5536),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_9));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g2085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g30151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_n_207),
    .B(n_19181),
    .Y(n_22841));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g30152 (.A(n_12066),
    .B(n_22843),
    .Y(n_22844));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g30153 (.B(n_22842),
    .Y(n_22843),
    .A(n_22841));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g30155 (.A1(n_22845),
    .A2(n_12066),
    .B(n_22846),
    .Y(n_22847));
 NOR2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_128_55_g30157 (.A(n_12066),
    .B(n_22843),
    .Y(n_22846));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_297),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_654));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g25535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_239),
    .Y(n_4349));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g25536 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_226),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_249));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g25537 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_239),
    .Y(n_17669));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g25538 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_271),
    .B(n_17670),
    .Y(n_17672));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_223),
    .B(n_22969),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_642));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2960 (.A(n_19039),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_648));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2964 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_29),
    .A2(n_13130),
    .B(n_22082),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_315));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_298),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_652));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2970 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_302),
    .A2(n_17673),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_306),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_29));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2971 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_282),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_312));
 OAI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2973 (.A1(n_13130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_305),
    .A3(n_14925),
    .B1(n_14925),
    .B2(n_22079),
    .C(n_14921),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_311));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_302),
    .B(n_17673),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_310));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2975 (.A(n_19219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_656));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2976 (.A(n_14925),
    .B(n_13130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_308));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_306));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2979 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_289),
    .A2(n_7283),
    .B(n_7282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_305));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2981 (.A(n_17673),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_304));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_282),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_302));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2989 (.A(n_7283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_298));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_297));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2992 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_295));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2993 (.A1(n_8639),
    .A2(n_17670),
    .B(n_8640),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_294));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_291));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2996 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_290));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2997 (.A(n_7282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_288));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g2998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_262),
    .B(n_14382),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_286));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3001 (.A(n_22820),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_289));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_660));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3008 (.A(n_22820),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_282));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_274));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_272));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3013 (.A(n_8625),
    .B(n_8639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_271));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3016 (.A(n_19235),
    .B(n_14928),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_275));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3019 (.A(n_3833),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_219),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_270));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3025 (.A(n_10102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_264));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_263));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3027 (.A(n_26177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_262));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3028 (.A(n_26177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_261));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_252),
    .B(n_4349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_662));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3038 (.A(n_17669),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_252));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_10),
    .B(n_7223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_242));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_664));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_239));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_235));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3055 (.A(n_9631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_238));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3058 (.A(n_4138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_149),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_234));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3060 (.A(n_10356),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_184),
    .C(n_15355),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_232));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_228));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_226));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_229));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_227));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_223));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3069 (.A1(n_4429),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_225));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_220));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3080 (.A(n_19440),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_113),
    .C(n_9799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120),
    .B(n_19076),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_666));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_215));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_119),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3101 (.A(n_9633),
    .B(n_9632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_201));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_205));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3105 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_200));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_199));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_161),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_45),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_193));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3120 (.A(n_10360),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_182));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_176));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_49),
    .B(n_10099),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_183));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_73),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_175));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3135 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_76),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_166));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_172));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3144 (.A(n_3882),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_167));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_161),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_162));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_156));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_164));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_101),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_161));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_19),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_34),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_155));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_64),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_154));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_21));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3172 (.A(n_21937),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_142));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_668));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_136));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3181 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_90),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_17),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_127));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3189 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_40),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_57),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_126));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_133));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3192 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_19),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_34),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_124));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3196 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_100),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_131));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_105),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_53),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_54),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_121));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_120));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_118));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3208 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_115));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3209 (.A(n_21936),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_114));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .A2(n_3168),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B2(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_107));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_105));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_102));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_19));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_92));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_90));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_86));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_77));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_74));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_108));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_103));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3239 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(n_6861),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_99));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3242 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3245 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3247 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3249 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3252 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_85));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3253 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3254 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(n_22743),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_83));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3260 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B(n_15192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3263 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_17));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_73));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_670));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_64));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_54));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_48));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_45));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_41));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_34));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3283 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B(n_3168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_70));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_69));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_65));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3289 (.A(n_15192),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3290 (.A(n_3181),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_59));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3293 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3297 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_51));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_49));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3304 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3306 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[32]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_42));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3307 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[35]),
    .B(n_6861),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[38]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_38));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3310 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3311 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[33]),
    .B(n_18041),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[36]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3313 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[34]),
    .B(n_4831),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_7),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3323 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_9));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_116),
    .B(n_21937),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3331 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_g3332 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[37]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_130_55_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_299),
    .B(n_9956),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_622));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22016 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_16772),
    .Y(n_13772));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22017 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(n_16772),
    .Y(n_13773));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22018 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(n_16763),
    .Y(n_13774));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22022 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(n_16763),
    .Y(n_13778));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22023 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .Y(n_13779));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22029 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(n_16769),
    .Y(n_13785));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g22039 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .Y(n_13795));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_225),
    .B(n_9805),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_610));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_298),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_616));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2963 (.A(n_7107),
    .B(n_22431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_614));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2964 (.A1(n_9957),
    .A2(n_9960),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_317));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2966 (.A(n_8391),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_620));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2971 (.A1(n_9956),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_284),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_314));
 OAI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2973 (.A1(n_9959),
    .A2(n_9697),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285),
    .B2(n_9961),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_282),
    .B(n_14944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_624));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285),
    .B(n_9959),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_310));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_303),
    .B(n_9960),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_309));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_303));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2987 (.A(n_9961),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_302));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_299));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2991 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_270),
    .A2(n_14415),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_298));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_293));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2996 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_292));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g2997 (.A(n_8392),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g29970 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .Y(n_22623));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g29972 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .Y(n_22625));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g29974 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B(n_22616),
    .Y(n_13133));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g29982 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(n_22616),
    .Y(n_22635));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3001 (.A(n_11127),
    .B(n_13040),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_291));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_280),
    .B(n_11124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_282));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3006 (.A(n_14415),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_281));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3007 (.A(n_14415),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_285));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3008 (.A(n_13040),
    .B(n_11127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_284));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3009 (.A(n_11126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_280));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_235),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_270));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3023 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_224),
    .C(n_4012),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_265));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3027 (.A(n_19077),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3028 (.A(n_19077),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3034 (.A(n_22428),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_630));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3037 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_235),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_188),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_226),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_249));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3045 (.A(n_14394),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_247));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_226),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_244));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3049 (.A(n_11389),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_243));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_632));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_237));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3058 (.A(n_18795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_147),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_236));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3059 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_187),
    .B(n_3562),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_235));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3062 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_202),
    .B(n_14418),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_232));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_230));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3064 (.A(n_22427),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_228));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_231));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_229));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_70),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_191),
    .B(n_9806),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_225));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_226));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3076 (.A(n_21524),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_5),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_223));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_44),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_220));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3082 (.A(n_9297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118),
    .B(n_19078),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_634));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3086 (.A(n_13142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_214));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_211));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_210));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3092 (.A(n_9298),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_207));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3097 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_201));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3101 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_5),
    .B(n_21524),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_199));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_149),
    .B(n_14645),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_202));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3105 (.A(n_22426),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3109 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_144),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_142),
    .B1(n_14645),
    .B2(n_11411),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_194));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_159),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_43),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_193));
 AOI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3111 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_152),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_111),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_22),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_191));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3115 (.A(n_10915),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_114),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3116 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_187));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3120 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_180));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_176));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_183));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3128 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3134 (.A(n_22422),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_71),
    .C(n_13133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_173));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3138 (.A(n_22635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_170));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_61),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_169));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3143 (.A(n_13778),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3144 (.A(n_3210),
    .B(n_18702),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_165));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_160));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_158));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_162));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_92),
    .B(n_13785),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_62),
    .C(n_13774),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_153));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3158 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3159 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_148));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3161 (.A(n_11411),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3163 (.A(n_22625),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_47),
    .C(n_13773),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_80),
    .B(n_9628),
    .C(n_14388),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_150));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3166 (.A(n_21929),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3167 (.A(n_13795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_106),
    .C(n_22635),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3168 (.A(n_22623),
    .B(n_13778),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_145));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3171 (.A(n_14645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_142));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_140));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_636));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3176 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3179 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_92),
    .B1(n_13785),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_134));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3182 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_46),
    .B1(n_13773),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_132));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_139));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3187 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3188 (.A(n_13795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_131));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_101),
    .B(n_22623),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_121));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_103),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_51),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_52),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_128));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_126));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_60),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_119));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_118));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_117));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_114));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3208 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_113));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3209 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_112));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_110));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .A2(n_18049),
    .B1(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B2(n_23276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_108));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_105));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3216 (.A(n_13785),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_92));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_97));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3242 (.A(n_3309),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3247 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(n_14674),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_89));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(n_3713),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3256 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_3709),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_71));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_638));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3266 (.A(n_13773),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_64));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_62));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_43));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3282 (.A(n_13779),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_32));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3283 (.A(n_19396),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[40]),
    .B(n_18049),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_68));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_67));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3289 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_61));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[41]),
    .B(n_23280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(n_19393),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[42]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[45]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[43]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[46]),
    .B(n_19395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_36));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3310 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[44]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_7),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_114),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_8));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3325 (.A(n_15158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_7));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_4),
    .B(n_22625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_5));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_g3331 (.A(n_13774),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_132_55_n_1));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14553 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_32),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_258),
    .Y(n_4780));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14555 (.A(n_10094),
    .B(n_5583),
    .Y(n_4782));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14556 (.A(n_4783),
    .Y(n_4784));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14557 (.A1(n_4780),
    .A2(n_5584),
    .B(n_4782),
    .Y(n_4783));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14559 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_277),
    .A2(n_4786),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_285),
    .Y(n_4787));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g14560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_293),
    .B(n_4786),
    .Y(n_4788));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_576));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1707 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_269),
    .B(n_14335),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_580));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1708 (.A(n_19240),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_584));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1709 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_315));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1711 (.A1(n_24979),
    .A2(n_6401),
    .B(n_6406),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_313));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1712 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_287),
    .B2(n_14336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_582));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1713 (.A(n_6404),
    .B(n_6401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_586));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1716 (.A(n_14336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_307));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1724_dup (.A1(n_4780),
    .A2(n_5584),
    .B(n_4782),
    .Y(n_4786));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_275),
    .B(n_4780),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_592));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1735 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_284),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_293));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_291));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_268),
    .B(n_3901),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_594));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_287));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_284));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_286));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1745 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_285));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1748 (.A(n_2793),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_596));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_274),
    .B(n_5584),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_275));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_277));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1754 (.A(n_4782),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_274));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_271));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_269));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_268));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_14),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_270));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1763 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_239),
    .B(n_19661),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_266));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_265));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1765 (.A(n_19667),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_264));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1767 (.A1(n_11310),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_31),
    .B(n_11309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_261));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1770 (.A(n_21928),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_598));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_246),
    .B(n_7974),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_243),
    .B(n_19079),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_260));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1773 (.A(n_7974),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1774 (.A(n_11309),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1775 (.A(n_19079),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_190),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_254));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_236),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_26),
    .C(n_23376),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_253));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1780 (.A(n_19667),
    .B(n_11743),
    .C(n_14208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_252));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1781 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_237),
    .B(n_13331),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_251));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1783 (.A(n_11310),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_248));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1786 (.A1(n_21927),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_13),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_31));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1787 (.A(n_26073),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_246));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1790 (.A1(n_11743),
    .A2(n_23685),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_222),
    .B2(n_14208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_243));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_238));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1799 (.A(n_5131),
    .B(n_11145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_237));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_207),
    .B(n_10739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_236));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_600));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1804 (.A(n_19662),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_233));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_3),
    .B(n_18809),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_228));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_30));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1819 (.A(n_11743),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_222));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1825 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_26));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_225));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1831 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_188),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_123),
    .B(n_19080),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_602));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_211));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_181),
    .B(n_9694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_201));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1850 (.A(n_9694),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_208));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_148),
    .C(n_14203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1854 (.A(n_21926),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_122),
    .B(n_10212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_200));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_195));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_197));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1860 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_196));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_190));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1875 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_121),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_134),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_120),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_181));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_51),
    .B(n_16063),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_188));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_184));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_138),
    .B(n_10208),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_180));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_172));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_166));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1906 (.A(n_13685),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_21),
    .C(n_22884),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_165));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_158));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_99),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_22));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_46),
    .B(n_22868),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_104),
    .C(n_9692),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_154));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1925 (.A(n_16062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_51),
    .C(n_22873),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_153));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_604));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1930 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_68),
    .A2(n_22885),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_69),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_146));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_144));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1933 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_78),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_79),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_143));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_148));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_135));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_127));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_126));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_46),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_132));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_124));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_93));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_88));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_79));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(n_2930),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(n_3592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(n_2377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_2711),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_89));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_78));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2014 (.A(n_2697),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_46));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2032 (.A(n_22885),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[55]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(n_3479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_45));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[48]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_40));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2065 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .B(n_22865),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_35));
 BUFx2_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2069 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_14));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_9));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2079 (.A(n_19172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_8));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_4));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2084 (.A(n_22868),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_3));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g2087 (.A(n_2927),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[51]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_0));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g21633 (.A(n_10299),
    .Y(n_13331));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g30178 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22868));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g30189 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(n_22880),
    .Y(n_22881));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g30194 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22884));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g30195 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22885));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g31873 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_34),
    .B(n_2927),
    .Y(n_24751));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g31874 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[50]),
    .B(n_3468),
    .Y(n_24752));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g31875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_n_35),
    .B(n_24753),
    .Y(n_24754));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_134_55_g31876 (.A(n_24752),
    .B(n_24751),
    .Y(n_24753));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g14652 (.A(n_13717),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_20),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_81),
    .Y(n_4902));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g14653 (.A(n_10283),
    .Y(n_4906));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g14655 (.A(n_4903),
    .B(n_4902),
    .Y(n_4904));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g14657 (.A(n_20017),
    .B(n_10283),
    .Y(n_4907));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_546));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1743 (.A(n_6787),
    .B(n_7980),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_552));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1746 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_298),
    .A2(n_11235),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_301),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_330));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1759 (.A(n_10585),
    .B(n_10582),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_560));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1769 (.A(n_19959),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_307));
 NOR2xp33_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_297),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_305));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1772 (.A(n_8696),
    .B(n_8691),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_304));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1775 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_281),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_301));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_562));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1778 (.A(n_8694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_296));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_294));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_291));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_298));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1784 (.A(n_14162),
    .B(n_9510),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_297));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1786 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_293));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1788 (.A(n_14162),
    .B(n_9510),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_290));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1798 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_282));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_17),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_283));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_281));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1801 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_278));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1804 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_252),
    .A2(n_9255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_277));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1808 (.A(n_6100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_273));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_269),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_270));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1812 (.A(n_4451),
    .B(n_4810),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_269));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_255),
    .B(n_14907),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_266));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1818 (.A(n_14907),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_264));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1820 (.A(n_2893),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_566));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1823 (.A(n_6100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_190),
    .C(n_3983),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_259));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1825 (.A1(n_4451),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_215),
    .B1(n_4810),
    .B2(n_6097),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_256));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_253));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_12),
    .B(n_20018),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_255));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1829 (.A(n_6771),
    .B(n_14908),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_254));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1830 (.A(n_6771),
    .B(n_14908),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_252));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_190),
    .B(n_10014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_247));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1838 (.A(n_10013),
    .B(n_14159),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_250));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_568));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1843 (.A(n_4906),
    .B(n_20017),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_240));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1844 (.A(n_4906),
    .B(n_20017),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_239));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_229),
    .B(n_9253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_238));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1849 (.A(n_13358),
    .B(n_9712),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_29),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_235));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1854 (.A(n_9254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_197),
    .B(n_5842),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_226));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1879 (.A(n_5842),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_27),
    .C(n_3436),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_215));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_210));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1886 (.A(n_14159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_129),
    .B(n_26178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_570));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_201));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_199));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_27),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_31),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_197));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1902 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_166),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_85),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_195));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_198));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_193));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1908 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_149),
    .B(n_13149),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1910 (.A(n_13149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_190));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_182));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_184));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_66),
    .C(n_13227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_180));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1940 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_135),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_171));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1942 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_166));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1949 (.A(n_13248),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_108),
    .C(n_11826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_160));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_158));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1959 (.A(n_5549),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_157));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1960 (.A(n_5549),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_156));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_113),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_31));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_26),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_30));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_126),
    .B(n_9638),
    .C(n_9639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_29));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_152));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_572));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_143));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1984 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_23),
    .A2(n_13243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_27),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_151));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_66),
    .B(n_13227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1994 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_96),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_114),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_135));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1997 (.A1(n_13238),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_138));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2 (.A(n_9256),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_564));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2002 (.A(n_13244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_128));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2010 (.A(n_13242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_126));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_23),
    .B(n_13243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_27));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_119),
    .B(n_12134),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2015 (.A(n_13238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_114));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_102));
 INVx2_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_97));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2026 (.A(n_13718),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_95));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_2657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_117));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_113));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_111));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_110));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_11770),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2054 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_98));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_67));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2086 (.A(n_5548),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_61));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_40),
    .B(n_2747),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_n_574));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2094 (.A(n_2820),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2099 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2107 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(n_3375),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2116 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_47),
    .B(n_4555),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2121 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_53));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2126 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_208),
    .B(n_10013),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_17));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_185),
    .B(n_14912),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_12));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_126),
    .B(n_9637),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2150 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_81),
    .B(n_13717),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_3));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21528 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_3528),
    .Y(n_13227));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21539 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(n_13231),
    .Y(n_13238));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_0));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21543 (.A(n_13231),
    .B(u_NV_NVDLA_cmac_u_core_wt0_actv_data[62]),
    .Y(n_13242));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21544 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[63]),
    .B(n_13231),
    .Y(n_13243));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21545 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(n_13231),
    .Y(n_13244));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21549 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_2657),
    .Y(n_13248));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21961 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(n_13707),
    .Y(n_13717));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21962 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[58]),
    .B(n_13707),
    .Y(n_13718));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g21971 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[57]),
    .B(n_3528),
    .Y(n_13727));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g22087 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[59]),
    .B(n_11770),
    .Y(n_13843));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g22088 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[60]),
    .B(n_13707),
    .Y(n_13844));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g22089 (.A(u_NV_NVDLA_cmac_u_core_wt0_actv_data[56]),
    .B(n_22019),
    .Y(n_13845));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g22092 (.A(n_13845),
    .B(n_13844),
    .Y(n_13846));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_g26369 (.A(u_NV_NVDLA_cmac_u_core_u_mac_0_mul_136_55_n_305),
    .B(n_11242),
    .Y(n_18578));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1_reg (.CLK(nvdla_core_clk),
    .D(n_17870),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d1));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2_reg (.CLK(nvdla_core_clk),
    .D(n_7),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d2));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_0_pp_pvld_d0_d3_reg (.CLK(nvdla_core_clk),
    .D(n_13),
    .QN(u_NV_NVDLA_cmac_u_core_out_mask[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_4417),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[0]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1238),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[10]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1237),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[11]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1236),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[12]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_17775),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[13]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_16616),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[14]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_22971),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[15]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_10054),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[16]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_20291),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[17]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_20071),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1249),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1247),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1246),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1245),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1243),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1242),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[6]));
 DFFHQNx1_ASAP7_75t_L \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1241),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1240),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[8]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_17873),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1230),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1217),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1216),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1215),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1214),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1213),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1212),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1211),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1210),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1209),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1229),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1228),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_855),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1226),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1224),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1222),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1221),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1220),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1218),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d2[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1208),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1197),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1196),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1195),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1194),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1193),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1192),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1191),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1190),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1189),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1207),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1206),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1205),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1204),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1203),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1202),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1201),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1200),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_0_sum_out_d0_d3_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1199),
    .QN(u_NV_NVDLA_cmac_u_core_out_data0[9]));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g2 (.A(n_22326),
    .B(n_23266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_180));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g24190 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_447),
    .B(n_10515),
    .Y(n_16255));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g24452 (.A(n_23895),
    .B(n_16561),
    .Y(n_16528));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g24463 (.A(n_21278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_494),
    .Y(n_16540));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g25530 (.A(n_17663),
    .Y(n_17665));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g30204 (.A1(n_13667),
    .A2(n_22889),
    .B1(n_6673),
    .B2(n_22894),
    .Y(n_22895));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g30205 (.A(n_22889),
    .Y(n_22894));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6015 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_466),
    .A2(n_16253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_473),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_496));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6017 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_488),
    .A2(n_23753),
    .B(n_20742),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_494));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6023 (.A(n_22323),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_488));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6029 (.A(n_23894),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_439),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_178));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_481),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_438),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_177));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_481));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6035 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_480));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6036 (.A(n_3212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_450),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_176));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_472),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_64));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_472),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_175));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6044 (.A1(n_7407),
    .A2(n_15153),
    .B(n_7408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_473));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6045 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_386),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_383),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_472));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_174));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6049 (.A(n_7408),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_455),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_468));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6051 (.A(n_10515),
    .B(n_7407),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_466));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6057 (.A(n_7407),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_455));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_453));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_432),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_450));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_430),
    .B(n_4365),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_449));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6070 (.A(n_15153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_447));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6071 (.A(n_10515),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_445));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_173));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6075 (.A(n_17665),
    .B(n_24166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_439));
 NAND2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6076 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_412),
    .B(n_24153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_438));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_379),
    .B(n_7410),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_437));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6082 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_381),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_443));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_432));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6085 (.A(n_8196),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_430));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_433));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6095 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_431));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6101 (.A(n_9972),
    .B(n_20023),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_62));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6107 (.A(n_21434),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_412));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_380),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_172));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6125 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_397));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_386),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_384),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_396));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_401));
 XOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6128 (.A(n_9111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_400),
    .B(n_22045));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6130 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_356),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_398));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6132 (.A(n_21134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_347),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_395));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_383),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_384));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_345),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_171));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_353),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_360),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_386));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_385));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_381));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6145 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_380));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_353),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_360),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_383));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_308),
    .B(n_6687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_379));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_342),
    .B(n_21372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_377));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6157 (.A(n_8928),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_372));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_356));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6169 (.A1(n_20794),
    .A2(n_8928),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_354));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_361));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_328),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_360));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_359));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_358));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_325),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_353));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6180 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_291),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .B2(n_12839),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_347));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_352));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6183 (.A1(n_26179),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_345));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_344));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6187 (.A(n_14299),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_299),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_342));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6196 (.A(n_8928),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_330));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_337));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_328));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6201 (.A(n_26179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_327));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_326));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6203 (.A(n_26179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_336));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6208 (.A(n_7311),
    .B(n_21669),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_58));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6213 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_325));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6214 (.A(n_20794),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_322));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6219 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_314));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_308));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_324));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .B(n_26126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_318));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6231 (.A(n_21131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .C(n_15651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_317));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6233 (.A(n_21947),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_315));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6234 (.A(n_19149),
    .B(n_8923),
    .C(n_8929),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_312));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6242 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_300));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6243 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_307));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6245 (.A1(n_10235),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .B1(n_13702),
    .B2(n_4246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_299));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6251 (.A(n_11832),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_298));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6255 (.A(n_12839),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_291));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6264 (.A(n_26079),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_292));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6266 (.A(n_21129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_289));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6272 (.A1(n_6673),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_281));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6274 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_217),
    .B(n_22895),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_279));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6278 (.A(n_13667),
    .B(n_21439),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_278));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6279 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_225),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .B2(n_15740),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_277));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_283));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6289 (.A(n_7311),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_267));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6290 (.A(n_21370),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_265));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_263));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6303 (.A(n_17024),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_126),
    .C(n_11913),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_262));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6304 (.A(n_19084),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .C(n_26181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_261));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6305 (.A(n_26180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_260));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6306 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_259));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6307 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_216),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_258));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6309 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_250));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_251));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_145),
    .B(n_21945),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_240));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_237));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6337 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_233));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6338 (.A(n_11105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_231));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_229));
 AOI21xp5_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6350 (.A1(n_22894),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_84),
    .B(n_21438),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6351 (.A(n_11833),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_232));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6353 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_697),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_228));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6354 (.A(n_20796),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_227));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6356 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6362 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_221));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6364 (.B(n_21152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .A(n_9370));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6365 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_218));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_216));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6374 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6376 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_204));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6379 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6380 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_215));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6382 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_661),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_629),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_213));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6383 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_156),
    .B(n_17587),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_212));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6388 (.A(n_14340),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_643),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_42));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6389 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_209));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_148),
    .B(n_5806),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_207));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6391 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_152),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_655),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_623),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_206));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6392 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_649),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_205));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6396 (.A(n_26079),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6405 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_200));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6412 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_663),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_699),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_190));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_633),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_185));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6419 (.A(n_12571),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_178));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6426 (.A(n_20833),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_162));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6428 (.A(n_20833),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6430 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_797),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6439 (.A(n_9735),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6441 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_168));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6444 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_729),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_165));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6447 (.A(n_23423),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_157));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6448 (.A(n_21152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_156));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6450 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_152));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6451 (.A(n_22180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_601),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_88),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_161));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6459 (.A(n_19058),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_767),
    .C(n_19057),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6463 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_785),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_721),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6465 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_563),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_787),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_723),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6466 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_733),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_637),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_797),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6467 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_691),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_145));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_639),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_671),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_143));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6472 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_743),
    .B(n_12540),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_583),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6474 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_135));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_131));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6477 (.A(n_20796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_129));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6493 (.A(n_14758),
    .B(n_14759),
    .C(n_14761),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6494 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_701),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6495 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_559),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_783),
    .C(n_9728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_793),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_729),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_130));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6499 (.A(n_13960),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_751),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_126));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6500 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_695),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_663),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_125));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_761),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_665),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_633),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_123));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_763),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_635),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_667),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_122));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_603),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_731),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_n_699),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_121));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_597),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_693),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_111));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6514 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_761),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_109));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_791),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_695),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_108));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_667),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_763),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_107));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_106));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6525 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_623),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_655),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_103));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6530 (.A(n_19059),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_575),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_115));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_565),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_98));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6544 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_629),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_661),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_97));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6545 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_731),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_96));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_637),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_733),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_91));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6553 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_90));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_691),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_89));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6556 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_571),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_102));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_795),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_575),
    .B(n_19059),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6561 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_73),
    .B(n_26252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_84));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6562 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_651),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_82));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6585 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_609),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_73));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6586 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_617),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_72));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6588 (.A(n_10595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_71));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6596 (.A(n_19264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_70));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6621 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_34));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6627 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_212),
    .B(n_5627),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_28));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6628 (.A(n_23670),
    .B(n_6411),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_27));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6629 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_26));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6630 (.A(n_26180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_25));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6631 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_140),
    .B(n_7821),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_24));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6632 (.A(n_8495),
    .B(n_21051),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_23));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6637 (.A(n_23668),
    .B(n_23666),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_18));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6642 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_13),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_619));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6647 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_785),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_561),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6649 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_n_787),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_n_563),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_g6650 (.A(n_12987),
    .B(n_12986),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_csa_tree_ADD_TC_OP_6_groupi_n_5));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g14720 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_69),
    .Y(n_4970));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_285),
    .B(n_10429),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_746));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g20807 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_6965),
    .Y(n_12263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_299),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_740));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2963 (.A1(n_12395),
    .A2(n_10318),
    .B(n_12382),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_299));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2964 (.A1(n_3795),
    .A2(n_10429),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_298));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_748));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2969 (.A1(n_13481),
    .A2(n_9388),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_294));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2975 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_274),
    .A2(n_21364),
    .B1(n_13482),
    .B2(n_9388),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_750));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2980 (.A(n_21368),
    .B(n_21362),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_752));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_277),
    .B(n_3796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_285));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_282));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2989 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_245),
    .B(n_10650),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_23));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_277));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2992 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_245),
    .B(n_10650),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_276));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2993 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_275));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g2994 (.A(n_13482),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_274));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3000 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_241),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_22));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_754));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_265));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_262));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3007 (.A(n_12382),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3009 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_261));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_257));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_256));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3015 (.A(n_21289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_259));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_230),
    .B(n_13480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_258));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3018 (.A(n_12395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_252));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_240),
    .B(n_12383),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_222),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_255));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3023 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_226),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_21));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_247));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_244));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3029 (.A(n_10865),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_249));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3031 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_213),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_213),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_20),
    .C(n_8131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_203),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_243));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_237));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_236));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3041 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_235));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3042 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_207),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_758));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3044 (.A(n_10865),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_173),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_232));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3045 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_170),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_231));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_4),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_185),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_216),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_229));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_228));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3049 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_216),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_227));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3051 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_207),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_161),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_224));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3055 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_222));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_203),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_221));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3057 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_20),
    .B(n_8131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_220));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3059 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_218));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_760));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_189),
    .B(n_19462),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_216));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3065 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_213));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3066 (.A(n_20114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_212));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3068 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_186),
    .B(n_19165),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_210));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_132),
    .C(n_3944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_208));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3073 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_179),
    .A2(n_19700),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_207));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_206));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3075 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3076 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_169),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_20));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_200));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_199));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_142),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_203));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_99),
    .C(n_4474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_201));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_18));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_147),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_198));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3087 (.A(n_19462),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_196));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3088 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106),
    .B(n_19085),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_762));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_192));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3091 (.A(n_12387),
    .B(n_12388),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3092 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_190));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_188));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3099 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_187));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3102 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_129),
    .C(n_4017),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_186));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_149),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_185));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3104 (.A(n_19700),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_182));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3105 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_179));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3107 (.A(n_19699),
    .B(n_19701),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_177));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_99),
    .A2(n_8134),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_100),
    .B2(n_4474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_176));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3113 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_130),
    .A2(n_4017),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_134),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_171));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3114 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_174));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_1),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_139),
    .C(n_2685),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_17));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3116 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_31),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_173));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_172));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3121 (.A(n_9750),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_167));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3123 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3125 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_162));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_170));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_169));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3128 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_30),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_168));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3129 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_16),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_66));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_158));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3136 (.A(n_21045),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_29),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_161));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3138 (.A(n_2685),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_74),
    .C(n_25976),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_159));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_44),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_157));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_156));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_155));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_154));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_153));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_146));
 MAJIxp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_63),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_48),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_145));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_27),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_56),
    .C(n_4970),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_141));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_81),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_140));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3162 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_12),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_37),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_137));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3166 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_30),
    .C(n_12262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3168 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_67),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_764));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_59),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_73),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_126));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3175 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_37),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_125));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3179 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_31),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_122));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_131));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_129));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3183 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_117));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_116));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_115));
 OAI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3186 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_39),
    .A2(n_12263),
    .B1(n_12262),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_114));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3187 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_26),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_113));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_121));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3189 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_112));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3190 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_43),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_110));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3193 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_118));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3195 (.A(n_21043),
    .B(n_21044),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_109));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3196 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_92),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_108));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3198 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_106));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_103));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_102));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_99));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_100));
 AOI22xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3206 (.A1(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .A2(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B1(n_3761),
    .B2(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_98));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_766));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3210 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_89));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3222 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_12));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3227 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B(n_3760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3228 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_90));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3229 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_88));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3231 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B(n_3275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3232 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3242 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3245 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_6972),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_68));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3247 (.A(n_2325),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_67));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(n_3275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(n_6972),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_59));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3255 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_51));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_42));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_39));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_37));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_33));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_58));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3266 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_57));
 NAND2x1p5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3267 (.A(n_2335),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3269 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3271 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_48));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3274 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_47));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3275 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[7]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3279 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3280 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3281 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(n_2335),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_36));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3283 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_35));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_32));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[3]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_31));
 NAND2x1p5_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3287 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_30));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[0]),
    .B(n_6973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_29));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3289 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[5]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_28));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_27));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[2]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[1]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_25));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3295 (.A(n_21289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_226),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_756));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3297 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_168),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_16),
    .B(n_19165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3299 (.A(n_3443),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_4));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[4]),
    .B(n_2337),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_122_55_n_0));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g14605 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(n_14523),
    .Y(n_4856));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g14718 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_101),
    .Y(n_4968));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_225),
    .B(n_19265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_770));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1743 (.A(n_26045),
    .B(n_22334),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_776));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1748 (.A(n_22332),
    .B(n_21527),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_778));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1749 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_305),
    .B(n_12110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_780));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_304),
    .B(n_13694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_782));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1767 (.A(n_21837),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_309));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1771 (.A(n_21846),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_305));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1772 (.A(n_21845),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_304));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_786));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1778 (.A(n_21828),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_296));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1780 (.A(n_21845),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_292));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1782 (.A(n_21835),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_291));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1791 (.A(n_21836),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_285));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1801 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_278));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1804 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_252),
    .A2(n_9884),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_277));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_233),
    .B(n_6940),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_275));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_255),
    .B(n_6930),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_266));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1818 (.A(n_6930),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_264));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1820 (.A(n_22041),
    .B(n_19086),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_790));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1823 (.A(n_19273),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_190),
    .C(n_3011),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_259));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1824 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_233),
    .A2(n_6942),
    .B(n_6941),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_258));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_253));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_12),
    .B(n_3279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_255));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1829 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_207),
    .B(n_6926),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_254));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_207),
    .B(n_6926),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_252));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_249));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_190),
    .B(n_10159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_247));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1838 (.A(n_20074),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_250));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1839 (.A(n_3279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_185),
    .C(n_20152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_248));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1840 (.A(n_9603),
    .B(n_9604),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_243));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1841 (.A(n_9604),
    .B(n_9603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_242));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_792));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_14),
    .B(n_10612),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_234));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1852 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_233));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_225));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_210));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_134),
    .B(n_20148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_212));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1888 (.A(n_22005),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_794));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1893 (.A(n_21211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_131),
    .C(n_21206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1897 (.A(n_22040),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_201));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_198));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1910 (.A(n_6579),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_190));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_184));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_180));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1939 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_172));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_168));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_169));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_167));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1952 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_33));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_26),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_30));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_118),
    .C(n_15324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_154));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_796));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_149));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1977 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_56),
    .A2(n_15325),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_104),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_148));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_143));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1994 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_113),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_96),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_114),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_135));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1997 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_115),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_138));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_262),
    .B(n_9885),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_788));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_134));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_128));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_127));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_126));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_119),
    .B(n_2718),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_114));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_97));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_123));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_113));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_112));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_110));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2054 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_98));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2062 (.A(n_14523),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_90));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(n_4275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_24));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2064 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2065 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(n_14523),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_67));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_56));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_40),
    .B(n_4528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_798));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2094 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2096 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_48));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2098 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2099 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .B(n_6576),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2102 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_77));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_73));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2105 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2116 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[12]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_47),
    .B(n_3113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_57));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2120 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2121 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[15]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_208),
    .B(n_20074),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_17));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_172),
    .B(n_8948),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_15));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_9),
    .B(n_7805),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_185),
    .B(n_20152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_112),
    .B(n_13324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g23553 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[13]),
    .Y(n_15585));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g31527 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_81),
    .B(n_24403),
    .Y(n_24404));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g31528 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[11]),
    .Y(n_24403));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_g31529 (.A(n_24403),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_20),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_124_55_n_81),
    .Y(n_24405));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g14537 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_234),
    .A2(n_21487),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_233),
    .Y(n_4762));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g14541 (.A(n_21534),
    .B(n_12531),
    .Y(n_4764));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g14542 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_249),
    .A2(n_4861),
    .B(n_4151),
    .Y(n_4767));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g14612 (.A1(n_4762),
    .A2(n_4764),
    .B(n_12532),
    .Y(n_4861));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g14614 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_257),
    .A2(n_4865),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_258),
    .B2(n_4864),
    .Y(n_4866));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1688 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_708));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1690 (.A1(n_4864),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_288));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1695 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_265),
    .B(n_4767),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_716));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_264),
    .B(n_4769),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_718));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1705_dup (.A1(n_4762),
    .A2(n_4764),
    .B(n_12532),
    .Y(n_4768));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_263),
    .B(n_4762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_720));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1712 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_268));
 AOI21xp5_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1715 (.A1(n_19472),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_265));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1716 (.A(n_4151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_264));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1717 (.A1(n_12531),
    .A2(n_21534),
    .B(n_12532),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_263));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_242),
    .B(n_21487),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_722));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1723 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1726 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_257));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1728 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_230),
    .B(n_19472),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_254));
 NOR2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1729 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_230),
    .B(n_19472),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_255));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1732 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1738 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_227),
    .B(n_19890),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_245));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_246));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_244));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_243));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_242));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1750 (.A(n_4487),
    .B(n_12402),
    .C(n_21951),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_238));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_237));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1752 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_235));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_236));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1754 (.A(n_6480),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_231));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1755 (.A(n_21530),
    .B(n_6483),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_234));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1756 (.A(n_6483),
    .B(n_21530),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_233));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_232));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1759 (.A(n_26011),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_191),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_230));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1760 (.A(n_26100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_25),
    .C(n_4224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_229));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1761 (.A(n_12424),
    .B(n_13546),
    .C(n_13552),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_228));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1762 (.A(n_12530),
    .B(n_12526),
    .C(n_5817),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_227));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1764 (.A(n_6479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_222));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_219));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_130),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_218));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_728));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1789 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_25));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1794 (.B(n_12397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_202),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_163));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_196));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1803 (.A(n_16140),
    .B(n_15921),
    .C(n_15920),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_195));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1806 (.A(n_13878),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_191));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_165),
    .B(n_14050),
    .C(n_14048),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_190));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1809 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_105),
    .B(n_19088),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_730));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_182));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_189));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_173));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_172));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_168));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1832 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_170));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1834 (.A(n_12398),
    .B(n_12400),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_163));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_72),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_167));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1837 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1838 (.A(n_12267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_5),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_165));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_159));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1853 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_153));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_149));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_147));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1869 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_141));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1874_dup26443 (.A(n_13873),
    .B(n_13874),
    .C(n_15795),
    .Y(n_13880));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_137));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_54),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_135));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_16),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_130));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1892 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_127));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1893 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_732));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_124));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1899 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_44),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_75),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_120));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1901 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_129));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1904 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_63),
    .B(n_12398),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_126));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_113));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_118));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_110));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1915 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_90),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_91),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_117));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1916 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_57),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_108));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_106));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_105));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_104));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_91));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .B(n_5737),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1945 (.A(n_16757),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_99));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1947 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1953 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1954 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1955 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(n_16749),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1957 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_23016),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_87));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_85));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_69));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1974 (.A(n_4386),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_68));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_58));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_48),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_49));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_44));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_66));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1987 (.A(n_2544),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_64));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_63));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_59));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_55));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_54));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2002 (.A(n_5737),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_45));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2007 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_40));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_35));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_34));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_33));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[23]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_32));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2023 (.A(n_12411),
    .B(n_12412),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_10));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2027 (.A(n_13874),
    .B(n_13873),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_6));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2028 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_5),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_0));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2031 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_2));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g2033 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_0));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g20810 (.A(n_12266),
    .Y(n_12267));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g20811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_59),
    .Y(n_12266));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g22117 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[20]),
    .Y(n_13873));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g22118 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(n_13874));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g22120 (.A1(n_13880),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_133),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_n_134),
    .B2(n_13877),
    .Y(n_13878));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_126_55_g23752 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[19]),
    .B(n_16757),
    .Y(n_15795));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_672));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_226),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_674));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_680));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1709 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_315));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1710 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_308),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_314));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1711 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_297),
    .A2(n_11043),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_313));
 OAI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1712 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_287),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_308),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_678));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_300),
    .B(n_11043),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_682));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1714 (.A(n_11045),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_684));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1715 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_277),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302),
    .B(n_4061),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_309));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1716 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_308),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_307));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1717 (.A1(n_11039),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_308));
 AOI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1720 (.A1(n_11041),
    .A2(n_20099),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278),
    .B1(n_20098),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_305));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_303));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1724 (.A1(n_17832),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_275),
    .B(n_17832),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_688));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1726 (.A(n_7883),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_300));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1728 (.A(n_20099),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_297));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1731 (.A(n_7883),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_295));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1735 (.A(n_4062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_293));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1736 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_292));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_291));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_268),
    .B(n_3819),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_690));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_287));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_286));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1744 (.A(n_10685),
    .B(n_11918),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_282));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1745 (.A(n_20088),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_285));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1747 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_280));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1748 (.A(n_2686),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_692));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_275));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_265),
    .B(n_7884),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_279));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1752 (.A(n_7884),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_278));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1753 (.A(n_20088),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_277));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_274));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_271));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_242),
    .B(n_22451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_273));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_259),
    .B(n_17829),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_268));
 NOR2x1_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_14),
    .B(n_20030),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1760 (.A(n_20030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_270));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1762 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_242),
    .B(n_22451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_267));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_223),
    .B(n_20034),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_265));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_12),
    .B(n_19901),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_264));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_261));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1769 (.A(n_17831),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1770 (.A(n_21411),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_694));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_260));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1779 (.A(n_21678),
    .B(n_19489),
    .C(n_19488),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_253));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_208),
    .B(n_9591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1784 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_208),
    .B(n_9591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_247));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1786 (.A1(n_21410),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_13),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_31));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1787 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_10),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_164),
    .C(n_11846),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1793 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_228),
    .B(n_8188),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_242));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_241));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1797 (.A(n_20095),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_238));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_228));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_224));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_225));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1827 (.A(n_23497),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_123),
    .B(n_19089),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_698));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_164),
    .B(n_11846),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_211));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_209));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1848 (.A1(n_24976),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_186),
    .B1(n_24977),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_202));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_153),
    .B(n_10856),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_201));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1850 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_208));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_148),
    .B(n_9389),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_195));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1858 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_132),
    .A2(n_20730),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_133),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_194));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_192));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_186));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1875 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_121),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_134),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_120),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_181));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_56),
    .B(n_19493),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_185));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1884 (.A(n_10856),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_176));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_179));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1891 (.B(n_21270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_178),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_91));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_174));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_171));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1909 (.A(n_19494),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_56),
    .C(n_19492),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1917 (.A(n_10982),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_156));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1918 (.A(n_20730),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_47),
    .B(n_11845),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1920 (.A(n_12806),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_99),
    .C(n_12802),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_22));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_157));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_153));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_149));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_700));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1930 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_68),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_41),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_69),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_146));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1934 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_44),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_43),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_142));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_148));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_135));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_133));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_131));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_130));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_128));
 AOI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_46),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_132));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1971 (.A(n_19892),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(n_14975),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(n_2958),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(n_14981),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_14179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_98));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_293),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_686));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(n_14186),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_85));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_81));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2014 (.A(n_2381),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_46));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_43),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_44));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_68));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(n_14987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[26]),
    .B(n_2944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[27]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_43));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2059 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[24]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[25]),
    .B(n_14179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_37));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_14));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2075 (.A(n_3946),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2077 (.A(n_8188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_10));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_9));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2080 (.A(n_10983),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_4));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_g2084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_128_55_n_3));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g14701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_75),
    .Y(n_4951));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_297),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_654));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g29214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_89),
    .Y(n_21805));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_223),
    .B(n_8178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_642));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_296),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_648));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2964 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_29),
    .A2(n_13364),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_315));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_307),
    .B(n_3642),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_650));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_298),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_652));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2970 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_302),
    .A2(n_12272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_306),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_29));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2971 (.A1(n_11064),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_312));
 OAI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2973 (.A1(n_13362),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_305),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_299),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_311));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_280),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_656));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_301),
    .B(n_13364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_307));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_306));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2979 (.A1(n_11065),
    .A2(n_21042),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_287),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_305));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2981 (.A(n_12272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_304));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2983 (.A(n_11064),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_302));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_301));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_299),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_300));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2988 (.A(n_7670),
    .B(n_20974),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_299));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2989 (.A(n_21042),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_298));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_290),
    .B(n_11064),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_297));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2991 (.A1(n_19487),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_296));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2993 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_260),
    .A2(n_5593),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_294));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2994 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_271),
    .B(n_5593),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_658));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_291));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2996 (.A(n_11065),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_290));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g2997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_287),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3002 (.A(n_26235),
    .B(n_21038),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_287));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_660));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_278),
    .B(n_7007),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_270),
    .B(n_19487),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_279));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_270),
    .B(n_19487),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_283));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3009 (.A(n_7008),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_278));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_272));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_271));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3018 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_248),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_27));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3019 (.A(n_20975),
    .B(n_26227),
    .C(n_20968),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_270));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_263));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3027 (.A(n_26183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_262));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3028 (.A(n_26183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_261));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3029 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_234),
    .B(n_22050),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_260));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_259));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3031 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_234),
    .B(n_22050),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_252),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_257));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_662));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3037 (.A(n_19485),
    .B(n_6606),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_253));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_252));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_210),
    .B(n_23398),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_210),
    .B(n_23398),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_250));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3041 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_249));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3042 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_226),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_248));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_247));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_242));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3050 (.A(n_6999),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_7),
    .C(n_22046),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_240));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_664));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_235));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3055 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_238));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3058 (.A(n_3746),
    .B(n_23394),
    .C(n_14951),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_234));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_228));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_226));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_229));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_227));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_223));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3069 (.A1(n_4434),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_225));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_224));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_150),
    .B(n_20884),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_26));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3076 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_5),
    .C(n_21804),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_25));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_220));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_666));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_215));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_212));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3092 (.A(n_9105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_208));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_119),
    .C(n_3955),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3099 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_183),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_202));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3101 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_5),
    .B(n_21804),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_201));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3103 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_205));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3105 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_199));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_46),
    .A2(n_10153),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_45),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_193));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3113 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_129),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_148),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_128),
    .B2(n_10646),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_188));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3115 (.A(n_7000),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_116),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_191));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3120 (.A(n_21866),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_182));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_178));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3122 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_177));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_176));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_49),
    .B(n_19136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_183));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_73),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_175));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3135 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_76),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_166));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_172));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_171));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3144 (.A(n_3229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_167));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_163));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3146 (.A(n_10153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_162));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3148 (.A(n_4951),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_158));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3150 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_165));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_164));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_64),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_154));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3158 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3160 (.A(n_10646),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_148));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3163 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3166 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_150));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_115),
    .B(n_21805),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_21));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_142));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_668));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_136));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_141));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3187 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_129));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_133));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3196 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_100),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_131));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_105),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_53),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_54),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_130));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_128));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_121));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_120));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_118));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3208 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_115));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3209 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_114));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3210 (.A(n_4965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_113));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .A2(n_3168),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B2(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_110));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_107));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_105));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_19));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_108));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_103));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_99));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3242 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3245 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_87));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3253 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_79));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3260 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3263 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_17));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_73));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_670));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_64));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_54));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3273 (.A(n_21856),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_45));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_41));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_34));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3283 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B(n_3168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_70));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_65));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3289 (.A(n_15192),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3290 (.A(n_3181),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_59));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_55));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3296 (.A(n_21861),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_51));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_49));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3304 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3306 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[32]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_42));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3307 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[35]),
    .B(n_6861),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3308 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[38]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_38));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3310 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3311 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[33]),
    .B(n_18041),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_36));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[36]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3313 (.A(n_4826),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_7));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3326 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_18),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3327 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_4),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_5));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3331 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_g3332 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[37]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_130_55_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_299),
    .B(n_19283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_622));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g22007 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .Y(n_13766));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g22034 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .Y(n_13790));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g22036 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .B(n_16772),
    .Y(n_13792));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g22040 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(n_16763),
    .Y(n_13796));
 AOI21xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2957 (.A1(n_19583),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_217),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_608));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2960 (.A(n_10793),
    .B(n_9880),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_616));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_309),
    .B(n_4029),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_618));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2966 (.A(n_22861),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_620));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2971 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_284),
    .A2(n_19283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_314));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2975 (.A(n_26210),
    .B(n_19289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_624));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2976 (.A(n_13952),
    .B(n_13082),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_310));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_303),
    .B(n_15079),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_309));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2978 (.A(n_22862),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_308));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_284),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_304));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2986 (.A(n_9879),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_303));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_299));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2992 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_264),
    .A2(n_12640),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_297));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2994 (.A(n_19291),
    .B(n_19288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_626));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_293));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2996 (.A(n_19594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_292));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g29966 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .B(n_22616),
    .Y(n_22619));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g29969 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .Y(n_22622));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2997 (.A(n_19595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_290));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g29975 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(n_22616),
    .Y(n_22628));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g2998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_264),
    .B(n_12639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g29980 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(n_22616),
    .Y(n_22633));
 NAND2x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g29981 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B(n_22616),
    .Y(n_22634));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3003 (.A(n_19274),
    .B(n_10860),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_628));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_267),
    .B(n_10754),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_284));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3010 (.A(n_12640),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_276));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g30167 (.A(n_22860),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_290),
    .Y(n_22861));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_207),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_9),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_267));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_265));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3027 (.A(n_19090),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3028 (.A(n_19090),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_630));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3037 (.A(n_6474),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_188),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_226),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_255));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3042 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_228),
    .A2(n_21025),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_249));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_226),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_244));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_632));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_237));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_156),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_233));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3063 (.A(n_21025),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_230));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_228));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3066 (.A(n_26228),
    .B(n_21028),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_231));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3069 (.A1(n_4435),
    .A2(n_6618),
    .B(n_6620),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_227));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_226));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_44),
    .C(n_13190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_220));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118),
    .B(n_19091),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_634));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3086 (.A(n_6620),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_214));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3087 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_213));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3088 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_168),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_185),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_167),
    .B2(n_9316),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_212));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3096 (.A(n_21015),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_117),
    .C(n_21013),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3101 (.A(n_20812),
    .B(n_20813),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_199));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3105 (.A(n_6618),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_159),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_43),
    .B2(n_13191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_191));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3116 (.A(n_22190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_188));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3118 (.A(n_9316),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_185));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_176));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_183));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_168));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3135 (.A(n_9180),
    .B(n_9179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_164));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_61),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_169));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3142 (.A(n_10423),
    .B(n_19304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_167));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3148 (.A(n_8019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_156));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_162));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_92),
    .B(n_13796),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_62),
    .C(n_13792),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_153));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3160 (.A(n_6710),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3163 (.A(n_22628),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3167 (.A(n_13790),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_106),
    .C(n_22633),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_147));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3172 (.A(n_9033),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_140));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_636));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3176 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_137),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_41));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3179 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_92),
    .B1(n_13796),
    .B2(n_22619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_134));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3187 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3188 (.A(n_13790),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_131));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_103),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_51),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_52),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_128));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_126));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_60),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_119));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_118));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_114));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3208 (.A(n_6949),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_113));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_110));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_67),
    .B(n_13936),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_109));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .A2(n_18049),
    .B1(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B2(n_23278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_108));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3216 (.A(n_13796),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_98));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3223 (.A(n_22619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_97));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3242 (.A(n_3309),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_96));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(n_3706),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_85));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3252 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_83));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_71));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_638));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3266 (.A(n_13766),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_64));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_62));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_59));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_43));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3283 (.A(n_19396),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[40]),
    .B(n_18049),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_68));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_67));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3289 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_61));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[41]),
    .B(n_23272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(n_19393),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[42]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[43]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3308 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[45]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[46]),
    .B(n_19395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_36));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3310 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[44]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_33));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3321 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_207),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_9),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_11));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3323 (.A(n_7874),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_9));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_114),
    .B(n_9033),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_g3331 (.A(n_13792),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_132_55_n_1));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_576));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_226),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_578));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1709 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_315));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1710 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_272),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_308),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_314));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1712 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_287),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_308),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_582));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_300),
    .B(n_12514),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_586));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1714 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_294),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_588));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1715 (.A1(n_19696),
    .A2(n_21577),
    .B(n_4286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_309));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1716 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_308),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_307));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1717 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_304),
    .A2(n_21577),
    .B(n_19503),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_308));
 NAND3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1721 (.A(n_12494),
    .B(n_19496),
    .C(n_19502),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_304));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_275),
    .B(n_21576),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_592));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1726 (.A(n_19504),
    .B(n_12512),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_300));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1734 (.A1(n_11762),
    .A2(n_8501),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_294));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1735 (.A(n_4287),
    .B(n_19696),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_293));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_291));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1738 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_32),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_290));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_268),
    .B(n_3860),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_594));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_287));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_286));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1744 (.A(n_8501),
    .B(n_11762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_282));
 NOR2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1746 (.A(n_8501),
    .B(n_11762),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_283));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1748 (.A(n_2781),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_596));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_275));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_274));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_271));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_242),
    .B(n_21284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_273));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_268));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_14),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_270));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1762 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_242),
    .B(n_21284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_267));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1763 (.A(n_22494),
    .B(n_21967),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_266));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_265));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1767 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_247),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_261));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1770 (.A(n_20965),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_598));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_243),
    .B(n_26184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_260));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1773 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1775 (.A(n_26184),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_190),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_254));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1784 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_247));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1786 (.A1(n_20965),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_13),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_31));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1787 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_10),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1793 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_228),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_5),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_242));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_241));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1795 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_240));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1803 (.A(n_20957),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_600));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1804 (.A(n_8951),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_233));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_216),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_154),
    .C(n_2873),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_231));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_3),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_228));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_30));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_224));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_225));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_29));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_602));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_199),
    .B(n_20966),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_211));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1840 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_210));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_215));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_209));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1850 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_208));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1854 (.A(n_20954),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_199));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_195));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1858 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_151),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_133),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_194));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_145),
    .B(n_10882),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_197));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1864 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_161),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_165),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_162),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1868 (.A(n_10882),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_190));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_186));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1873 (.A(n_25979),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_183));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1874 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_149),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_117),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_182));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1875 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_121),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_134),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_120),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_181));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_184));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_138),
    .B(n_2398),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_180));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1891 (.B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_178),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_91));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_177));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_172));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_166));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_161),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_163));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1903 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_161),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_162));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1904 (.A(n_17244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_170));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_74),
    .B(n_17250),
    .C(n_22869),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_165));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_164));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_161));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_160));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_156));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_93),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_99),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_22));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_103),
    .B(n_22882),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_18),
    .C(n_17249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_155));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_104),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_154));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1926 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_75),
    .B(n_17246),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_151));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_149));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1929 (.A1(n_17243),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_604));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1930 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_68),
    .A2(n_22877),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_69),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_146));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_144));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1933 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_78),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_79),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_143));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1934 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_44),
    .B1(n_22867),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_142));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1935 (.A(n_17249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_150));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1937 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_109),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_48),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_110),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_141));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_148));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_135));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_133));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1945 (.A(n_2398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_131));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1947 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_104),
    .B(n_17248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_129));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1948 (.A(n_22869),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_128));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_89),
    .B(n_17245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_127));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_46),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_132));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_124));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_72),
    .B(n_17243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_123));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_119));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_118));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_93));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1978 (.A(n_17248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_88));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_84));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_79));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_2930),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(n_3592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(n_3190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(n_2377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_2711),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2009 (.A(n_3479),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_78));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2014 (.A(n_2697),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_48),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_49));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_46));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2030 (.A(n_22867),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_44));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2032 (.A(n_22877),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2054 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(n_3479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_48));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(n_3479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_45));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[48]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_40));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_35));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_14));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_5),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_10));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_9));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_124),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_4));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2084 (.A(n_22882),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2085 (.A(n_17246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_2));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g2087 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[51]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25124 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(n_20459),
    .Y(n_17243));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25127 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(n_3408),
    .Y(n_17244));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25128 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(n_17245));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25129 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(n_2927),
    .Y(n_17246));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25130 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(n_22886),
    .Y(n_2398));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25131 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(n_3468),
    .Y(n_17248));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25132 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(n_17249));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g25133 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(n_17250));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g30174 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22867));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g30179 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22869));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g30187 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22877));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_134_55_g30192 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22882));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1743 (.A(n_6205),
    .B(n_6203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_552));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1746 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_298),
    .A2(n_21656),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_301),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_330));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1748 (.A(n_6201),
    .B(n_6199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_554));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1749 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_305),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_556));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1750 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_285),
    .A2(n_9746),
    .B(n_13172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_326));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_319),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_558));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1757 (.A(n_9746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_319));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_303),
    .B(n_20078),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_560));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1763 (.A(n_5617),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_313));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1769 (.A(n_10162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_307));
 NOR2xp33_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1771 (.A(n_5616),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_305));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1772 (.A(n_13173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_304));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1773 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_296),
    .B(n_9744),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_303));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1775 (.A1(n_21224),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_301));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1777 (.A(n_20082),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_562));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1778 (.A(n_9745),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_296));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_291));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1783 (.A(n_21222),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_298));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1788 (.A(n_22489),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_290));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1791 (.A(n_22488),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_285));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1798 (.A(n_21222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_282));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1801 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_280));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1803 (.A(n_8304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_278));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_233),
    .B(n_9430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_275));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1810 (.A(n_22221),
    .B(n_22480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_271));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_268));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1817 (.A(n_12576),
    .B(n_10888),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_266));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_263));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1823 (.A(n_11072),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_190),
    .C(n_3953),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_259));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1824 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_233),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_258));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_253));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1829 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_207),
    .B(n_6917),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_254));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_207),
    .B(n_6917),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_252));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1833 (.A(n_21293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_249));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_223),
    .B(n_20116),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_250));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1840 (.A(n_11763),
    .B(n_5575),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_243));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1841 (.A(n_5575),
    .B(n_11763),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_242));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1843 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_205),
    .B(n_21311),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_240));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1844 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_205),
    .B(n_21311),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_239));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1852 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_233));
 AOI21x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1864 (.A(n_11936),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_36));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1874 (.A(n_11936),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_223));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_214));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1886 (.A(n_20116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_208));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1888 (.A(n_10623),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_129),
    .B(n_19093),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_570));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_131),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_201));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_199));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1902 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_166),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_85),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_193));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1908 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_149),
    .B(n_21243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1910 (.A(n_21243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_190));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_182));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_188));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_184));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1934 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_179));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1939 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_0),
    .B(n_8320),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_172));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1942 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_166));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_165));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1949 (.A(n_13250),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1950 (.A(n_21218),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_108),
    .C(n_21220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_164));
 AOI21x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1952 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_33));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1969 (.A(n_4031),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_111),
    .C(n_13723),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_28));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1971 (.A(n_21157),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_107),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_153));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_572));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_146));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1980 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_93),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_91),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_25),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_145));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_143));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1997 (.A1(n_13236),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_138));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2002 (.A(n_13245),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_128));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2010 (.A(n_13241),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_126));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_23),
    .B(n_13247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_27));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_119),
    .B(n_12134),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2015 (.A(n_13236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_116));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_97));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2026 (.A(n_13710),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_95));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_25));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_2657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_110));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_108));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_11770),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(n_11770),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_98));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_92));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_43),
    .B(n_4549),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_90));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2064 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_67));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_40),
    .B(n_2747),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_n_574));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2094 (.A(n_2820),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2099 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(n_2820),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2107 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_21));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_66));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2111 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(n_2820),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(n_3375),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2116 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_47),
    .B(n_4555),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_57));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2121 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_53));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2126 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2137 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_17));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_188),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_107),
    .B(n_21157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2150 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_81),
    .B(n_14652),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_65),
    .B(n_13720),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_1));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21537 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .B(n_13231),
    .Y(n_13236));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_n_0));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21542 (.A(n_13231),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[62]),
    .Y(n_13241));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21546 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(n_13231),
    .Y(n_13245));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21548 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[63]),
    .B(n_13231),
    .Y(n_13247));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21551 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .B(n_2657),
    .Y(n_13250));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21954 (.A(n_13707),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[58]),
    .Y(n_13710));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g21964 (.A(u_NV_NVDLA_cmac_u_core_wt1_actv_data[60]),
    .B(n_13707),
    .Y(n_13720));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_mul_136_55_g23213 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt1_actv_data[57]),
    .Y(n_15157));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1_reg (.CLK(nvdla_core_clk),
    .D(n_5332),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d1));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2_reg (.CLK(nvdla_core_clk),
    .D(n_15),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d2));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_1_pp_pvld_d0_d3_reg (.CLK(nvdla_core_clk),
    .D(n_10),
    .QN(u_NV_NVDLA_cmac_u_core_out_mask[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1188),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1178),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_16477),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1176),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[12]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_16541),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[13]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_17940),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[14]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_5432),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[15]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_16259),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[16]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_5874),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[17]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_11165),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1187),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1186),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1185),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1184),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1183),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1182),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1181),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[7]));
 DFFHQNx1_ASAP7_75t_L \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1180),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[8]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_16529),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1169),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1159),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1158),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1157),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1156),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1154),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1153),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1152),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1151),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1150),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1168),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1167),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1166),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1165),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1164),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1163),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1162),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1161),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1160),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d2[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1148),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1136),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1135),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1133),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1132),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1131),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1130),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1129),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1127),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1126),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1147),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1146),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1144),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1142),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1141),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1140),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1139),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1138),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_1_sum_out_d0_d3_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1137),
    .QN(u_NV_NVDLA_cmac_u_core_out_data1[9]));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_448),
    .B(n_20637),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_180));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g24957 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(n_17072));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g24959 (.A(n_16782),
    .B(n_16785),
    .Y(n_17074));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g24960 (.A(n_17076),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_439),
    .Y(n_17077));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g24962 (.A1(n_17072),
    .A2(n_17073),
    .B(n_17074),
    .Y(n_17075));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g24963 (.A1(n_17075),
    .A2(n_6731),
    .B(n_23790),
    .Y(n_17078));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g25294 (.A(n_17416),
    .Y(n_17417));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g25295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_10),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_705),
    .Y(n_17416));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g25296 (.A(n_8886),
    .B(n_17419),
    .Y(n_17420));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g25297 (.A1(n_17417),
    .A2(n_21978),
    .B1(n_17418),
    .B2(n_17416),
    .Y(n_17419));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g25298 (.A(n_21978),
    .Y(n_17418));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g30069 (.A(n_22719),
    .B(n_22720),
    .Y(n_22721));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6011 (.A1(n_3649),
    .A2(n_5421),
    .B(n_3679),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_500));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_465),
    .B(n_24203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_186));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_451),
    .B(n_5421),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_184));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6021 (.A1(n_4842),
    .A2(n_20637),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_424),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_490));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_481),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_438),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_177));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6034 (.A(n_17072),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_481));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6036 (.A(n_3231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_450),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_176));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .C(n_14772),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_64));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6040 (.A(n_14773),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_175));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6046 (.A(n_14774),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_174));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6052 (.A(n_20629),
    .B(n_25447),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_465));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6057 (.A(n_20630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_455));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_453));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6062 (.A(n_3679),
    .B(n_3650),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_451));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_432),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_433),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_450));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6071 (.A(n_20629),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_445));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_173));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6075 (.A(n_6731),
    .B(n_23789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_439));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6076 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_412),
    .B(n_17074),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_438));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6077 (.A(n_4842),
    .B(n_10627),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_448));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_432));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_430));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6089 (.A(n_10627),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_424));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_433));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6095 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_372),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_431));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6096 (.A(n_20111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_399),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_429));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6101 (.A(n_11865),
    .B(n_9536),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_62));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6107 (.A(n_17073),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_412));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_380),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_172));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6125 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_397));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6126 (.A(n_14769),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_384),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_396));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6127 (.A(n_10696),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_401));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6129 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_346),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_399));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6130 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_356),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_398));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_347),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_395));
 MAJIxp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6139 (.A(n_17440),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_52),
    .C(n_3456),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_387));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6140 (.A(n_14771),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_384));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_345),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_171));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_385));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_381));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6145 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_380));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_308),
    .B(n_11334),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_379));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_305),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_375));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_343),
    .B(n_16059),
    .C(n_5433),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_373));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6157 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_331),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .C(n_10696),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_372));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_22),
    .B(n_12659),
    .C(n_4095),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_362));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6166 (.A(n_11246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_357));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_356));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6169 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_331),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_354));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_361));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_359));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_358));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6177 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .A2(n_6351),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_314),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_349));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6180 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_291),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_313),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_347));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_352));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6182 (.A1(n_15227),
    .A2(n_17420),
    .B1(n_15068),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_316),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_346));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6183 (.A1(n_19096),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_345));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_344));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6186 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_297),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_343));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6196 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_330));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_337));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_328));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6201 (.A(n_19096),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_327));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_326));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6203 (.A(n_19096),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_336));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6208 (.A(n_15553),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_58));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6210 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_276),
    .B(n_10694),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_332));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_273),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_331));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6213 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_325));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_322));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6219 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_314));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_308));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_324));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_321));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6227 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_214),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_320));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6228 (.A(n_21972),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_243),
    .C(n_23466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_319));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_318));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6231 (.A(n_10693),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_317));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6232 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_264),
    .B(n_23467),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_316));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6233 (.A(n_12887),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .C(n_2442),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_315));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6234 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_211),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_312));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6239 (.A(n_6351),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_305));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6242 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_300));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6243 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_307));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6251 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_298));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6255 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_291));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6257 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_52));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6260 (.A(n_6296),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_297));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_290));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6267 (.A(n_6296),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118),
    .C(n_8886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_288));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6272 (.A1(n_2582),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_281));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_280));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6274 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_217),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_279));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6278 (.A(n_2580),
    .B(n_14110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_278));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6279 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .A2(n_2442),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .B2(n_2441),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_277));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_276));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_275));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_283));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6289 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_267));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6290 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_265));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6292 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6293 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_254));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6294 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_273));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6297 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_138),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_270));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6300 (.A(n_2275),
    .B(n_5494),
    .C(n_14683),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_266));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_140),
    .C(n_21056),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_264));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_263));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6304 (.A(n_19097),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .C(n_19098),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_261));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6305 (.A(n_26186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_260));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6306 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_259));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6307 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_216),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_258));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6308 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_120),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_256));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6309 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6315 (.A(n_17552),
    .B(n_5393),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_247));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_251));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6324 (.A(n_13097),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_243));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6327 (.A(n_12884),
    .B(n_12882),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_240));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6328 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_137),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_164),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_138),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_239));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_237));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6333 (.A1(n_8886),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_234));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6337 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_233));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6338 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_231));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6350 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37),
    .A2(n_14109),
    .B(n_14108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6351 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_232));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6352 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_230));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6353 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_697),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_228));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6357 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_224));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6358 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_223));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6360 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_222),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6362 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_221));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_216));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6374 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6376 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_204));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6377 (.A1(n_2580),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118),
    .B1(n_2582),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_203));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6379 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6380 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_215));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6381 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_659),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_627),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_214));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6382 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_129),
    .B(n_22720),
    .C(n_22719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_213));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6385 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_631),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6386 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_653),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_621),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_210));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6388 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_643),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_739),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_42));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6389 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_209));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_657),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_207));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6405 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_200));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6412 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_663),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_699),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_190));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_633),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_185));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6423 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_169),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_170));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6424 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6428 (.A(n_17416),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6430 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_797),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6435 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_713),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_175));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6436 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6437 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_757),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_173));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6439 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_745),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6440 (.A(n_5492),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_169));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6441 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_168));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6442 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_167));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6444 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_729),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_165));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6445 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_723),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_163),
    .A(n_12996));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6449 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_154));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6452 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_148));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_601),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_88),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_161));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6458 (.A(n_23445),
    .B(n_23014),
    .C(n_21052),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6459 (.A(n_19061),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_767),
    .C(n_19060),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6462 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_565),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_789),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_725),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6465 (.A(n_12997),
    .B(n_14812),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_723),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6466 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_733),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_637),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_797),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_713),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_553),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_639),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_671),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_143));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6471 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_745),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_585),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_141));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6472 (.A(n_8850),
    .B(n_8853),
    .C(n_13676),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6473 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_138));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6475 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_133));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_131));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6477 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_129));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6486 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_118));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6492 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_757),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_693),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_597),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_137));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6494 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_701),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6495 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_559),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_783),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_793),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_729),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_130));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6497 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_599),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_727),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_567),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_128));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6500 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_695),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_663),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_125));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_761),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_665),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_633),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_123));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_763),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_635),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_667),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_122));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_603),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_731),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_n_699),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_121));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6505 (.A(n_8670),
    .B(n_5399),
    .C(n_5400),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_120));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6508 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_705),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_70),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_37));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_597),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_693),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_111));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6514 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_761),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_109));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_791),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_695),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_108));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_667),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_763),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_107));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_106));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6530 (.A(n_19063),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_575),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_115));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_625),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_100));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_565),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_98));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6545 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_731),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_96));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6546 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_659),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_627),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_95));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6551 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_567),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_599),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_92));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_637),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_733),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_91));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6553 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_90));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_691),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_89));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6556 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_571),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_102));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_795),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6559 (.A(n_23424),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_575),
    .B(n_19063),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_82));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6578 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_613),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_76));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6579 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_75));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6588 (.A(n_10262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_71));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6622 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .A(n_15361));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6623 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_32));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6627 (.A(n_23467),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_28));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6629 (.A(n_8956),
    .B(n_8954),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_26));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6630 (.A(n_26186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_25));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6632 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_23));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6633 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_22));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6634 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_21));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6636 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_777),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_19));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6637 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_621),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_653),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_18));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6638 (.A(n_9650),
    .B(n_9652),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_17));
 XOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6640 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_643),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_15),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_739));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6641 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_581),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_677),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_14));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6642 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_13),
    .A(n_23424));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6643 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_591),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_12));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6645 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_10),
    .A(n_10262));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6648 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_559),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_783),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6650 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_n_585),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_5));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_g6651 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_n_673),
    .B(n_12550),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_csa_tree_ADD_TC_OP_6_groupi_n_4));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_285),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_746));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2959 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_268),
    .A2(n_11857),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_270),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_197),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_736));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_738));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_299),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_740));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_271),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_298),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_744));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2963 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_293),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_299));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2964 (.A1(n_4074),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_298));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2965 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_268),
    .A2(n_11857),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_297));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2966 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_264),
    .A2(n_11857),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_265),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_742));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_748));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2969 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_263),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_287),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_294));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2970 (.A(n_11857),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_293));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_281),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_292));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2975 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_274),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_288),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_273),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_287),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_750));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_289));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2978 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_287));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2979 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_256),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_22),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_288));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_752));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_277),
    .B(n_4075),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_285));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_284));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_283));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2985 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_281));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2986 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_258),
    .A2(n_14836),
    .B(n_14835),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2989 (.A(n_14837),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_23));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_278));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_277));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2992 (.A(n_14837),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_276));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2993 (.A(n_14836),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_275));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2994 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_274));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_273));
 AOI21xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2996 (.A1(n_12606),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2997 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_271));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g2998 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_239),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_270));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3000 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_241),
    .A2(n_10481),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_22));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_250),
    .B(n_6960),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_754));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_265));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3003 (.A(n_14835),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_262));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_268));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_231),
    .B(n_12606),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_266));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_264));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_263));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3012 (.A(n_14838),
    .B(n_19195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_260));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_231),
    .B(n_12606),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_256));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3015 (.A(n_13586),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_259));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_258));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3018 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_252));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_240),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_250));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_254));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_253));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3029 (.A(n_11175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_249));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3030 (.B(n_20336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_248),
    .A(n_8442));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_240));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3037 (.A(n_26187),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_239));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3038 (.A(n_26187),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_238));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_237));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_236));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3044 (.A(n_11175),
    .B(n_11177),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_232));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3045 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_170),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_231));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3046 (.A(n_12597),
    .B(n_12603),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_216),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_229));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_224));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3054 (.A(n_11177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_223));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_219));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_760));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_189),
    .B(n_19712),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_216));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3066 (.A(n_8442),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_212));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_132),
    .C(n_4331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_208));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3072 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_197),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_204));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_178),
    .B(n_12929),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_206));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3075 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_177),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_205));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3078 (.A(n_6242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_200));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3080 (.A(n_19185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_199));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3082 (.A(n_8233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_142),
    .C(n_5398),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_203));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_35),
    .C(n_6305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_202));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3087 (.A(n_19712),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_196));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3088 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106),
    .B(n_19099),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_762));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_180),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_192));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3091 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3092 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_190));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_189));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_197));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_188));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_182));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3105 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_179));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3106 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_181));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_35),
    .B(n_6305),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_177));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_175));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3123 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3125 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_162));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_117),
    .B(n_9060),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_170));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_158));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_74),
    .C(n_25982),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_159));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_44),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_157));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_155));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_153));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_63),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_48),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_145));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3154 (.A(n_9060),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_33),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_81),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_140));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3168 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3169 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_10),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_13));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_764));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_126));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3177 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_76),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_10),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3180 (.A(n_18751),
    .B(n_9059),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_131));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3183 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_117));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_116));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_115));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_121));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_81),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_110));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3192 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_120));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3193 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_118));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_109));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3197 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_107));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3198 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_106));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_103));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_102));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3203 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_101));
 AOI22xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3206 (.A1(n_4463),
    .A2(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B1(n_3761),
    .B2(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_98));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_766));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_77));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_10));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_73));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3221 (.A(n_3150),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3222 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3227 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(n_3760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3228 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_87));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3231 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(n_3275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3232 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_85));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_82));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_80));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3237 (.A(n_3148),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3239 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_11));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3242 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_68));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3247 (.A(n_2325),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(n_6972),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_63));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3255 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_51));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_42));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3260 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_37));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_33));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_62));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3266 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_57));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3269 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3270 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3271 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3274 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_47));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3275 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[7]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3279 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_36));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3283 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_35));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_32));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[3]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_31));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[0]),
    .B(n_6973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_29));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3289 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[5]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_28));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_27));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[1]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_25));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3295 (.A(n_13586),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3297 (.A(n_8233),
    .B(n_5398),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_2));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[4]),
    .B(n_2337),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_122_55_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1743 (.A(n_19132),
    .B(n_10816),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_776));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1748 (.A(n_10814),
    .B(n_14802),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_778));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1767 (.A(n_19732),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_309));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1771 (.A(n_5487),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_305));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_285),
    .B(n_7342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_304));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1775 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_281),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_301));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1778 (.A(n_8826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_296));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_294));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1780 (.A(n_7342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_292));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_291));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_283),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_298));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1786 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_281),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_293));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1788 (.A(n_7343),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_290));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1791 (.A(n_11858),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_285));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1798 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_282));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_17),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_283));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_281));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1801 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_265),
    .B(n_8821),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_279));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_233),
    .B(n_10129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_275));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1808 (.A(n_10071),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_273));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_271));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1811 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_269),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_270));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1812 (.A(n_2735),
    .B(n_12661),
    .C(n_12665),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_269));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1814 (.A(n_8823),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1815 (.A(n_21452),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_267));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_193),
    .B(n_21452),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1820 (.A(n_2634),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_790));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1823 (.A(n_10071),
    .B(n_19967),
    .C(n_3030),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_259));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1824 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_233),
    .A2(n_10131),
    .B(n_10130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_258));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1834 (.A(n_19967),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_247));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1836 (.A1(n_22735),
    .A2(n_3553),
    .B1(n_22734),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_245));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1842 (.A(n_22980),
    .B(n_26059),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_792));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_229),
    .B(n_8661),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_14),
    .B(n_20306),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_234));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1852 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_33),
    .B(n_20200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_233));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1854 (.A(n_8665),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1864 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_36));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1874 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_186),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_223));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_171),
    .C(n_10777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_222));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_151),
    .B(n_20304),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_218));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_211));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_213));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1888 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_204),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1889 (.A(n_22978),
    .B(n_26207),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_794));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_131),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_207));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_11),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_204));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1900 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_27),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_31),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_197));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1902 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_86),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_166),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_85),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_193));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_5),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_127),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_191));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_182));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1920 (.A(n_9912),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_187));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_186));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_170));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1934 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1937 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_50),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_174));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1939 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_172));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1940 (.A(n_15289),
    .B(n_15588),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_171));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1942 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_166));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_165));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1950 (.A(n_25335),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_108),
    .C(n_20514),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_164));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1952 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_33));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1953 (.A(n_22840),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_20),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_81),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1958 (.A(n_11943),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1959 (.A(n_11090),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_156));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1964 (.A(n_15290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_113),
    .C(n_15588),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_31));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_159));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_93),
    .C(n_15239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_29));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_118),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_154));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_152));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_122),
    .B(n_22978),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_796));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_149));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1977 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_56),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_103),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_104),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_148));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1978 (.A1(n_9905),
    .A2(n_22954),
    .B1(n_22953),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_147));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_143));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1984 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_23),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_27),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_151));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1997 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_115),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_138));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2 (.A(n_8667),
    .B(n_14814),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_788));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_134));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_128));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_127));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_126));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_23),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_27));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_103));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_123));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_113));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_112));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_110));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .B(n_6576),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_98));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_92));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_43),
    .B(n_3107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(n_14537),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2064 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_67));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_56));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_40),
    .B(n_4528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_798));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2094 (.A(n_6576),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2095 (.A(n_18692),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2096 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_48));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2098 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2099 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_73));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2105 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[15]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2116 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_47),
    .B(n_3113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_58));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2120 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2122 (.A(n_18692),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2124 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_50));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_43));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2137 (.A(n_21448),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_17));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_29),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_171),
    .B(n_10777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_127),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_11));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_112),
    .B(n_18947),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_107),
    .B(n_15590),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_5));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2150 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_81),
    .B(n_22840),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g2154 (.A(n_11942),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_0));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23199 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(n_9349),
    .Y(n_15142));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23201 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(n_15144));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23204 (.A(n_15144),
    .B(n_15142),
    .Y(n_15145));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23294 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_96),
    .Y(n_15290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23556 (.A(n_24402),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[13]),
    .Y(n_15588));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g23558 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[9]),
    .B(n_24402),
    .Y(n_15590));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g30080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_187),
    .Y(n_22735));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g30150 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[11]),
    .B(n_22834),
    .Y(n_22840));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_g30262 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_124_55_n_218),
    .Y(n_22952));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1688 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_708));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1689 (.A(n_6991),
    .B(n_6993),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_712));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1690 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_246),
    .A2(n_16564),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_288));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1694 (.A(n_6988),
    .B(n_24916),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_714));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1695 (.A(n_6366),
    .B(n_21256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_716));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1699 (.A(n_24916),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_279));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1701 (.A(n_21255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_718));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1704 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_273));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1705 (.A1(n_16327),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_274));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_263),
    .B(n_10247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_720));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1712 (.A(n_6354),
    .B(n_24912),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_268));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1717 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_13),
    .A2(n_20108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_263));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1719 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_244),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_261));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1722 (.A(n_10248),
    .B(n_8351),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_722));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1723 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_258));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_259));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1726 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_244),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_257));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1727 (.A(n_20108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_256));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1732 (.A(n_6354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_248));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1734 (.A(n_20108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_247));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_245));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_246));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_244));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_243));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1747 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_216),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_241));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1750 (.A(n_22738),
    .B(n_22737),
    .C(n_12218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_238));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_237));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1752 (.A(n_16324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_235));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_236));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_232));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_203),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_726));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_11),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_191),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_230));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1761 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_164),
    .C(n_8881),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_228));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1764 (.A(n_8347),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_222));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1766 (.A(n_26119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_204),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_224));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_164),
    .B(n_8881),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_216));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1773 (.A(n_12900),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_215));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_130),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_218));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_152),
    .B(n_5411),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_213));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_728));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1781 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1783 (.A(n_12899),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_208));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1787 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_131),
    .C(n_5385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1792 (.A(n_9467),
    .B(n_5512),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_204));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1793 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_170),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_203));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_196));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1799 (.A(n_12900),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_139),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_146),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_197));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1803 (.A(n_8878),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_195));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_162),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1809 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_105),
    .B(n_19101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_730));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_185));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1812 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_183));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_182));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_189));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_187));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1819 (.A(n_12893),
    .B(n_12894),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_177));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1823 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_139),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1824 (.A(n_19164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_134),
    .C(n_5378),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_178));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_173));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_172));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1831 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_171));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1832 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_170));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1835 (.A1(n_5378),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_133),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_138),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_162));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_72),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_167));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1837 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_78),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1844 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_154));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_159));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1852 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1853 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_152));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1857 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_69),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_150));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_147));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1862 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_145));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1866 (.A(n_5378),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_138));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1869 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1870 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_141));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1871 (.A(n_12214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_49),
    .C(n_20488),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_140));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1873 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_45),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_95),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_139));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_137));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_134));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_19));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1885 (.A(n_9842),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_55),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_20));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_16),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_98),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1888 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_94),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_131));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_33),
    .B(n_8872),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_130));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1891 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_128));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1892 (.A(n_19164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_127));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1893 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_732));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_124));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1895 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_39),
    .A2(n_14353),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_38),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_84),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_122));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_121));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_114));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_113));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_118));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_110));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1915 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_90),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_91),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_117));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1916 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_57),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_116));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1917 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_115),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_108));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_106));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_105));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_104));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_91));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1935 (.A(n_14353),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1936 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_81));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .B(n_5737),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1945 (.A(n_16757),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_99));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_98));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1947 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_95));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_94));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1951 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1953 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1954 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(n_16749),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1957 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_88));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_86));
 NAND2x1_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_78));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1974 (.A(n_4386),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_68));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_58));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1981 (.A(n_12215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_49));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_44));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_66));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1987 (.A(n_2544),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_64));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_63));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_59));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_55));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_54));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(n_16757),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_51));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2 (.A(n_5413),
    .B(n_8352),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_724));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_50));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2002 (.A(n_5737),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2004 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_45));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_42));
 NAND2x1p5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2009 (.A(n_16749),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[16]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_35));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_33));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[23]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_32));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_208),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_12),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_9),
    .B(n_5517),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2022 (.A(n_8512),
    .B(n_18974),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_11));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2024 (.A(n_21251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_93),
    .B(n_5375),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_6));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2028 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_5),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_0));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2031 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_2));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g2033 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20759 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(n_12213));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20760 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[21]),
    .B(n_16749),
    .Y(n_12214));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20761 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(n_12215));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20763 (.A(n_12214),
    .B(n_12216),
    .Y(n_12217));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20764 (.A(n_12213),
    .B(n_12215),
    .Y(n_12216));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g20765 (.A(n_11534),
    .B(n_12217),
    .Y(n_12219));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g23754 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[19]),
    .B(n_16753),
    .Y(n_15798));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g30082 (.A(n_10078),
    .Y(n_22737));
 INVx1_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_g30083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_126_55_n_209),
    .Y(n_22738));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_672));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_226),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_315),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_674));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1707 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_269),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_676));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_292),
    .B(n_10479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_680));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1709 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_315));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1710 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_272),
    .A2(n_13605),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_314));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1712 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_287),
    .B2(n_13605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_678));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1714 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_294),
    .B(n_13609),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_684));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1716 (.A(n_13605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_307));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1726 (.A(n_12681),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_300));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1728 (.A(n_19377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_297));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1731 (.A(n_12681),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_295));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1734 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252),
    .B(n_19382),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_294));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1735 (.A(n_4251),
    .B(n_19381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_293));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1736 (.A(n_19378),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_292));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_291));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_268),
    .B(n_3815),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_690));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_287));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_286));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1748 (.A(n_2689),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_692));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_274));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_271));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_269));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1757 (.A(n_25602),
    .B(n_25603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_273));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_268));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_14),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_270));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_12),
    .B(n_22731),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_264));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1766 (.B(n_9451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_263),
    .A(n_25504));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1767 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_247),
    .A2(n_17474),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_261));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_259));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_246),
    .B(n_7335),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_260));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1773 (.A(n_7335),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_258));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1777 (.A(n_13575),
    .B(n_21160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_250));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1778 (.A(n_18786),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_190),
    .C(n_19803),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_254));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1780 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_12),
    .B(n_3877),
    .C(n_26033),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_252));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1782 (.A(n_7572),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1784 (.A(n_7572),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_247));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1787 (.A(n_18884),
    .B(n_22989),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_243));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1794 (.A(n_6639),
    .B(n_18868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_241));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1795 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_215),
    .B(n_7332),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_240));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1796 (.A(n_21160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_239));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1799 (.A(n_22726),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_237));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1803 (.A(n_17470),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_696));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1807 (.A(n_6639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_230));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_226));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1826 (.A(n_19801),
    .B(n_12281),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_225));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1828 (.A(n_25499),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_29));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_123),
    .B(n_19102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_698));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_199),
    .B(n_17472),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_211));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_215));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1843 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_206));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1847 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_187),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_156),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_25),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_203));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1848 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_173),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_186),
    .B1(n_13577),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1852 (.A(n_22988),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_132),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_205));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1854 (.A(n_17471),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_199));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1858 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_132),
    .A2(n_7336),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_133),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_194));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1864 (.A1(n_14785),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_165),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_162),
    .B2(n_25500),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_190));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1871 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_187));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_186));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1878 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_25));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1884 (.A(n_21162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_176));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1886 (.A(n_13577),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_138),
    .B(n_2642),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_174));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1903 (.A(n_14785),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_162));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_74),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_165));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_156));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1918 (.A(n_7336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_93),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_99),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_155));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_149));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_700));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1930 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_68),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_41),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_69),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_146));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_144));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1933 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_78),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_79),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_143));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1934 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_44),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_43),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_142));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_140));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_135));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_133));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_131));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_130));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_128));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_126));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_46),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_103),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_132));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_119));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_118));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_116));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_114),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1971 (.A(n_14784),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_108));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_84));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(n_14981),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(n_2944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_111));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_14987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(n_21990),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_14179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_100));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(n_14987),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_95));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2003 (.A(n_12800),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_2392),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_89));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_80));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2013 (.A(n_21990),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_78));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2014 (.A(n_2381),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_46));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_43),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_44));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(n_14978),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(n_2944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_47));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[27]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_45));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_43));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2059 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[24]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_39));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .B(n_3504),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34),
    .B(n_14183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2065 (.A(n_14975),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_36));
 BUFx2_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2069 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_34));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_190),
    .B(n_19802),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2075 (.A(n_3971),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2076 (.A(n_22727),
    .B(n_22725),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_11));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_6));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g20825 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_76),
    .Y(n_12281));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_4));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25341 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_168),
    .Y(n_17470));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25342 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_122),
    .Y(n_17471));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25343 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_179),
    .Y(n_17472));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25344 (.A1(n_17473),
    .A2(n_18868),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_230),
    .Y(n_17474));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25345 (.A1(n_17471),
    .A2(n_17470),
    .B(n_17472),
    .Y(n_17473));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g25346 (.A(n_17473),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_241),
    .Y(n_17475));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g30071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_21),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_128),
    .Y(n_22725));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g30074 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_29),
    .A2(n_22728),
    .B1(n_3878),
    .B2(n_26033),
    .Y(n_22731));
 MAJIxp5_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g30075 (.A(n_22725),
    .B(n_22726),
    .C(n_22727),
    .Y(n_22728));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32579 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_115),
    .Y(n_25499));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32580 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_165),
    .Y(n_25500));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32582 (.A(n_14785),
    .B(n_25500),
    .C(n_25499),
    .Y(n_25502));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32584 (.A(n_25502),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_203),
    .Y(n_25504));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32659 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_237),
    .B(n_7459),
    .Y(n_25603));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32661 (.A(n_25603),
    .B(n_25602),
    .Y(n_25604));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_g32663 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_128_55_n_274),
    .B(n_25604),
    .Y(n_25607));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g21630 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_40),
    .Y(n_13328));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_272),
    .B(n_10185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_644));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2960 (.A(n_23072),
    .B(n_23070),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_648));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_285),
    .B(n_23058),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_646));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2965 (.A(n_23071),
    .B(n_3647),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_650));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_298),
    .B(n_10038),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_652));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2975 (.A(n_6230),
    .B(n_6235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_656));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2989 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_292),
    .B(n_25983),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_298));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_297));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2992 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_295));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_291));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2996 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_290));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_262),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_286));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g2999 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_285));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3000 (.A(n_19808),
    .B(n_6589),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_292));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_265),
    .B(n_19367),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_289));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_660));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_232),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_12),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_284));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_265),
    .B(n_19367),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_282));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_272));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_275));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_273));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3019 (.A(n_20401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_219),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_270));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3021 (.B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_268),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_233));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3023 (.A(n_19804),
    .B(n_3905),
    .C(n_8846),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_266));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3024 (.A(n_6592),
    .B(n_19360),
    .C(n_9322),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_265));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_263));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3027 (.A(n_19103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_262));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3028 (.A(n_19103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_261));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_252),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_662));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3036 (.A(n_9321),
    .B(n_6592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_254));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3037 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_233),
    .B(n_14826),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_253));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_252));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_210),
    .B(n_8840),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_210),
    .B(n_8840),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_250));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3041 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_249));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3042 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_226),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_248));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_247));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3046 (.A(n_14826),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_244));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_10),
    .B(n_7685),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_242));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3049 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_241));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3050 (.A(n_7685),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_7),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_240));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_664));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_235));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3056 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_189),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_211),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_237));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3059 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_189),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_151),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_233));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3060 (.A(n_18748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_184),
    .C(n_26200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_232));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_228));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_226));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_229));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_227));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_72),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_223));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3069 (.A1(n_4438),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_225));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_224));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_150),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_26));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_220));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3080 (.A(n_23035),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_113),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120),
    .B(n_19104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_666));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_215));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_154),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_212));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_151),
    .B(n_11941),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_119),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_209));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3105 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_199));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3109 (.A1(n_15071),
    .A2(n_15462),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_143),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_196));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_46),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_161),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_45),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_195));
 AOI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3111 (.A1(n_6284),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_111),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_22),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_194));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_193));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3113 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_129),
    .A2(n_19355),
    .B1(n_19353),
    .B2(n_19354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_152),
    .B(n_14825),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_189));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3120 (.A(n_11941),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_182));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_176));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_183));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_73),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_175));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_172));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_171));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3144 (.A(n_3233),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_77),
    .C(n_9269),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_167));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_161),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_162));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3149 (.A(n_7686),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_156));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_164));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3152 (.A(n_19615),
    .B(n_19612),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_161));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_64),
    .C(n_22745),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_154));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3158 (.A(n_6284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_22));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_49),
    .C(n_8738),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_86),
    .B(n_23033),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3166 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_150));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3169 (.A(n_9274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_57),
    .C(n_13328),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_145));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_142));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_668));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_136));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3182 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_66),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_48),
    .B1(n_8738),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_134));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3184 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_69),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_143));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_141));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3187 (.A(n_19353),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_129));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_133));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3196 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_100),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_131));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_105),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_53),
    .B1(n_13699),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_121));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_120));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_116));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3210 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_113));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_112));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_69),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_111));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .A2(n_3168),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B2(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_110));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_105));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3220 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_19));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_90));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_86));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_77));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_74));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_31),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_104));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_103));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_99));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3242 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3252 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3253 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3260 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3263 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_17));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_73));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_670));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3266 (.A(n_8738),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_66));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_64));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_48));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_45));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3282 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_34));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3283 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B(n_3168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_70));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_69));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3289 (.A(n_15192),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3290 (.A(n_3181),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_59));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3293 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[36]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3297 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_51));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_49));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3306 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[32]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_42));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3307 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[35]),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3308 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[37]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[38]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_38));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3310 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3311 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[33]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3313 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[34]),
    .B(n_4826),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_33));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3314 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[36]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_32));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3315 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[36]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_31));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3320 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_219),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_12));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_7),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_7));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3326 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_18),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_g3331 (.A(n_22744),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_130_55_n_1));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_299),
    .B(n_20345),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_622));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22015 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_16763),
    .Y(n_13771));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22020 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_16772),
    .Y(n_13776));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22021 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_16769),
    .Y(n_13777));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22031 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .B(n_16763),
    .Y(n_13787));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .B(n_16769),
    .Y(n_13791));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g22038 (.A(n_16772),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .Y(n_13794));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_225),
    .B(n_7906),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_610));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2964 (.A1(n_7618),
    .A2(n_20346),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_317));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2966 (.A(n_13091),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_620));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2971 (.A1(n_10561),
    .A2(n_20345),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_314));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2975 (.A(n_7060),
    .B(n_7064),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_624));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2976 (.A(n_23031),
    .B(n_7618),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_310));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2983 (.A(n_10561),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_304));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_303));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2987 (.A(n_7619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_302));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_292),
    .B(n_10561),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_299));
 AOI21xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2991 (.A1(n_15353),
    .A2(n_9126),
    .B(n_23031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_298));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_293));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2996 (.A(n_11790),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_292));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g29965 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_22616),
    .Y(n_22618));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g29967 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .Y(n_22620));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g2997 (.A(n_13089),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g29976 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .Y(n_22629));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g29978 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .B(n_22616),
    .Y(n_22631));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g29979 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_22616),
    .Y(n_22632));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_250),
    .B(n_22511),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_628));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3006 (.A(n_9126),
    .B(n_15353),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_281));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3012 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_274));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3022 (.A(n_23450),
    .B(n_14211),
    .C(n_11791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_269));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_265));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3027 (.A(n_19105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3028 (.A(n_19105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_630));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3037 (.A(n_10999),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_188),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_226),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_255));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3042 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_228),
    .A2(n_8861),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_249));
 XOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3046 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_188),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_246),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_10),
    .B(n_11327),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_244));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3049 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3050 (.A(n_11327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_7),
    .C(n_3611),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_242));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_632));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_237));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3063 (.A(n_8861),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_230));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_228));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3066 (.A(n_8855),
    .B(n_20222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_231));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_70),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_225));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3069 (.A1(n_4439),
    .A2(n_7352),
    .B(n_7354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_227));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_226));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_44),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_220));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118),
    .B(n_19106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_634));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3086 (.A(n_7354),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_214));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_211));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3095 (.A(n_22521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_203));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3105 (.A(n_7352),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_44),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_159),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_43),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_160),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_191));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3113 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_127),
    .A2(n_8866),
    .B1(n_8864),
    .B2(n_8865),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_186));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3116 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_86),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_188));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_187));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_176));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_61),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_169));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_160));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_156));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_162));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_92),
    .B(n_13791),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_157));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3154 (.A(n_7166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_155));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_62),
    .C(n_13787),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_153));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3158 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3161 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3163 (.A(n_22618),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_79),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_152));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_47),
    .C(n_13777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_84),
    .C(n_14675),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_150));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3166 (.A(n_21911),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3167 (.A(n_13794),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_106),
    .C(n_22632),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3169 (.A(n_15081),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_55),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_143));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3170 (.A(n_18771),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_88),
    .C(n_20480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_21));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3172 (.A(n_22741),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_140));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_636));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3176 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_86),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3179 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_92),
    .B1(n_13791),
    .B2(n_22629),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_134));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3181 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_88),
    .A2(n_20481),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_17),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_133));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3182 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_46),
    .B1(n_13777),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3187 (.A(n_8864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_131));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_60),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_119));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_118));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_114));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3211 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_110));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_67),
    .B(n_13771),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_109));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .A2(n_18049),
    .B1(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .B2(n_23278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_108));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3216 (.A(n_13791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3223 (.A(n_22629),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_92));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_88));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_101));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3242 (.A(n_3309),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_87));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_3706),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3252 (.A(n_3317),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3256 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_3713),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3263 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_17));
 NAND2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_71));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_638));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3266 (.A(n_13777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_64));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_62));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_43));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3283 (.A(n_19396),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .B(n_18049),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_68));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_67));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3289 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_61));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3293 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_2990),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_55));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[41]),
    .B(n_23272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_19393),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[42]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[45]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3304 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[40]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[43]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[46]),
    .B(n_19395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_36));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3310 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[44]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_7),
    .B(n_3611),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3324 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_114),
    .B(n_22741),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3325 (.A(n_7166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_g3331 (.A(n_13787),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_132_55_n_1));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_288),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_291),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_213),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_576));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1707 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_269),
    .B(n_23436),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_580));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1708 (.A(n_19243),
    .B(n_11483),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_584));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1712 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_286),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_287),
    .B2(n_23434),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_582));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1714 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_294),
    .B(n_11489),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_588));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1716 (.A(n_23434),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_307));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1728 (.A(n_9206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_297));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1731 (.A(n_9209),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_295));
 AOI21xp5_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1734 (.A1(n_15380),
    .A2(n_14105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_294));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1737 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_270),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_257),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_291));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_268),
    .B(n_3880),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_594));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_287));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_270),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_286));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1744 (.A(n_14105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_282));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1745 (.A(n_8214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_285));
 NOR2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1746 (.A(n_14105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_283));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1748 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_255),
    .B(n_2785),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_596));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1755 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_272),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_271));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_269));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_268));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_14),
    .B(n_13107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_272));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1760 (.A(n_13107),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_14),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_270));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1765 (.A(n_13401),
    .B(n_14103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_264));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1766 (.B(n_12594),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_263),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_236));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1767 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_247),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_261));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1769 (.A(n_22061),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1770 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_598));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1771 (.A(n_26147),
    .B(n_7471),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_260));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_236),
    .B(n_12583),
    .C(n_12595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_253));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1782 (.A(n_10378),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1784 (.A(n_10378),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_247));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1786 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_227),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_13),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_31));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1792 (.A(n_13112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_243));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_241));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1795 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_215),
    .B(n_7469),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_240));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_207),
    .B(n_21690),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_236));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_600));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_180),
    .B(n_10379),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_226));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1814 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_196),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_227));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1817 (.A(n_13598),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1819 (.A(n_18915),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_222));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_123),
    .B(n_19108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_602));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_211));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1841 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_215));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1851 (.A(n_8739),
    .B(n_12906),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_76),
    .A2(n_21588),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_195));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1860 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_196));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_190));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1875 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_134),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_120),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_181));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_188));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_184));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_138),
    .B(n_2400),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_174));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_128),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_171));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1902 (.A(n_12905),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_163));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_36),
    .B(n_25984),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1913 (.A(n_21588),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_156));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_68),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_22));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_155));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_153));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_604));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_144));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1934 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_44),
    .B1(n_22872),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_142));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_150));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1937 (.A1(n_12903),
    .A2(n_12901),
    .B1(n_12902),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_141));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_140));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_131));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_130));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1948 (.A(n_22870),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_128));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1951 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_46),
    .B1(n_20512),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_134));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1971 (.A(n_12903),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_110));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_84));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1987 (.A(n_20504),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1988 (.A(n_20504),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1994 (.A(n_2922),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(n_3592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(n_2377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_2711),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2009 (.A(n_3479),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_80));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2014 (.A(n_2697),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_46));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2030 (.A(n_22872),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_44));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2032 (.A(n_22878),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2039 (.A(n_20504),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_56));
 AND2x4_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2056 (.A(n_3479),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[51]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_45));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[48]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_40));
 AND2x4_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[49]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2065 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_36));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_211),
    .B(n_13112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_14));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_180),
    .B(n_10379),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2076 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_11));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_6));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g20820 (.A(n_9209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_297),
    .Y(n_12276));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g2086 (.A(n_12904),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_1));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_n_92),
    .Y(n_22733));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30180 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22870));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30182 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[55]),
    .Y(n_22872));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30188 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22878));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30193 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22883));
 INVx1_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_134_55_g30259 (.A(n_11469),
    .Y(n_22949));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1743 (.A(n_7704),
    .B(n_7708),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_552));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1748 (.A(n_7709),
    .B(n_7703),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_554));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1749 (.A(n_12547),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_556));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1750 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_285),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_318),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_326));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_304),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_319),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_558));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_318),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_319));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1758 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_300),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_289),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_318));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1759 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_303),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_560));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1769 (.A(n_9616),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_307));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1772 (.A(n_14089),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_304));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1773 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_296),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_289),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_303));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1775 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_281),
    .A2(n_14688),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_301));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1776 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_266),
    .A2(n_10544),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_300));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_562));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_296));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1780 (.A(n_14089),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_292));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1783 (.A(n_12923),
    .B(n_14688),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_298));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1784 (.A(n_14091),
    .B(n_11945),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_297));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1785 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_295));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1791 (.A(n_14090),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_285));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1793 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_248),
    .B(n_4197),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_289));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1798 (.A(n_12923),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_282));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1800 (.A(n_19189),
    .B(n_12922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_281));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1803 (.A(n_10544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_278));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1806 (.A(n_19332),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_275));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_250),
    .B(n_14687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1816 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_262));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_255),
    .B(n_7452),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_266));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1818 (.A(n_7452),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_264));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1820 (.A(n_2883),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_566));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_253));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_227),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_255));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1829 (.A(n_19134),
    .B(n_7451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_254));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1830 (.A(n_19134),
    .B(n_7451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_252));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_249));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1837 (.A(n_19333),
    .B(n_19335),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_244));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1838 (.A(n_12917),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_154),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_250));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_185),
    .C(n_7453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_248));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_568));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_238));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_225));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1860 (.A(n_6742),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_230));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_181),
    .B(n_6742),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_228));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1862 (.A(n_6796),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_227));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1863 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_198),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_37));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1864 (.A(n_21497),
    .B(n_21545),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_36));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1865 (.A(n_20215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_226));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1871 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_216));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1875 (.A(n_20296),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_171),
    .C(n_12580),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_222));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1879 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_187),
    .B(n_20214),
    .C(n_3454),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_215));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_210));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1885 (.A(n_6749),
    .B(n_6799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_129),
    .B(n_19109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_570));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_201));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_199));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_198));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1906 (.A(n_18794),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1908 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_163),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_163),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_190));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_182));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_1),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_111),
    .B(n_10892),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_187));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_184));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1926 (.A(n_6799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_178));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_66),
    .C(n_13728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_20),
    .B(n_26122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_173));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1939 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_172));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1940 (.A(n_18822),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_171));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1949 (.A(n_13251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1951 (.A(n_8719),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_112),
    .C(n_8725),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_163));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1952 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_132),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_133),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_33));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1958 (.A(n_12252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_158));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_113),
    .C(n_12581),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_31));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1968 (.A(n_12578),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_93),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_29));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1970 (.A(n_12278),
    .B(n_21493),
    .C(n_11771),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_154));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_572));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_146));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1980 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_93),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_91),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_25),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_145));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_143));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_66),
    .B(n_13728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1997 (.A1(n_13239),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_138));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2002 (.A(n_13234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_128));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_80),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_127));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_119),
    .B(n_12134),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2015 (.A(n_13239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_116));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_25));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_2657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_113));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_111));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_110));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_109));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_11770),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2054 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_92));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_43),
    .B(n_4549),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_22));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g20800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_14),
    .B(n_12257),
    .Y(n_12258));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_67));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g20822 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_55),
    .Y(n_12278));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_40),
    .B(n_2747),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_n_574));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2107 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_69));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(n_12129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_66));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2111 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .B(n_2820),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(n_3375),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_62));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2116 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_20));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_59));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_47),
    .B(n_4555),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_57));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2120 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[63]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2124 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_3374),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_50));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2126 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_188),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_15));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_9),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_29),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_185),
    .B(n_7453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_12));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_112),
    .B(n_18914),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_9));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_106),
    .B(n_13240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_3));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2152 (.B(n_13234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_2),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_79));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_65),
    .B(n_13721),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_1));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21535 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(n_13231),
    .Y(n_13234));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21540 (.A(n_13231),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[58]),
    .Y(n_13239));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21541 (.A(n_13231),
    .B(u_NV_NVDLA_cmac_u_core_wt2_actv_data[62]),
    .Y(n_13240));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21552 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(n_2657),
    .Y(n_13251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21956 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[59]),
    .B(n_13707),
    .Y(n_13712));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21963 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[57]),
    .B(n_13707),
    .Y(n_13719));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21965 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[60]),
    .B(n_13707),
    .Y(n_13721));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g21972 (.A(u_NV_NVDLA_cmac_u_core_wt2_actv_data[56]),
    .B(n_3528),
    .Y(n_13728));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_g28139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_2_mul_136_55_n_101),
    .Y(n_20591));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1_reg (.CLK(nvdla_core_clk),
    .D(n_17882),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d1));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2_reg (.CLK(nvdla_core_clk),
    .D(n_4),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d2));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_2_pp_pvld_d0_d3_reg (.CLK(nvdla_core_clk),
    .D(n_5),
    .QN(u_NV_NVDLA_cmac_u_core_out_mask[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_4418),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[0]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1115),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_17868),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[11]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_23935),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[12]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_17886),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[13]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1111),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[14]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_5510),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[15]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_10329),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[16]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_22092),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[17]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_5347),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1124),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1123),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1122),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1121),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1120),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1119),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1118),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[7]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1117),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[8]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1116),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1107),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1097),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1096),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1095),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1094),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1093),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1092),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1223),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1091),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1089),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1106),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1149),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1105),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1104),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1102),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1101),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1100),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1099),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1098),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d2[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1088),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1078),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1077),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1076),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1075),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1074),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1073),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1072),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1071),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1070),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1087),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1086),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1085),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1084),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1083),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1082),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1081),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1080),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_2_sum_out_d0_d3_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1079),
    .QN(u_NV_NVDLA_cmac_u_core_out_data2[9]));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g20787 (.A(n_19530),
    .Y(n_12245));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g24385 (.A(n_16456),
    .Y(n_16458));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g24386 (.A1(n_16456),
    .A2(n_10200),
    .B(n_10202),
    .Y(n_16459));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g25773 (.A(n_17907),
    .B(n_17908),
    .Y(n_17909));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g25774 (.A(n_13687),
    .B(n_16456),
    .Y(n_17907));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g26222 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_167),
    .B(n_21170),
    .C(n_21169),
    .Y(n_18430));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g26223 (.A(n_26024),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_659),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_627),
    .Y(n_18431));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g26224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .Y(n_18432));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g30065 (.A(n_22717),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_144),
    .Y(n_22718));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6011 (.A1(n_23582),
    .A2(n_3654),
    .B(n_3685),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_500));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6013 (.A(n_23582),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_184));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6017 (.A1(n_10340),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_488),
    .B(n_2562),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_494));
 OAI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6019 (.A1(n_18828),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .B1(n_17438),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_488),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_182));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_452),
    .B(n_5457),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_181));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6023 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_488));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6024 (.A1(n_5456),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_440),
    .B(n_16459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_489));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6029 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_439),
    .B(n_16070),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_178));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6030 (.A(n_7362),
    .B(n_16069),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_483));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6033 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_481),
    .B(n_7364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_177));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_481));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6035 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_64),
    .A2(n_11541),
    .B(n_11540),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_480));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6036 (.A(n_3237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_450),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_176));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6038 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .C(n_12705),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_64));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6040 (.A(n_12706),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_453),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_175));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6044 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_446),
    .A2(n_14151),
    .B(n_14152),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_473));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6046 (.A(n_12707),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6051 (.A(n_14151),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_444),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_466));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_444),
    .B(n_4082),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_465));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6057 (.A(n_14151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_455));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_352),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_401),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_453));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6061 (.A(n_10201),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_435),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_452));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6062 (.A(n_3686),
    .B(n_3655),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_451));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6064 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_432),
    .B(n_11541),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_450));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_444),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_445));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6072 (.A1(n_23095),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_391),
    .B(n_7716),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_442));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_398),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_173));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6074 (.A(n_13688),
    .B(n_10200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_440));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6075 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_406),
    .B(n_16069),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_439));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6078 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_379),
    .B(n_6254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_437));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_408),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_404),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_436));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_418),
    .B(n_14125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_446));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_417),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_366),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_444));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6083 (.A(n_10202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_435));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6084 (.A(n_11540),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_432));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_429),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_430));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6096 (.A(n_10091),
    .B(n_14122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_429));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6101 (.A(n_10090),
    .B(n_9625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_62));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6104 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_417),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_418));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6109 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_407),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_408));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6111 (.A(n_7716),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_406));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_380),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_172));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6113 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_391),
    .B(n_23095),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_404));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6114 (.A(n_7371),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_417));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6121 (.A(n_23095),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_407));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6125 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_397));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6126 (.A(n_12701),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_384),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_396));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6127 (.A(n_13619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_354),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_401));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6128 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_357),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_400));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6130 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_358),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_356),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_398));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6136 (.A(n_18823),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_391));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6140 (.A(n_12704),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_384));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_345),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_171));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_385));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_337),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_381));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6145 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_361),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_380));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_308),
    .B(n_6257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_379));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6154 (.A(n_14125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_366));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6157 (.A(n_13412),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .C(n_13619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_372));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6165 (.A(n_9618),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_54),
    .C(n_4101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_362));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6166 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_309),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_357));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_356));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6169 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .A2(n_13412),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_322),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_354));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6170 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_307),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_344),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_361));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_326),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_359));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_261),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_327),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_358));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6176 (.A(n_20357),
    .B(n_20719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_350));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6181 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_352));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6183 (.A1(n_19112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_336),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_345));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_300),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_344));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6186 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_278),
    .B(n_5637),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_343));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_285),
    .B(n_17492),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_340));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6196 (.A(n_13412),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_330));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_337));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_258),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_328));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6201 (.A(n_19112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_327));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_283),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_326));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6203 (.A(n_19112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_336));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6212 (.A(n_14118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_329));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6213 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_324),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_325));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_321),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_322));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6222 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_311));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_279),
    .B(n_26189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_308));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_324));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6226 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_321));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6229 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_272),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_56));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_318));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6231 (.A(n_13617),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .C(n_21177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_317));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6233 (.A(n_10274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .C(n_2445),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_315));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6235 (.A(n_17808),
    .B(n_9410),
    .C(n_9408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_54));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6237 (.A(n_14118),
    .B(n_3661),
    .C(n_2312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_309));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6242 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_300));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6243 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_307));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6251 (.A(n_5637),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_298));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_294));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6257 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_288),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_52));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6262 (.A(n_8771),
    .B(n_12246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_293));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6264 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_187),
    .B(n_10271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_292));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6267 (.A(n_23835),
    .B(n_17414),
    .C(n_8772),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_288));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_285));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6271 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_44),
    .B(n_22247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_282));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6274 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_217),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_203),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_279));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6278 (.A(n_2591),
    .B(n_7379),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_278));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6279 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .A2(n_2445),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_208),
    .B2(n_2444),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_277));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6280 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_213),
    .B(n_21177),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_276));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6282 (.A(n_18431),
    .B(n_18432),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_275));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6283 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_274));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6284 (.A(n_21920),
    .B(n_22718),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_284));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6285 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_204),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_283));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6289 (.A(n_23175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_267));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6293 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_221),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_254));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6294 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_273));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6295 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_193),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_142),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_272));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6302 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_263));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6304 (.A(n_19113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_116),
    .C(n_19114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_261));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6305 (.A(n_26190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_260));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6306 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_259));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6307 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_216),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_258));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6308 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_171),
    .B(n_7097),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_256));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6309 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_255));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6312 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_143),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6314 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_248));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_251));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_237));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6339 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_229));
 AOI21xp5_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6350 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .A2(n_20784),
    .B(n_20783),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_217));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6353 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_697),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_228));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6362 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_221));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6364 (.B(n_12001),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_219),
    .A(n_19657));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6365 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_218));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6366 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_216));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6374 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_207),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6376 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_204));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6377 (.A1(n_2591),
    .A2(n_17414),
    .B1(n_2592),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_203));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6379 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_161),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6380 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_215));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6382 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_661),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_629),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_213));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6384 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_83),
    .A2(n_9074),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_44));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6385 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_631),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6389 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_209));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6390 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_657),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_625),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_207));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6391 (.A(n_18790),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_655),
    .C(n_13467),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_206));
 BUFx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6393 (.A(n_11998),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_197));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6396 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_187),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_188));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6402 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_183));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6405 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_635),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_200));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6410 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_751),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_12),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6412 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_663),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6413 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_699),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_190));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6415 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_753),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_187));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6417 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_633),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_109),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_185));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6419 (.A(n_8689),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_178));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6430 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_797),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_181));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6431 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_180),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_719));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6435 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_713),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_175));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6436 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_727),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_174));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6439 (.A(n_22712),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6441 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_725),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_168));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6442 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_755),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_167));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6444 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_729),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6448 (.A(n_12001),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_156));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6451 (.A(n_22243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_150));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6452 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_148));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6456 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_601),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_139));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6457 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_601),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_88),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_161));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6459 (.A(n_19062),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_767),
    .C(n_19056),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6465 (.A(n_16230),
    .B(n_9978),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_723),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6466 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_733),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_637),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_797),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6468 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_713),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_553),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_777),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6469 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_639),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_671),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_799),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_143));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6470 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_753),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_689),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_593),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_142));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6475 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_133));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6476 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_131));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6477 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_129));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6494 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_701),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_605),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_134));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6495 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_559),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_783),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6496 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_793),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_729),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_130));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6497 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_599),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_727),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_567),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_128));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6500 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_695),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_663),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_125));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6502 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_761),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_665),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_633),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_123));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6503 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_763),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_635),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_667),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_122));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6504 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_603),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_731),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_n_699),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_121));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6512 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_597),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_693),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_111));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6514 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_665),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_761),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_109));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6515 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_791),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_695),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_108));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6516 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_667),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_763),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_107));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6519 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_106));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6530 (.A(n_19055),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_575),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6531 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_115));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6535 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_625),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_100));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6543 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_565),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_98));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6545 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_731),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_603),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_96));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6551 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_567),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_599),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_92));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6552 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_637),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_733),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_91));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6553 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_631),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_90));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6555 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_691),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_595),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_89));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6556 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_795),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_571),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_102));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6557 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6558 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_571),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_795),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6559 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6560 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_575),
    .B(n_19055),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_85));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6562 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_651),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_619),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6563 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_669),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_765),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_82));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6585 (.A(n_23829),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_73));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6596 (.A(n_22154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_70));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6603 (.A(n_15579),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_69));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6605 (.A(n_22802),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_68));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6620 (.A(n_25598),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_343),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_35));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6621 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_317),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_34));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6622 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_33),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_272));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6629 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_206),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_26));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6630 (.A(n_26190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_250),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_25));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6632 (.A(n_7097),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_23));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6635 (.B(n_21377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_20),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_549));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6636 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_777),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_19));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6637 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_621),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_653),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_18));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6642 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_619),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_651),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_13));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6643 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_591),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_687),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_12));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6648 (.B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_783),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_7),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_559));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6650 (.A(n_22714),
    .B(n_22713),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_g6652 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_n_593),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_n_689),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_csa_tree_ADD_TC_OP_6_groupi_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_285),
    .B(n_11597),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_746));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_204),
    .B(n_11585),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_738));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_299),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_740));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2962 (.A(n_11599),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_298),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_744));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2963 (.A1(n_11583),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_299));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2964 (.A1(n_4079),
    .A2(n_11597),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_298));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_275),
    .B(n_11592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_748));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2980 (.A(n_18903),
    .B(n_24035),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_752));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_277),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_285));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2989 (.A(n_20385),
    .B(n_13437),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_23));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_277));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2992 (.A(n_20385),
    .B(n_13437),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_276));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2993 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_267),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_275));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g2998 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_239),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_270));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_265));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3003 (.A(n_11596),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_262));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_253),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_268));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3005 (.A(n_22120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_267));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3007 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_254),
    .B(n_15358),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_249),
    .B(n_26231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_259));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_240),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_251));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_250));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_254));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_253));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3026 (.A(n_5780),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_247));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3029 (.A(n_11209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_249));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3035 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_225),
    .B(n_21464),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3036 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_240));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3037 (.A(n_26191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_239));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3038 (.A(n_26191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_219),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_238));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3039 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_237));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3040 (.A(n_21464),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_236));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3042 (.A(n_20905),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_758));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3044 (.A(n_11209),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_173),
    .C(n_22113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_232));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_225));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_224));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_173),
    .B(n_22112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_223));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3056 (.A(n_10569),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3058 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_202),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_140),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3059 (.A(n_20909),
    .B(n_20912),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_218));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3060 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_760));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3065 (.A(n_10355),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_213));
 OAI21xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3072 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_197),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_204));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3074 (.A(n_21918),
    .B(n_26138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_206));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3083 (.A(n_22110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_35),
    .C(n_8035),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_202));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3085 (.A(n_19168),
    .B(n_7726),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_18));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3088 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106),
    .B(n_19115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_762));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3089 (.A(n_20904),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_182),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3090 (.A(n_11200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_192));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3091 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3092 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_165),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_190));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_189));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3094 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_197));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_109),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_188));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3101 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_152),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_167),
    .B1(n_11277),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_183));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3104 (.A(n_20903),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_182));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_43),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3116 (.A(n_8260),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_31),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_173));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3117 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_122),
    .B(n_8260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_172));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_167));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3123 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_164));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3125 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_109),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_162));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3130 (.A(n_11195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_166));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3132 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_165));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3133 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3135 (.A(n_11277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_152));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3139 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_115),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3140 (.A(n_22025),
    .B(n_22023),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_159));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3141 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_44),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_157));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_25),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_153));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_146));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_48),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_145));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_91),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_144));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_51),
    .C(n_22105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_140));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3165 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_58),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3168 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3169 (.A(n_11195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_10),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_13));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3171 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_764));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3173 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_59),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_73),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_126));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3177 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_11),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_76),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_10),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3179 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_28),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_31),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3183 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_41),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_33),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_42),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_117));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3184 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_116));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_29),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_115));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_121));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3192 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_120));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3193 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_87),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_119));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_118));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_109));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3197 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_107));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3198 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_95),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3199 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_105));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_0),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_102));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3205 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_0),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_100));
 AOI22xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3206 (.A1(n_4463),
    .A2(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B1(n_3761),
    .B2(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_98));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_766));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3212 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_11),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_77));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_10));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3216 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_73));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3221 (.A(n_3150),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3222 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_12));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(n_21183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3226 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3227 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(n_3760),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3228 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_90));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_87));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3232 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3234 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .B(n_19342),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3239 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_11));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[6]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3242 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_74));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_68));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3247 (.A(n_2325),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3249 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(n_2855),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_64));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(n_6972),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3253 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_59));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3255 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_51));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_42));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_33));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_58));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3269 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3270 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3271 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_50));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3273 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_48));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3274 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[0]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_47));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3275 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[6]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(n_2864),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3278 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[7]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3279 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3280 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(n_6965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_40));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3283 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(n_3266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_35));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[5]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_32));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[3]),
    .B(n_3148),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_31));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[0]),
    .B(n_6973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_29));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3289 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[5]),
    .B(n_19340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_28));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_3260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_27));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[2]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[1]),
    .B(n_2325),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_25));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3298 (.A(n_9549),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_5));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_3));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_71),
    .B(n_21184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_2));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[4]),
    .B(n_2337),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_122_55_n_0));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1743 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_302),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_776));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1745 (.A1(n_5065),
    .A2(n_23230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_331));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1748 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_316),
    .B(n_23230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_778));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1749 (.A(n_23236),
    .B(n_13622),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_780));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1759 (.A(n_13627),
    .B(n_5301),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_784));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1760 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_307),
    .B(n_7960),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_316));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1767 (.A(n_23220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_309));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1769 (.A(n_7531),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_307));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1774 (.A(n_5300),
    .B(n_15235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_302));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_786));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1778 (.A(n_21559),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_296));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1791 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_284),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_285));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1797 (.A(n_7749),
    .B(n_13530),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_284));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1798 (.A(n_22138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_282));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1799 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_17),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_283));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_281));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1801 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_268),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_280));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_265),
    .B(n_12717),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1803 (.A(n_21624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_278));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_234),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_271));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_268));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1814 (.A(n_12719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1815 (.A(n_21385),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_267));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_193),
    .B(n_21385),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_263));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1820 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_790));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1822 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_234),
    .B(n_2965),
    .C(n_3557),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_260));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1823 (.A(n_23195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_190),
    .C(n_3032),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_259));
 INVxp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_253));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_207),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_252));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1832 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_251));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_190),
    .B(n_21340),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_247));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1836 (.A1(n_9682),
    .A2(n_3558),
    .B1(n_2966),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_245));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_792));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_238));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1848 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_212),
    .B(n_21332),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_236));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_14),
    .B(n_20139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_234));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_229));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1860 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_230));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_228));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1863 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_198),
    .A2(n_20922),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_37));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_10),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_171),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_222));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_214));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_212));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_794));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_131),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1897 (.A(n_20922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1898 (.A(n_20916),
    .B(n_20921),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_201));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_198));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_193));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1908 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_149),
    .B(n_21573),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_192));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_5),
    .B(n_23573),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_191));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1910 (.A(n_21573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_21),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_190));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_183));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_182));
 XNOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_132),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_170));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1932 (.A(n_20917),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1934 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1937 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_50),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1940 (.A(n_20925),
    .B(n_21069),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_171));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_168));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_169));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1953 (.A(n_22837),
    .B(n_17709),
    .C(n_17707),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_158));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_155),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_156));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1964 (.A(n_20923),
    .B(n_20924),
    .C(n_21069),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_31));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1965 (.A(n_14029),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_26),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_30));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1967 (.A(n_21201),
    .B(n_21199),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_155));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1968 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_93),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_25),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_29));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_56),
    .B(n_21335),
    .C(n_13204),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_154));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1971 (.A(n_15591),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_107),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_153));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_152));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_796));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1976 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_21),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_149));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1977 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_56),
    .A2(n_13203),
    .B1(n_9350),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_148));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_146));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1980 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_93),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_91),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_25),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_145));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1982 (.A(n_14029),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_143));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1984 (.A1(n_9571),
    .A2(n_9570),
    .B(n_3206),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_151));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1986 (.A(n_26173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_140));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_139));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_138));
 XOR2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2 (.A(n_21622),
    .B(n_21626),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_788));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_134));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_133));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_132));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_128));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_126));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_116));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_25));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_123));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(n_2499),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .B(n_4521),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_115));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_110));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_108));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(n_9349),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2055 (.A(n_6576),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_92));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_43),
    .B(n_3107),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(n_14537),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2064 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_88));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_21),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_67));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2090 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_55),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_56));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2092 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_51));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_40),
    .B(n_4528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_798));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2095 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(n_15045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(n_2728),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_48));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2098 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_73));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2105 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[9]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2109 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[15]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_66));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2111 (.A(n_9349),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_62));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_46),
    .B(n_14372),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_59));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_57));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2120 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[13]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2121 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2122 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[15]),
    .B(n_3112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2123 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[14]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[11]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2124 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .B(n_3868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_50));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[8]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2137 (.A(n_21382),
    .B(n_21339),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_17));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2140 (.A(n_9677),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_29),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2142 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2143 (.A(n_23573),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_5),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_11));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2144 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_145),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_10));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_107),
    .B(n_15591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_8));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2149 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_82),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2152 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g23559 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[9]),
    .B(n_24402),
    .Y(n_15591));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g25576 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[10]),
    .B(n_9349),
    .Y(n_17707));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g25578 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[10]),
    .Y(n_17709));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g25581 (.A(n_17709),
    .B(n_22837),
    .Y(n_17710));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g30147 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[11]),
    .B(n_22834),
    .Y(n_22837));
 AND2x4_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_124_55_g30149 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[12]),
    .B(n_22834),
    .Y(n_22839));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g14562 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(n_4790));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g14563 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .Y(n_4791));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g14564 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_126),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_134),
    .C(n_18663),
    .Y(n_4793));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g14566 (.A1(n_18663),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_133),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_134),
    .B2(n_4795),
    .Y(n_4796));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g14567 (.A(n_18663),
    .Y(n_4795));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1689 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_262),
    .B(n_15962),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_712));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1694 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_271),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_714));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1695 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_716));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1696 (.A1(n_14147),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_274),
    .B(n_20868),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_282));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1700 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_268),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_273),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_270),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_278));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1701 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_264),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_718));
 AOI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1702 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_270),
    .A2(n_21552),
    .A3(n_21118),
    .B1(n_21554),
    .B2(n_21118),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_276));
 NAND3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1703 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_268),
    .B(n_21552),
    .C(n_21118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_275));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1704 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_274),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_273));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1705 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_28),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_247),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_274));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1706 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_263),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_720));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1707 (.A(n_15960),
    .B(n_21553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_271));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1708 (.A1(n_20868),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_270));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1712 (.A(n_14147),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_268));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1715 (.A1(n_4565),
    .A2(n_7188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_265));
 NAND2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1716 (.A(n_20868),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_264));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1717 (.A1(n_9480),
    .A2(n_18458),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_256),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_263));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1718 (.A(n_21118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_252),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_262));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1721 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_234),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_26),
    .B(n_12745),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_28));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_26),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_722));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1727 (.A(n_18458),
    .B(n_9480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_256));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1728 (.A(n_7188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_254));
 NOR2x1p5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1729 (.A(n_7188),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_255));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1731 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_251),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_252));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1732 (.A(n_14147),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_248));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1734 (.A(n_18458),
    .B(n_9480),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_247));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1736 (.A(n_21117),
    .B(n_21111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_251));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1742 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_232),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_243));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1743 (.A(n_12745),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_242));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1745 (.A1(n_7478),
    .A2(n_8760),
    .B(n_7479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_26));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1749 (.B(n_5910),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_239),
    .A(n_15570));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_236),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_237));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1752 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_235));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1753 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_236));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1754 (.A(n_7479),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_231));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1755 (.A(n_12744),
    .B(n_12738),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_234));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_232));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1758 (.A(n_8748),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_726));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1760 (.A(n_15570),
    .B(n_10490),
    .C(n_5903),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_229));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1761 (.A(n_21112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_164),
    .C(n_21110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_228));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1764 (.A(n_7478),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_222));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_219));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_130),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_218));
 XNOR2xp5_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1777 (.A(n_8752),
    .B(n_8759),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_213));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_728));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_196));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1799 (.A(n_20234),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_193));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1801 (.A(n_7189),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_24));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1803 (.A(n_12945),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_82),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_19),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1804 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_1),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_129),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_194));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1806 (.A(n_4796),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_191));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1809 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_105),
    .B(n_19117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_730));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_173),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1813 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_182));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_65),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_189));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1818 (.A(n_8757),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_180));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1819 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_177));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1823 (.A(n_22159),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_145),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_175));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_173));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_174));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_172));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1830 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_168));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1832 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_105),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_170));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_72),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_167));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1837 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_111),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1839 (.A(n_10346),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_78),
    .C(n_5742),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_164));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1843 (.A1(n_19829),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_128),
    .B1(n_25963),
    .B2(n_19835),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_155));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1847 (.A(n_15449),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_161));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_159));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1850 (.A(n_15796),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_6),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_158));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1853 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1857 (.A(n_23471),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_69),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_16),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_113),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_149));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1860 (.A(n_20771),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_148));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_147));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1862 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_145));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1869 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_142));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1874_dup26444 (.A(n_15796),
    .B(n_4790),
    .C(n_4791),
    .Y(n_18663));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1875 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_137));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1877 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_134));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_19));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_136));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_71),
    .B(n_15794),
    .C(n_21058),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_135));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_16),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_133));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_98),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_132));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_33),
    .B(n_12939),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_130));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1891 (.A(n_19835),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_128));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1892 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_126),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_127));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1893 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_100),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_732));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_94),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_124));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1895 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_39),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_83),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_38),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_84),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_122));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1902 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_129));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1904 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_126));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_114));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_42),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_113));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_72),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_111));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_118));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1912 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_35),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_110));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1916 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_57),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_52),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_58),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_116));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1917 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_115));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1918 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_108));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1921 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_97),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_106));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_105));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1923 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_56),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_17));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_83),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_84));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1936 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_81));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(n_5737),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1945 (.A(n_16757),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_98));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1947 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1953 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_16));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(n_16749),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1957 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_23016),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_87));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1961 (.A(n_22156),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_78));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1970 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(n_15014),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1971 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .B(n_2466),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_69));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1974 (.A(n_4386),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_68));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_58));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1981 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_48),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_49));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1984 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_38));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_66));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1987 (.A(n_2544),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_4314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_64));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_63));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_59));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1993 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[17]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_55));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_53));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_51));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2 (.A(n_8761),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_724));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2002 (.A(n_5737),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_47));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[20]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[21]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_40));
 NAND2x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .B(n_16753),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[18]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .B(n_2544),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[16]),
    .B(n_22156),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_35));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[22]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_33));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[23]),
    .B(n_2827),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_32));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_155),
    .B(n_19833),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2025 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_69),
    .B(n_23471),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2027 (.A(n_4790),
    .B(n_4791),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2029 (.A(n_15450),
    .B(n_15451),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2031 (.A(n_15794),
    .B(n_21058),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g2032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_43),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_1));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g23421 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[23]),
    .Y(n_15450));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g23422 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[18]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[22]),
    .Y(n_15451));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g23750 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[17]),
    .B(n_16757),
    .Y(n_15794));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g23753 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[19]),
    .B(n_16757),
    .Y(n_15796));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g26250 (.A(n_12746),
    .B(n_20235),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_n_150),
    .Y(n_18458));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_126_55_g26445 (.A(n_15449),
    .B(n_15450),
    .C(n_15451),
    .Y(n_18664));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1706 (.A(n_22808),
    .B(n_22805),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_674));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1707 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_269),
    .B(n_22807),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_676));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_680));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1711 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_297),
    .A2(n_9338),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_300),
    .B(n_9338),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_682));
 AOI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1720 (.A1(n_9336),
    .A2(n_20046),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278),
    .B1(n_20044),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_305));
 NAND3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1721 (.A(n_9334),
    .B(n_20046),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_304));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1725 (.A(n_21509),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_688));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1726 (.A(n_20045),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_300));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1728 (.A(n_20046),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_297));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1731 (.A(n_20045),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_295));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1735 (.A(n_11968),
    .B(n_11965),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_293));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1736 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_292));
 AO21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1738 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_262),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_32),
    .B(n_21984),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_290));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_268),
    .B(n_3817),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_690));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1740 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_286),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_287));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1743 (.A(n_9483),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_271),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_286));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1747 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_280));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1748 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_692));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_265),
    .B(n_8387),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_279));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1752 (.A(n_8387),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_278));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_274));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1755 (.A(n_9481),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_271));
 NOR2xp67_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_269));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_242),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_16),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_273));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_268));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_265));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1765 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_12),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_264));
 OAI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1767 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_247),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_31),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_32));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_261));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1769 (.A(n_21984),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1770 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_227),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_694));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1771 (.A(n_21983),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_243),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_260));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1774 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_255));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1775 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_192),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_257));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_190),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_254));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1780 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_12),
    .B(n_4403),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_252));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1782 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_208),
    .B(n_19816),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_249));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1783 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_247),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_248));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1784 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_208),
    .B(n_19816),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_247));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1786 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_227),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_13),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_31));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1790 (.A1(n_8376),
    .A2(n_19746),
    .B1(n_4404),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_28),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1793 (.A(n_20400),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_5),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_242));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1794 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_13),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1796 (.A(n_20900),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1803 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_196),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_696));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1806 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_216),
    .B(n_19809),
    .C(n_19810),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_231));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1807 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_230));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1810 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_180),
    .B(n_26110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_229));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1814 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_196),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_227));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_30));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1821 (.A(n_19746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_28));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_77),
    .C(n_20421),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_225));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1827 (.A(n_20901),
    .B(n_20896),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_223));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1833 (.A(n_19815),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_216));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_698));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_212));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_211));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1843 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_205),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_206));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1848 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_173),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_186),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_172),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_202));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1850 (.A(n_19737),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_121),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_208));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1852 (.A(n_22064),
    .B(n_20395),
    .C(n_20397),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_205));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_200));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1856 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_179),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_77),
    .B2(n_20422),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_195));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1860 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_196));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_193));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1866 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_130),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_192));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1867 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_4),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_118),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_191));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1868 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_167),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_190));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_186));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1873 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_183));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1874 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_118),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_149),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_117),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_182));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1884 (.A(n_20895),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_176));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_179));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_177));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1895 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_136),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1896 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_172));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_169));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1904 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_170));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1905 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_113),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_36),
    .B(n_25990),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_20),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_160));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_93),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_99),
    .C(n_21991),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1922 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_81),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_103),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_157));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1928 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_4),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_149));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_700));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1930 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_68),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_41),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_69),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_146));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_144));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1933 (.A1(n_21991),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_79),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_143));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1940 (.A1(n_21987),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_71),
    .B(n_21988),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_148));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_131));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1946 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_130));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_128));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1949 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_89),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_80),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_127));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1950 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_126));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_137));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1954 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_52),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_53),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_136));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_134));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_124));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1959 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_72),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_123));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_119));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1964 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_117),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_118));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1974 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_93));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_84));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1982 (.A(n_21991),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_79));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(n_2958),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_112));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(n_14981),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_14179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1998 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_21));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_98));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_293),
    .B(n_21508),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_686));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(n_14984),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2003 (.A(n_12800),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(n_14186),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_91));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_2392),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_82));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2011 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_80));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2014 (.A(n_2381),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2015 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(n_12800),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_69));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2022 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_59));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2024 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_52),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_53));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_46));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2030 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_43),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_44));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2032 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_41),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_3331),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_68));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(n_14985),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_65));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[24]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(n_2307),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(n_2944),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2049 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[25]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_52));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[28]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(n_2293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[31]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(n_2381),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(n_19645),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[26]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[30]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2058 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[31]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_43));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2059 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[30]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[24]),
    .B(n_3491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_40));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2061 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[26]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_39));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .B(n_3504),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_38));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[25]),
    .B(n_14183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2065 (.A(n_14975),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[29]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[27]),
    .B(n_14179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_35));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2071 (.A(n_10085),
    .B(n_21985),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_16));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_14));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_180),
    .B(n_26110),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_13));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2075 (.A(n_19985),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_5),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_10));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_40),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2082 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_127),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_5));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2083 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_4));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g2085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_64),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_100),
    .Y(n_20395));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28002 (.A(n_20396),
    .Y(n_20397));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_75),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_67),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_n_35),
    .Y(n_20396));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28004 (.A(n_22064),
    .B(n_20399),
    .Y(n_20400));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28005 (.A1(n_20395),
    .A2(n_20396),
    .B1(n_20397),
    .B2(n_20398),
    .Y(n_20399));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_128_55_g28006 (.A(n_20395),
    .Y(n_20398));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_297),
    .B(n_19175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_654));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2960 (.A(n_18970),
    .B(n_12036),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_648));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_285),
    .B(n_13634),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_646));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_298),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_312),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_652));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2971 (.A1(n_10348),
    .A2(n_19175),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_291),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_312));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2975 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_280),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_294),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_656));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2989 (.A(n_10954),
    .B(n_17560),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_298));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_290),
    .B(n_10348),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_297));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2992 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_262),
    .A2(n_9866),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_261),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_295));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2993 (.A1(n_9506),
    .A2(n_10902),
    .B(n_9507),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_294));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2994 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_271),
    .B(n_4408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_658));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_291));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_262),
    .B(n_9865),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_286));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g2999 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_274),
    .B(n_9865),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_285));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3003 (.A(n_19543),
    .B(n_10904),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_660));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_278),
    .B(n_10492),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_280));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3009 (.A(n_9503),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_278));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3010 (.A(n_9866),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_274));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3013 (.A(n_9501),
    .B(n_9506),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_271));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3020 (.A(n_9281),
    .B(n_7925),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_269));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3024 (.A(n_22021),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_208),
    .C(n_5719),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_265));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_263));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3027 (.A(n_26194),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_262));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3028 (.A(n_26194),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_261));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3034 (.A(n_19540),
    .B(n_26193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_662));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3035 (.A(n_22022),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_255));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3037 (.A(n_14868),
    .B(n_19200),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_224),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_253));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3040 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_210),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_239),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_250));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_247));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_10),
    .B(n_21612),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_221),
    .B(n_21607),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_242));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3049 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_241));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3050 (.A(n_21612),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_7),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_240));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_178),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_215),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_664));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3053 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_9),
    .B(n_9821),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3055 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_191),
    .B(n_23112),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_238));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3070 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_195),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3079 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_171),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_46),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_220));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120),
    .B(n_19120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_666));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3086 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_215));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3089 (.A(n_21607),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_212));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3092 (.A(n_21613),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_208));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_172),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_119),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_209));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3105 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_200));
 NOR2xp33_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3107 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_199));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3108 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3110 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_46),
    .A2(n_20377),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_45),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_195));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_87),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_193));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3113 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_129),
    .A2(n_13023),
    .B1(n_13021),
    .B2(n_13022),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_188));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3115 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_155),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_116),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_191));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_164),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_178));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_119),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_176));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_185));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_73),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_175));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3136 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3138 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_127),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_172));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3140 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_63),
    .B(n_26140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_171));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3143 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_168));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3144 (.A(n_3239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_77),
    .C(n_9819),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_167));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3146 (.A(n_20377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_162));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_160));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_51),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_133),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_164));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3155 (.A(n_4671),
    .B(n_5137),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_155));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3166 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_39),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_18),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_150));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3167 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_108),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3169 (.A(n_12930),
    .B(n_12932),
    .C(n_12935),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_145));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_142));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_668));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_136));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_96),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_141));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3187 (.A(n_13021),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_129));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3188 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_108),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_127));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_133));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3192 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_33),
    .A2(n_5137),
    .B1(n_4671),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_124));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3194 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_123));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_73),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_42),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_122));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3196 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_99),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_61),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_100),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_131));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_105),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_53),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_54),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3200 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_121));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_120));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_118));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3210 (.A(n_7265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_113));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .A2(n_3168),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .B2(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_110));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_107));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_105));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3223 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_92));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3230 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_108));
 NAND2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_103));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_99));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3242 (.A(n_3218),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3243 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3247 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .B(n_18039),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_93));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_91));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3250 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_87));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3253 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_84));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3254 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(n_22743),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_83));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_81));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_79));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3260 (.A(n_18039),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3261 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .B(n_15192),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_73));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_70),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_670));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3266 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_67),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_66));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_64));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_61));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_54));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_47),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_48));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3277 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_46),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_45));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3283 (.A(n_9273),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .B(n_3168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_70));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_68));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3287 (.A(n_22743),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_65));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3289 (.A(n_15192),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3290 (.A(n_3181),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[33]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_59));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(n_3218),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_56));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(n_3396),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_51));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[32]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[38]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_49));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3303 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(n_4123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_46));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[35]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_43));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3306 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[32]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_42));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3308 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[37]),
    .B(n_3214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_39));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[38]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_38));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3310 (.A(n_15201),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[39]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3311 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[33]),
    .B(n_18031),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_36));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[36]),
    .B(n_9273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3313 (.A(n_4826),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[34]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_7),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3323 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_9));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_7));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3326 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_18),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_39),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_6));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_79),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_g3330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_130_55_n_2));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_299),
    .B(n_6030),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_622));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22028 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(n_16763),
    .Y(n_13784));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22030 (.A(n_16763),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .Y(n_13786));
 NAND2x1p5_ASAP7_75t_R u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22032 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(n_16772),
    .Y(n_13788));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22033 (.A(n_16769),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .Y(n_13789));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22037 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .B(n_16763),
    .Y(n_13793));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g22041 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .B(n_16772),
    .Y(n_13797));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_319),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_610));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2960 (.A(n_21391),
    .B(n_13016),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_616));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2962 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_288),
    .A2(n_13522),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_319));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_309),
    .B(n_4410),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_618));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_300),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_314),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_620));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2971 (.A1(n_14135),
    .A2(n_6030),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_314));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2975 (.A(n_6031),
    .B(n_6033),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_624));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2976 (.A(n_21392),
    .B(n_13012),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_310));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_303),
    .B(n_13013),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_309));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2986 (.A(n_13015),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_303));
 NOR2xp33_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2989 (.A(n_23103),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_300));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_292),
    .B(n_14135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_299));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2992 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_264),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_277),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_263),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_297));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2995 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_292),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_293));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2996 (.A(n_14136),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_292));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g29963 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(n_22616),
    .Y(n_22617));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g29968 (.A(n_22616),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .Y(n_22621));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2997 (.A(n_23102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_290));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g29971 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .B(n_22616),
    .Y(n_22624));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g29977 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B(n_22616),
    .Y(n_22630));
 OR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2998 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_264),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_288));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g29983 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(n_22616),
    .Y(n_22636));
 NOR2x1_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g2999 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_276),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_275),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_287));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_251),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_259),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_628));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3010 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_277),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_276));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3016 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_249),
    .B(n_11644),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_277));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3017 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_249),
    .B(n_11644),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_275));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3026 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_265));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3027 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_264));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_263));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3032 (.A(n_18165),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3034 (.A(n_21084),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_630));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3038 (.A(n_18167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_254));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3041 (.A(n_18166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_251));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3043 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_249));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3047 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_10),
    .B(n_22100),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_245));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3048 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_221),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_244));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3049 (.A(n_22101),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_243));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3052 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_176),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_632));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3054 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_231),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_237));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3060 (.A(n_26035),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_182),
    .C(n_20223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_234));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3063 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_229),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_230));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3064 (.A(n_21083),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_228));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3066 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_231));
 NOR2xp67_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3067 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_173),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_208),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_229));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3068 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_70),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_191),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_225));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3071 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_149),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_24));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3072 (.A(n_19249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_224));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_220),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_221));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3079 (.A(n_20931),
    .B(n_20933),
    .C(n_20934),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_220));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3080 (.A(n_9685),
    .B(n_24678),
    .C(n_19644),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_219));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3084 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118),
    .B(n_19122),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_634));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_191),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_217));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3086 (.A(n_21082),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_198),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_214));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3089 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_211));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3096 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_170),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_117),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3098 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_174),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_208));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3105 (.A(n_21078),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_198));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3109 (.A1(n_26267),
    .A2(n_4230),
    .B1(n_4231),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_194));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3112 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_158),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_85),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_36),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_191));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3114 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_190));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3119 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_182));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3120 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_180));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3121 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_162),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_176));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3124 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_117),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_128),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_174));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3126 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_183));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3127 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_181));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3128 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_135),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3134 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_71),
    .C(n_22630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_173));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3138 (.A(n_22636),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_125),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_170));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_157),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_158));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3151 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_49),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_131),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_162));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3153 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_35),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3155 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_90),
    .B(n_13697),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_32),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_154));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3156 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_33),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_62),
    .C(n_13793),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_153));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3164 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_46),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_47),
    .C(n_13789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_151));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3166 (.A(n_20675),
    .B(n_20674),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_63),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_149));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3167 (.A(n_13786),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_106),
    .C(n_22636),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_147));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3169 (.A(n_23659),
    .B(n_23658),
    .C(n_23660),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_143));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3170 (.A(n_18760),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_88),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_21));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3172 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_139),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_140));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3174 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_108),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_636));
 AOI22xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3179 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_92),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_100),
    .B1(n_13797),
    .B2(n_22624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_135));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3180 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_134));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3181 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_88),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_72),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_17),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_133));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3182 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_64),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_46),
    .B1(n_13789),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_132));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3185 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_104),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_139));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3188 (.A(n_13786),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_106),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_125));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3190 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_36),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_123));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3191 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_96),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_131));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3195 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_71),
    .B(n_22630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_120));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3196 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_97),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_59),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_98),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_129));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3198 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_103),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_51),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_52),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_128));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3201 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_68),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_49),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_118));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3202 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_117));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3204 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3207 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_20),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_114));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3213 (.A1(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .A2(n_18049),
    .B1(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B2(n_23276),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_108));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3214 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_104),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_105));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3215 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_102),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_103));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3216 (.A(n_13797),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_100));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3217 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_98));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3223 (.A(n_22624),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_92));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3224 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_89),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_90));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3225 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_87),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_88));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3233 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_17),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_72));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3235 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_106));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3236 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_104));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3237 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_102));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3238 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_101));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g32386 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_114),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_139),
    .Y(n_25299));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3240 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_97));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3241 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_20));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3242 (.A(n_3309),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3243 (.A(n_2985),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3244 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_94));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3246 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3248 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3249 (.A(n_19391),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_87));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3250 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(n_3713),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3251 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3252 (.A(n_3317),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3256 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(n_3706),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3257 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_79));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3258 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_78));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3259 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[45]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3262 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_73));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3263 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_17));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3264 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(n_3309),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_71));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3265 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_68),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_638));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3266 (.A(n_13789),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_64));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3267 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_62));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3268 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_58),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_59));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3272 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_51),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_52));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3276 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3282 (.A(n_13784),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_32));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3283 (.A(n_19396),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_70));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3284 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[40]),
    .B(n_18049),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_68));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3285 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_67));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3286 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3288 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_63));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3289 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_61));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3290 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3291 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3292 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[41]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_57));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3294 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .B(n_3317),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3295 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3296 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3298 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[41]),
    .B(n_23280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_49));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3299 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[40]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_15));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3300 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[45]),
    .B(n_19393),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3301 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(n_9154),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3302 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[42]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3305 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[43]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_41));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3309 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[46]),
    .B(n_19395),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_36));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3310 (.A(n_3713),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[47]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_35));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3312 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[44]),
    .B(n_19391),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_33));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3322 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_7),
    .B(n_3615),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_10));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3325 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_3),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_7));
 XOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3328 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_79),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_4),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_54));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3329 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_77),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_3));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3330 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_53),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_2));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_g3331 (.A(n_13793),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_33),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_132_55_n_1));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1708 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_292),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_584));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1711 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_297),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_306),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_295),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_313));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1713 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_300),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_306),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_586));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1718 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_296),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_303),
    .B(n_21477),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_306));
 AOI321xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1720 (.A1(n_21477),
    .A2(n_21426),
    .A3(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278),
    .B1(n_21429),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_305));
 NAND3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1721 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_296),
    .B(n_21426),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_304));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1722 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_303));
 AOI21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1724 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_267),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_290),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1725 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_275),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_290),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_592));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1726 (.A(n_21430),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_297),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_300));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1728 (.A(n_21426),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_297));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1730 (.A(n_7491),
    .B(n_20680),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_296));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1731 (.A(n_21430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_295));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1735 (.A(n_21474),
    .B(n_7491),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_293));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1736 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_280),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_292));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1738 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_262),
    .A2(n_22567),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_290));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1739 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_268),
    .B(n_3893),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_594));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1747 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_279),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_280));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1748 (.A(n_2789),
    .B(n_22565),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_596));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1750 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_274),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_275));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1751 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_279));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1752 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_266),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_265),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_278));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1754 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_273),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_274));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1756 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_261),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_257),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_269));
 NOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1757 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_242),
    .B(n_7493),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_273));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1758 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_259),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_262),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_268));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1762 (.A(n_7493),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_242),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_267));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1763 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_239),
    .B(n_19135),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_233),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_266));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1764 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_223),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_15),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_265));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1768 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_260),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_261));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1769 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_258),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_259));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1770 (.A(n_21980),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_241),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_598));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1771 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_246),
    .B(n_22568),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_262));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1772 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_243),
    .B(n_19123),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_260));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1773 (.A(n_22568),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_246),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_258));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1775 (.A(n_19123),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_243),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_257));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1777 (.A(n_19135),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_250));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1778 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_224),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_190),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_254));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1780 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_12),
    .B(n_11121),
    .C(n_9231),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_252));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1783 (.A(n_22566),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_248));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1786 (.A1(n_21980),
    .A2(n_26166),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_31));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1787 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_10),
    .B(n_22779),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_246));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1792 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_164),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_243));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1793 (.A(n_22779),
    .B(n_21618),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_242));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1794 (.A(n_23083),
    .B(n_26166),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_241));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1796 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_239));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1797 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_238));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1800 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_207),
    .B(n_19137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_236));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1803 (.A(n_8975),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_212),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_600));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1804 (.A(n_6896),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_233));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1807 (.A(n_23083),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_230));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1812 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_193),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_217),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_226));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1815 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_195),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_185),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_30));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_223),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_224));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1826 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_185),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_77),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_225));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1827 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_197),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_176),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_223));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1834 (.A(n_8973),
    .B(n_19124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_602));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1835 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_213));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1836 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_200),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_212));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1838 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_70),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_193),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_217));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1839 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_164),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_211));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1848 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_173),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_186),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_172),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_202));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1849 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_153),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_201));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1851 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_148),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_166),
    .C(n_11359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_207));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1854 (.A(n_21979),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_199));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1855 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_200));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1857 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_76),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_23),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_77),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_158),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_195));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1859 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_145),
    .B(n_6902),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_197));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1865 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_96),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_50),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1868 (.A(n_6902),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_90),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_190));
 INVx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1872 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_186));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1880 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_56),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_144),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_185));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_140),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_184));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_175),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_176));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1886 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_172),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_173));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_138),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_37),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1890 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_131),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_179));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1893 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_35),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_177));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1894 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_175));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1895 (.A(n_20928),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_40),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1896 (.A(n_18827),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_172));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1899 (.A(n_10908),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_166));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1909 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_83),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_56),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_164));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1911 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1913 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_23),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_158));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1919 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_57),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1920 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_78),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_99),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_23));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1924 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_88),
    .B(n_9472),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_91),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_154));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_85),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_51),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_44),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_153));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1929 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_112),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_72),
    .B(n_8973),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_604));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_90),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_38),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_145));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1932 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_82),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_95),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_83),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_94),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_144));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1933 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_78),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_92),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_79),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_93),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_143));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1934 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_84),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_44),
    .B1(n_22871),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_142));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1935 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_19),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_18),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_150));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1938 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_47),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_97),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_140));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1940 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_114),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_115),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_148));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_137),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_138));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1943 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_135));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1944 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_132),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_133));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1945 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_37),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_86),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_131));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1948 (.A(n_22875),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_128));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1952 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_139));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1953 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_106),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_60),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_105),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_137));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1955 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_63),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_65),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_62),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_134));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_100),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_132));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1960 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_101),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_54),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_122));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1961 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_121),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1962 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_106),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_61),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_121));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1963 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_63),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_66),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_119));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1967 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_55),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_111),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_116));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1969 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_71),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_114),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_115));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1973 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_106));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1976 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_95),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_94));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1977 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_92),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_93));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1978 (.A(n_9470),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_88));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_84));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1980 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_82),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_83));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_78),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_79));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1983 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_77));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1986 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_114));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_113));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1988 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_112));
 NAND2x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1989 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_111));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1992 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1994 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(n_2922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_102));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1995 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_3190),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_101));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1996 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_100));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1997 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g1999 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_98));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_293),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_302),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_590));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(n_3592),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_97));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_96));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2002 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_95));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(n_3474),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_92));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(n_22865),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_91));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(n_2377),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_2711),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_89));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2008 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_3468),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2009 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(n_3479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_85));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2010 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_82));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2012 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_80));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2013 (.A(n_2922),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_78));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2014 (.A(n_2697),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_76));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2015 (.A(n_3468),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2016 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2019 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_65),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_66));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2020 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_63));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2021 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_60),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_61));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2028 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_45),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_46));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2030 (.A(n_22871),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_44));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_3408),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_72));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2036 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_70));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_68));
 NAND2x1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_67));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2040 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_65));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2041 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2042 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2043 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[48]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_60));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2045 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(n_2359),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_56));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[49]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_55));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2048 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(n_20459),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2050 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[53]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_51));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2051 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(n_2364),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_50));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_20));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2053 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[55]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_19));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2055 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[54]),
    .B(n_2697),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_47));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .B(n_3479),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_45));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[54]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_18));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2060 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[48]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_40));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .B(n_3591),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_38));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2063 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[49]),
    .B(n_22886),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_37));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2065 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .B(n_2927),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_36));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2066 (.A(n_22886),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[51]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_35));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2072 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_190),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_15));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_211),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_225),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_14));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2075 (.A(n_19253),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_202),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_12));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2076 (.A(n_22258),
    .B(n_26153),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_11));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_174),
    .B(n_21617),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_10));
 XNOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2080 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_150),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_116),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_7));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2081 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_40),
    .B(n_20928),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_6));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2084_dup26446 (.A(n_22874),
    .B(n_13319),
    .Y(n_18665));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g2085 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_67),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_2));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g21624 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_102),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_46),
    .B1(n_12154),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_n_45),
    .Y(n_13319));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g30181 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[55]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22871));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g30184 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[52]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .Y(n_22874));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_134_55_g30185 (.A(u_NV_NVDLA_cmac_u_core_dat0_actv_data[50]),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[53]),
    .Y(n_22875));
 A2O1A1O1Ixp25_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1740 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_298),
    .A2(n_14140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_301),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_211),
    .D(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_544));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1741 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_225),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_330),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_546));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1743 (.A(n_6017),
    .B(n_21699),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_552));
 AO21x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1746 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_298),
    .A2(n_14140),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_301),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_330));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1767 (.A(n_11343),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_309));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1772 (.A(n_19254),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_285),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_304));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1775 (.A1(n_20653),
    .A2(n_20639),
    .B(n_20660),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_301));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1777 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_279),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_278),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_562));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1779 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_293),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_294));
 INVxp67_ASAP7_75t_SRAM u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1780 (.A(n_19254),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_292));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1783 (.A(n_20659),
    .B(n_20639),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_298));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1786 (.A(n_20653),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_282),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_293));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1790 (.A(n_9992),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_286));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1791 (.A(n_7947),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_285));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1798 (.A(n_20659),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_282));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1802 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_265),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_266),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_279));
 HB1xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1803 (.A(n_11267),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_278));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1806 (.A(n_12715),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_244),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_275));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1810 (.A(n_9142),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_245),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_271));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1814 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_264),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_265));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1817 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_255),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_266));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1818 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_237),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_255),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_264));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1820 (.A(n_2887),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_238),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_566));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1822 (.A(n_9142),
    .B(n_3516),
    .C(n_3922),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_260));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1824 (.A1(n_12715),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_239),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_240),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_258));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1828 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_12),
    .B(n_25431),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_255));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1832 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_37),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_230),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_251));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1833 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_248),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_249));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1834 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_190),
    .B(n_25313),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_247));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1836 (.A1(n_26167),
    .A2(n_3923),
    .B1(n_3516),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_222),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_245));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1837 (.A(n_21424),
    .B(n_25430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_244));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1838 (.A(n_20765),
    .B(n_21395),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_250));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1839 (.A(n_25431),
    .B(n_11116),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_248));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1842 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_198),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_210),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_568));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1843 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_205),
    .B(n_25430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_240));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1844 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_205),
    .B(n_25430),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_239));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1845 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_229),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_230),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_238));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1847 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_212),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_153),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_178),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_237));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1854 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_229));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1859 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_194),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_213),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_225));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1860 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_214),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_181),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_230));
 NOR2xp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1861 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_181),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_214),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_228));
 OAI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1863 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_198),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_199),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_37));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1875 (.A(n_21422),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_171),
    .C(n_21505),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_222));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1881 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_211));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1882 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_200),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_201),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_210));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1883 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_182),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_179),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_214));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1884 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_84),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_194),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_213));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1885 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_153),
    .B(n_9929),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_209));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1886 (.A(n_21395),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_184),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_208));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1887 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_134),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_170),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_212));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1888 (.A(n_21424),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_205));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1889 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_183),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_570));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1897 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_199),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_200));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1898 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_201));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1899 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_125),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_180),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_199));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1903 (.A1(one_),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_129),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_198));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1906 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_160),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_53),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_98),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_194));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1907 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_146),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_193));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1910 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_163),
    .B(n_22020),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_190));
 NAND2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1916 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_169),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_168),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_183));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1918 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_130),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_139),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_131),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_182));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1925 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_110),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_143),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_184));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1926 (.A(n_9929),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_178));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1931 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_50),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_2),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_170));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1932 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_141),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_66),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_181));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1933 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_137),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_141),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_180));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1934 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_88),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_8),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_179));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1937 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_2),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_50),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_134),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_174));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1940 (.A(n_19754),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_105),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_171));
 INVxp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1941 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_167),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_168));
 NAND2xp5_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1948 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_142),
    .B(n_13249),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_169));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1949 (.A(n_13249),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_142),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_167));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1951 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_54),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_112),
    .C(n_5948),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_163));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1956 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_159),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_160));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1958 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_158));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1959 (.A(n_20993),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_157));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1965 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_110),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_159));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1966 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_62),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_26),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_57),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_30));
 MAJx2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1968 (.A(n_13233),
    .B(n_20006),
    .C(n_9818),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_29));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1971 (.A(n_13716),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_107),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_88),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_153));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1972 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_151),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_152));
 AOI21xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1974 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_124),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_129),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_572));
 OAI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1976 (.A1(n_22020),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_71),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_67),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_22),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_149));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1979 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_98),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_53),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_146));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1982 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_58),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_64),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_143));
 OA21x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1984 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_23),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_83),
    .B(n_19821),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_151));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1987 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_138),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_139));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1990 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_66),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_90),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_137));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1991 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_48),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_119),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_142));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1997 (.A1(n_13237),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_75),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_116),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_76),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_141));
 AOI22xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g1999 (.A1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_120),
    .A2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_74),
    .B1(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_121),
    .B2(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_138));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2 (.A(n_11264),
    .B(n_11268),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_564));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2000 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_121),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_74),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_134));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2001 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_133));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2003 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_130),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_131));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2004 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_130));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2005 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_122),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_129));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2006 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_99),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_59),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_128));
 NOR3xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2013 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_119),
    .B(n_12134),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_40),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_125));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2014 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_120),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_121));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2015 (.A(n_13237),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_116));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2026 (.A(n_13711),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_95));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2034 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_85),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_86));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2035 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_124));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2037 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(n_2657),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_122));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2038 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_120));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2039 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(n_2746),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_119));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2044 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(n_22019),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_112));
 NAND2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2046 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_26));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2047 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_110));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2050 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_107));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2052 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_105));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2056 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_99));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2057 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[62]),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_98));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2062 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(n_3528),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_90));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2064 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(n_12124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_88));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2066 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_85));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2073 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_75),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_76));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2074 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_73),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_74));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2077 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_71),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_22));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2082 (.A(n_22020),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_67));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2093 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_40),
    .B(n_2747),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_n_574));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2094 (.A(n_2820),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_23));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2095 (.A(n_4263),
    .B(n_3630),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_84));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2096 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_83));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2097 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(n_12124),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_48));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2100 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(n_13228),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_80));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2101 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2103 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_75));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2104 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_73));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2106 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_71));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2110 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_66));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2112 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[63]),
    .B(n_3375),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_64));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2114 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[61]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_62));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2117 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_59));
 NOR2xp33_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2118 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_47),
    .B(n_4555),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_58));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2119 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[61]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_57));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2121 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[62]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_54));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2122 (.A(n_4263),
    .B(n_4553),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_53));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2124 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .B(n_3374),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_50));
 INVx1_ASAP7_75t_L u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2126 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_46));
 INVx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2129 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_43));
 INVxp67_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2136 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[56]),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_40));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2142 (.A(n_11116),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_174),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_12));
 XOR2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2145 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_112),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_7),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_9));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2146 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_107),
    .B(n_13716),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_8));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2147 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_54),
    .B(n_5948),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_7));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2148 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_59),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_99),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_6));
 XNOR2x1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2152 (.B(n_13235),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_2),
    .A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_79));
 AND2x2_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g21536 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .B(n_13231),
    .Y(n_13235));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g21538 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(n_13231),
    .Y(n_13237));
 XNOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g2154 (.A(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_57),
    .B(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_62),
    .Y(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_0));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g21550 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(n_2657),
    .Y(n_13249));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g21955 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .B(n_13707),
    .Y(n_13711));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g21959 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[57]),
    .B(n_3528),
    .Y(n_13716));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g32504 (.A(n_11770),
    .B(u_NV_NVDLA_cmac_u_core_wt3_actv_data[58]),
    .Y(n_25425));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g32505 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[59]),
    .B(n_13707),
    .Y(n_25426));
 NAND2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g32506 (.A(u_NV_NVDLA_cmac_u_core_wt3_actv_data[60]),
    .B(u_NV_NVDLA_cmac_u_core_dat0_actv_data[58]),
    .Y(n_25427));
 MAJIxp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g32507 (.A(n_25429),
    .B(n_22524),
    .C(u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_n_157),
    .Y(n_25430));
 XOR2xp5_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_mul_136_55_g32509 (.A(n_25427),
    .B(n_25426),
    .Y(n_25428));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1_reg (.CLK(nvdla_core_clk),
    .D(n_17876),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d1));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2_reg (.CLK(nvdla_core_clk),
    .D(n_18),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d2));
 DFFHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_mac_3_pp_pvld_d0_d3_reg (.CLK(nvdla_core_clk),
    .D(n_12),
    .QN(u_NV_NVDLA_cmac_u_core_out_mask[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_4419),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[0]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_17910),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[10]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1059),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[11]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1058),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[12]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_17880),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1056),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[14]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_5444),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[15]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_5454),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[16]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_6044),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[17]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_21197),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1068),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1067),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1264),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1066),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1065),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1064),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1063),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1061),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[8]));
 DFFHQNx2_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_16536),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1050),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1277),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1040),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1039),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1038),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1037),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1036),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1035),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1034),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1032),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1049),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1048),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1047),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1046),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1045),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1044),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1043),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1042),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1276),
    .QN(u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d2[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1031),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_992),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1020),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1019),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1018),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1017),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1016),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1015),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1014),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1013),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1030),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1029),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1028),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1027),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1026),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1024),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1023),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1022),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_mac_3_sum_out_d0_d3_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1021),
    .QN(u_NV_NVDLA_cmac_u_core_out_data3[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1587),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1586),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1585),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1584),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1471),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1583),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1582),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1581),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1439),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1438),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1437),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1362),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1436),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1435),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1434),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1433),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data0[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1579),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1578),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1577),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1576),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1575),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1574),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1573),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1572),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1432),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1430),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1429),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1428),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1427),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1425),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1424),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data1_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1423),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1570),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1569),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1568),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1567),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1566),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1565),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1564),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1563),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1421),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1420),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1419),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1418),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1417),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1416),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1453),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data2_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1414),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1562),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1561),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1560),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1559),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1558),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1557),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1556),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1555),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1598),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1411),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1409),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1408),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1407),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1406),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1405),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data3_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1404),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data3[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1554),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1553),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1552),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1595),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1551),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1550),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1548),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1547),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1402),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1401),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1400),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1399),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1398),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1397),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1396),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data4_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1395),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data4[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1545),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1544),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1543),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1542),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1596),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1541),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1540),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1539),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1394),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1393),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1392),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1390),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1389),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1452),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1387),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data5_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1386),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data5[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1537),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1536),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1535),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1534),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1533),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1532),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1531),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1530),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1383),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1330),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1381),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1380),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1379),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1378),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1377),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data6_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1375),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data6[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1529),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1528),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1527),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1526),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1589),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1525),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1524),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1523),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1373),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1371),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1369),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1368),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1367),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1366),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1447),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_data7_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1448),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_data7[7]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1607),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1606),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1605),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1604),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1603),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1602),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1601),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1600),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d1[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2063),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2062),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2061),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2060),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2059),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2058),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2057),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_mask_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2056),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_mask[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2055),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2054),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2053),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2052),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2051),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2050),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2049),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2048),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_2047),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d1[8]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2046),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2045),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2044),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2043),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2042),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2041),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_stripe_st),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2040),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_stripe_end),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2039),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_2038),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pd_d2[8]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1_reg (.CLK(nvdla_core_clk),
    .D(n_2126),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d1),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_dat_pvld_d2_reg (.CLK(nvdla_core_clk),
    .D(n_2132),
    .QN(u_NV_NVDLA_cmac_u_core_in_dat_pvld),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1522),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1597),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1521),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1520),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1519),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1518),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1517),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1516),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1361),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1360),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1359),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1358),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1357),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1356),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1355),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1315),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data0[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1514),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1513),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1512),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1470),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1511),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1510),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1509),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1508),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1354),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1316),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1353),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1352),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1351),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1350),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1349),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data1_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1317),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1505),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1504),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1503),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1502),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1501),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1500),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1499),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1498),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1347),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1346),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1345),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1344),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1342),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1341),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1340),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data2_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1325),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1497),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1496),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1495),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1494),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1493),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1492),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1491),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1490),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1338),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1335),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1337),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1336),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1339),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1343),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1348),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data3_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1334),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data3[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1489),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1506),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1507),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1488),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1515),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1487),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1486),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1485),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1403),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1370),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1374),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1441),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1333),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1332),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1382),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data4_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1384),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data4[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1484),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1538),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1483),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1482),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1546),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1549),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1481),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1480),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1410),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1413),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1331),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1329),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1415),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1431),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1422),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data5_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1426),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data5[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1571),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1479),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1478),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1594),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1580),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1477),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1476),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1588),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1440),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1328),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1327),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1326),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1324),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1323),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1442),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data6_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1322),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data6[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1475),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1474),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1592),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1590),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1591),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1473),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1472),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1593),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1321),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1445),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1443),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1320),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1444),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1319),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1446),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_data7_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1318),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_data7[7]));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1615),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1614),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1613),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1612),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1611),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1610),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1609),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1608),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d1[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2079),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2078),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2077),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2076),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_2075),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_2074),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_2073),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_mask_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_2072),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_mask[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1_reg (.CLK(nvdla_core_clk),
    .D(n_2125),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d1),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_pvld_d2_reg (.CLK(nvdla_core_clk),
    .D(n_2133),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_pvld),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2071),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2070),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2069),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2068),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2067),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_sel[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2066),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_sel[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_2065),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_sel[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_in_in_rt_wt_sel_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_2064),
    .QN(u_NV_NVDLA_cmac_u_core_in_wt_sel[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_990),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_984),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_983),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1268),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_981),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_980),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1278),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1279),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_979),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1280),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_989),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_982),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1012),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1009),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_986),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1244),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1248),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1254),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_985),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1010),
    .QN(mac2accu_data0[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_975),
    .QN(mac2accu_data0[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_974),
    .QN(mac2accu_data0[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_973),
    .QN(mac2accu_data0[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_972),
    .QN(mac2accu_data0[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_971),
    .QN(mac2accu_data0[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_970),
    .QN(mac2accu_data0[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_969),
    .QN(mac2accu_data0[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_968),
    .QN(mac2accu_data0[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_967),
    .QN(mac2accu_data0[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_917),
    .QN(mac2accu_data0[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_905),
    .QN(mac2accu_data0[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_909),
    .QN(mac2accu_data0[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_913),
    .QN(mac2accu_data0[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_919),
    .QN(mac2accu_data0[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_923),
    .QN(mac2accu_data0[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_978),
    .QN(mac2accu_data0[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_977),
    .QN(mac2accu_data0[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data0_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_976),
    .QN(mac2accu_data0[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_966),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_959),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1090),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1057),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_993),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_957),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_956),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_955),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_997),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_994),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_965),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_964),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_963),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_962),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_988),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_961),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1155),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_960),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1143),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_999),
    .QN(mac2accu_data1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_951),
    .QN(mac2accu_data1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1003),
    .QN(mac2accu_data1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1004),
    .QN(mac2accu_data1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_950),
    .QN(mac2accu_data1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_991),
    .QN(mac2accu_data1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1005),
    .QN(mac2accu_data1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_987),
    .QN(mac2accu_data1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1006),
    .QN(mac2accu_data1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1007),
    .QN(mac2accu_data1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_954),
    .QN(mac2accu_data1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_998),
    .QN(mac2accu_data1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_996),
    .QN(mac2accu_data1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_953),
    .QN(mac2accu_data1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_958),
    .QN(mac2accu_data1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1002),
    .QN(mac2accu_data1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_952),
    .QN(mac2accu_data1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1000),
    .QN(mac2accu_data1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data1_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1001),
    .QN(mac2accu_data1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_949),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_944),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_943),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1033),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_942),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1041),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_941),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1055),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1062),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_940),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_948),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1011),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_947),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1008),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_946),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1283),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_945),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_995),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1025),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_939),
    .QN(mac2accu_data2[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_931),
    .QN(mac2accu_data2[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1134),
    .QN(mac2accu_data2[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_930),
    .QN(mac2accu_data2[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_929),
    .QN(mac2accu_data2[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_928),
    .QN(mac2accu_data2[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_927),
    .QN(mac2accu_data2[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_926),
    .QN(mac2accu_data2[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_925),
    .QN(mac2accu_data2[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_924),
    .QN(mac2accu_data2[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_938),
    .QN(mac2accu_data2[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_937),
    .QN(mac2accu_data2[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_936),
    .QN(mac2accu_data2[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_935),
    .QN(mac2accu_data2[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1103),
    .QN(mac2accu_data2[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_934),
    .QN(mac2accu_data2[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_933),
    .QN(mac2accu_data2[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_932),
    .QN(mac2accu_data2[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data2_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1128),
    .QN(mac2accu_data2[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1198),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_918),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_1255),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_916),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1256),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_1258),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1257),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_915),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_1259),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_914),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1282),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1219),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1225),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_922),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1252),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_921),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1251),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_920),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1253),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d1[9]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1261),
    .QN(mac2accu_data3[0]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[10]  (.CLK(nvdla_core_clk),
    .D(n_1267),
    .QN(mac2accu_data3[10]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[11]  (.CLK(nvdla_core_clk),
    .D(n_908),
    .QN(mac2accu_data3[11]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_1271),
    .QN(mac2accu_data3[12]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_1270),
    .QN(mac2accu_data3[13]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[14]  (.CLK(nvdla_core_clk),
    .D(n_907),
    .QN(mac2accu_data3[14]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[15]  (.CLK(nvdla_core_clk),
    .D(n_1273),
    .QN(mac2accu_data3[15]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_1274),
    .QN(mac2accu_data3[16]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_906),
    .QN(mac2accu_data3[17]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[18]  (.CLK(nvdla_core_clk),
    .D(n_1275),
    .QN(mac2accu_data3[18]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1260),
    .QN(mac2accu_data3[1]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_912),
    .QN(mac2accu_data3[2]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1262),
    .QN(mac2accu_data3[3]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1263),
    .QN(mac2accu_data3[4]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_911),
    .QN(mac2accu_data3[5]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1265),
    .QN(mac2accu_data3[6]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1281),
    .QN(mac2accu_data3[7]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_910),
    .QN(mac2accu_data3[8]));
 DFFHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_data3_d2_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1266),
    .QN(mac2accu_data3[9]));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d1_reg (.CLK(nvdla_core_clk),
    .D(n_2150),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d1),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d2_reg (.CLK(nvdla_core_clk),
    .D(n_2191),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d2),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_done_d3_reg (.CLK(nvdla_core_clk),
    .D(n_2196),
    .QN(u_NV_NVDLA_cmac_dp2reg_done),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_11),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_22),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_19),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_21),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_6),
    .QN(mac2accu_mask[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_14),
    .QN(mac2accu_mask[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_23),
    .QN(mac2accu_mask[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_mask_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_17),
    .QN(mac2accu_mask[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1449),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1469),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1468),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1467),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1466),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1465),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1464),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1463),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1450),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d1[8]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1462),
    .QN(mac2accu_pd[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1461),
    .QN(mac2accu_pd[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1460),
    .QN(mac2accu_pd[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1459),
    .QN(mac2accu_pd[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1458),
    .QN(mac2accu_pd[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1457),
    .QN(mac2accu_pd[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1456),
    .QN(mac2accu_pd[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1455),
    .QN(mac2accu_pd[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pd_d2_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1454),
    .QN(mac2accu_pd[8]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1_reg (.CLK(nvdla_core_clk),
    .D(n_28),
    .QN(u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d1),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_core_u_rt_out_out_rt_pvld_d2_reg (.CLK(nvdla_core_clk),
    .D(n_29),
    .QN(mac2accu_pvld),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2121),
    .QN(cmac_a2csb_resp_pd[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[12]  (.CLK(nvdla_core_clk),
    .D(n_2120),
    .QN(cmac_a2csb_resp_pd[12]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[13]  (.CLK(nvdla_core_clk),
    .D(n_2119),
    .QN(cmac_a2csb_resp_pd[13]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[16]  (.CLK(nvdla_core_clk),
    .D(n_2117),
    .QN(cmac_a2csb_resp_pd[16]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[17]  (.CLK(nvdla_core_clk),
    .D(n_2112),
    .QN(cmac_a2csb_resp_pd[17]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2109),
    .QN(cmac_a2csb_resp_pd[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_pd_reg[33]  (.CLK(nvdla_core_clk),
    .D(n_2037),
    .QN(cmac_a2csb_resp_pd[33]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_cmac_a2csb_resp_valid_reg (.CLK(nvdla_core_clk),
    .D(u_NV_NVDLA_cmac_u_reg_n_1258),
    .QN(cmac_a2csb_resp_valid),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_dp2reg_consumer_reg (.CLK(nvdla_core_clk),
    .D(n_19236),
    .QN(u_NV_NVDLA_cmac_u_reg_dp2reg_consumer),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en_reg (.CLK(nvdla_core_clk),
    .D(n_2105),
    .QN(u_NV_NVDLA_cmac_u_reg_reg2dp_d0_op_en),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en_reg (.CLK(nvdla_core_clk),
    .D(n_2104),
    .QN(u_NV_NVDLA_cmac_u_reg_reg2dp_d1_op_en),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_1298),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_1286),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[1]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[22]  (.CLK(nvdla_core_clk),
    .D(n_1293),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[22]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[2]  (.CLK(nvdla_core_clk),
    .D(n_1292),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[2]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[34]  (.CLK(nvdla_core_clk),
    .D(n_1296),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[34]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[35]  (.CLK(nvdla_core_clk),
    .D(n_1290),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[35]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[3]  (.CLK(nvdla_core_clk),
    .D(n_1287),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[3]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[4]  (.CLK(nvdla_core_clk),
    .D(n_1288),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[4]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[54]  (.CLK(nvdla_core_clk),
    .D(n_1294),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[54]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[55]  (.CLK(nvdla_core_clk),
    .D(n_1289),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[55]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[5]  (.CLK(nvdla_core_clk),
    .D(n_1291),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[5]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[6]  (.CLK(nvdla_core_clk),
    .D(n_1297),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[6]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[7]  (.CLK(nvdla_core_clk),
    .D(n_1285),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[7]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[8]  (.CLK(nvdla_core_clk),
    .D(n_1284),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[8]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_req_pd_reg[9]  (.CLK(nvdla_core_clk),
    .D(n_1295),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pd[9]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_req_pvld_reg (.CLK(nvdla_core_clk),
    .D(n_24),
    .QN(u_NV_NVDLA_cmac_u_reg_req_pvld),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_conv_mode_reg (.CLK(nvdla_core_clk),
    .D(n_2103),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_proc_precision_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2108),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .RESETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_proc_precision_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2107),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d0_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_conv_mode_reg (.CLK(nvdla_core_clk),
    .D(n_2113),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[0]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_proc_precision_reg[0]  (.CLK(nvdla_core_clk),
    .D(n_2114),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[12]),
    .RESETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_SL \u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_proc_precision_reg[1]  (.CLK(nvdla_core_clk),
    .D(n_2111),
    .QN(u_NV_NVDLA_cmac_u_reg_u_dual_reg_d1_nvdla_cmac_a_d_misc_cfg_0_out[13]),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_NV_NVDLA_cmac_u_reg_u_single_reg_producer_reg (.CLK(nvdla_core_clk),
    .D(n_2099),
    .QN(u_NV_NVDLA_cmac_u_reg_reg2dp_producer),
    .RESETN(one_),
    .SETN(u_NV_NVDLA_cmac_u_reg_n_1228_BAR));
 DFFASRHQNx1_ASAP7_75t_SL u_partition_m_reset_sync_reset_synced_rstn_NV_GENERIC_CELL_d0_reg (.CLK(nvdla_core_clk),
    .D(n_2123),
    .QN(u_partition_m_reset_sync_reset_synced_rstn_NV_GENERIC_CELL_d0),
    .RESETN(one_),
    .SETN(n_2130));
 DFFASRHQNx1_ASAP7_75t_SL u_partition_m_reset_sync_reset_synced_rstn_NV_GENERIC_CELL_q_reg (.CLK(nvdla_core_clk),
    .D(n_2131),
    .QN(u_partition_m_reset_sync_reset_synced_rstn_reset_),
    .RESETN(one_),
    .SETN(n_2130));
endmodule
