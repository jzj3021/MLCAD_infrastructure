module ac97_top (ac97_reset_pad_o_,
    bit_clk_pad_i,
    clk_i,
    int_o,
    rst_i,
    sdata_pad_i,
    sdata_pad_o,
    suspended_o,
    sync_pad_o,
    wb_ack_o,
    wb_cyc_i,
    wb_stb_i,
    wb_we_i,
    wb_err_o,
    dma_ack_i,
    dma_req_o,
    wb_addr_i,
    wb_data_i,
    wb_data_o,
    wb_sel_i);
 output ac97_reset_pad_o_;
 input bit_clk_pad_i;
 input clk_i;
 output int_o;
 input rst_i;
 input sdata_pad_i;
 output sdata_pad_o;
 output suspended_o;
 output sync_pad_o;
 output wb_ack_o;
 input wb_cyc_i;
 input wb_stb_i;
 input wb_we_i;
 output wb_err_o;
 input [8:0] dma_ack_i;
 output [8:0] dma_req_o;
 input [31:0] wb_addr_i;
 input [31:0] wb_data_i;
 output [31:0] wb_data_o;
 input [3:0] wb_sel_i;

 wire ac97_rst_force;
 wire crac_rd_done;
 wire crac_wr;
 wire i3_empty;
 wire i3_full;
 wire i3_re;
 wire i4_empty;
 wire i4_full;
 wire i4_re;
 wire i6_empty;
 wire i6_full;
 wire i6_re;
 wire ld;
 wire n_0;
 wire n_1;
 wire n_10000;
 wire n_10001;
 wire n_10005;
 wire n_10007;
 wire n_10009;
 wire n_10013;
 wire n_10014;
 wire n_10017;
 wire n_10018;
 wire n_10019;
 wire n_10022;
 wire n_10025;
 wire n_10026;
 wire n_10030;
 wire n_10034;
 wire n_10036;
 wire n_10038;
 wire n_10042;
 wire n_10043;
 wire n_10046;
 wire n_10047;
 wire n_10048;
 wire n_10050;
 wire n_10054;
 wire n_10057;
 wire n_10058;
 wire n_10061;
 wire n_10065;
 wire n_10069;
 wire n_10071;
 wire n_10072;
 wire n_10075;
 wire n_10076;
 wire n_10079;
 wire n_10083;
 wire n_10089;
 wire n_10092;
 wire n_10094;
 wire n_10099;
 wire n_101;
 wire n_10100;
 wire n_10103;
 wire n_10104;
 wire n_10105;
 wire n_10107;
 wire n_10112;
 wire n_10119;
 wire n_10122;
 wire n_10124;
 wire n_10128;
 wire n_10129;
 wire n_10132;
 wire n_10133;
 wire n_10134;
 wire n_10138;
 wire n_10140;
 wire n_10143;
 wire n_10146;
 wire n_10151;
 wire n_10156;
 wire n_10157;
 wire n_10160;
 wire n_10161;
 wire n_10162;
 wire n_10165;
 wire n_10168;
 wire n_1017;
 wire n_10171;
 wire n_10175;
 wire n_10177;
 wire n_10182;
 wire n_10183;
 wire n_10186;
 wire n_10187;
 wire n_10188;
 wire n_10192;
 wire n_10194;
 wire n_10195;
 wire n_10196;
 wire n_10198;
 wire n_10202;
 wire n_10203;
 wire n_10204;
 wire n_10209;
 wire n_10210;
 wire n_10213;
 wire n_10214;
 wire n_10215;
 wire n_10218;
 wire n_10227;
 wire n_10230;
 wire n_10231;
 wire n_10234;
 wire n_10238;
 wire n_10240;
 wire n_10241;
 wire n_10242;
 wire n_10244;
 wire n_10247;
 wire n_10254;
 wire n_10257;
 wire n_10259;
 wire n_10260;
 wire n_10265;
 wire n_10267;
 wire n_10268;
 wire n_10269;
 wire n_10272;
 wire n_10276;
 wire n_10288;
 wire n_1029;
 wire n_10292;
 wire n_103;
 wire n_10302;
 wire n_10303;
 wire n_10306;
 wire n_10310;
 wire n_10315;
 wire n_10317;
 wire n_1032;
 wire n_10321;
 wire n_10323;
 wire n_10324;
 wire n_10326;
 wire n_10327;
 wire n_10329;
 wire n_1033;
 wire n_10330;
 wire n_10335;
 wire n_10336;
 wire n_10339;
 wire n_10344;
 wire n_10346;
 wire n_10350;
 wire n_10351;
 wire n_10352;
 wire n_10356;
 wire n_10363;
 wire n_10366;
 wire n_10369;
 wire n_10370;
 wire n_10372;
 wire n_10376;
 wire n_10377;
 wire n_10378;
 wire n_10379;
 wire n_104;
 wire n_1040;
 wire n_10408;
 wire n_1041;
 wire n_10413;
 wire n_10414;
 wire n_1042;
 wire n_10420;
 wire n_10422;
 wire n_10426;
 wire n_10429;
 wire n_10430;
 wire n_10431;
 wire n_10434;
 wire n_10439;
 wire n_1044;
 wire n_10442;
 wire n_10446;
 wire n_10452;
 wire n_10455;
 wire n_10456;
 wire n_10457;
 wire n_10460;
 wire n_10464;
 wire n_10467;
 wire n_10470;
 wire n_10471;
 wire n_10473;
 wire n_10477;
 wire n_10481;
 wire n_10482;
 wire n_10483;
 wire n_10486;
 wire n_10490;
 wire n_10493;
 wire n_10496;
 wire n_10497;
 wire n_10499;
 wire n_105;
 wire n_10503;
 wire n_10506;
 wire n_10507;
 wire n_10509;
 wire n_1051;
 wire n_1054;
 wire n_10563;
 wire n_10565;
 wire n_10576;
 wire n_1058;
 wire n_1059;
 wire n_106;
 wire n_10613;
 wire n_10614;
 wire n_10615;
 wire n_10617;
 wire n_10620;
 wire n_10621;
 wire n_10622;
 wire n_10623;
 wire n_10624;
 wire n_10626;
 wire n_10627;
 wire n_10628;
 wire n_10629;
 wire n_10631;
 wire n_10633;
 wire n_10635;
 wire n_10636;
 wire n_10637;
 wire n_10638;
 wire n_10640;
 wire n_10641;
 wire n_10642;
 wire n_10644;
 wire n_10649;
 wire n_10651;
 wire n_10654;
 wire n_10656;
 wire n_10657;
 wire n_10659;
 wire n_10660;
 wire n_10661;
 wire n_10665;
 wire n_10666;
 wire n_10669;
 wire n_10670;
 wire n_10676;
 wire n_10679;
 wire n_10680;
 wire n_10681;
 wire n_10683;
 wire n_10684;
 wire n_107;
 wire n_10709;
 wire n_10735;
 wire n_10761;
 wire n_10787;
 wire n_108;
 wire n_10813;
 wire n_1082;
 wire n_1083;
 wire n_10839;
 wire n_1084;
 wire n_1086;
 wire n_10867;
 wire n_10869;
 wire n_10870;
 wire n_10871;
 wire n_10873;
 wire n_10877;
 wire n_10878;
 wire n_1088;
 wire n_10881;
 wire n_10882;
 wire n_10884;
 wire n_10885;
 wire n_10887;
 wire n_10888;
 wire n_10889;
 wire n_1089;
 wire n_10890;
 wire n_10891;
 wire n_10892;
 wire n_10894;
 wire n_10895;
 wire n_10896;
 wire n_10902;
 wire n_10906;
 wire n_10910;
 wire n_10916;
 wire n_10918;
 wire n_10919;
 wire n_10921;
 wire n_10922;
 wire n_10923;
 wire n_10924;
 wire n_10929;
 wire n_10935;
 wire n_10936;
 wire n_10937;
 wire n_10941;
 wire n_10942;
 wire n_10943;
 wire n_10944;
 wire n_10959;
 wire n_10960;
 wire n_10961;
 wire n_10962;
 wire n_10963;
 wire n_10969;
 wire n_10970;
 wire n_10971;
 wire n_11000;
 wire n_11003;
 wire n_11004;
 wire n_11006;
 wire n_11007;
 wire n_11008;
 wire n_11009;
 wire n_11010;
 wire n_11011;
 wire n_11012;
 wire n_11013;
 wire n_11015;
 wire n_11017;
 wire n_11019;
 wire n_11046;
 wire n_111;
 wire n_11124;
 wire n_11125;
 wire n_11126;
 wire n_11127;
 wire n_11128;
 wire n_11129;
 wire n_1113;
 wire n_11130;
 wire n_11131;
 wire n_11132;
 wire n_11133;
 wire n_11134;
 wire n_11135;
 wire n_11136;
 wire n_11137;
 wire n_11138;
 wire n_11139;
 wire n_11140;
 wire n_11141;
 wire n_11142;
 wire n_11143;
 wire n_11144;
 wire n_11183;
 wire n_11184;
 wire n_11185;
 wire n_11186;
 wire n_11187;
 wire n_11188;
 wire n_11190;
 wire n_11191;
 wire n_11197;
 wire n_112;
 wire n_11204;
 wire n_11212;
 wire n_11259;
 wire n_11295;
 wire n_113;
 wire n_11312;
 wire n_1145;
 wire n_11477;
 wire n_11478;
 wire n_11512;
 wire n_11513;
 wire n_1153;
 wire n_11548;
 wire n_11550;
 wire n_11551;
 wire n_11552;
 wire n_11553;
 wire n_11554;
 wire n_11555;
 wire n_11556;
 wire n_11557;
 wire n_11558;
 wire n_11559;
 wire n_11560;
 wire n_11561;
 wire n_11562;
 wire n_11563;
 wire n_11564;
 wire n_11565;
 wire n_11566;
 wire n_11567;
 wire n_11568;
 wire n_11569;
 wire n_11570;
 wire n_11571;
 wire n_11572;
 wire n_11573;
 wire n_11574;
 wire n_11575;
 wire n_11576;
 wire n_11577;
 wire n_11578;
 wire n_11579;
 wire n_11580;
 wire n_11583;
 wire n_11584;
 wire n_11585;
 wire n_11586;
 wire n_11587;
 wire n_11588;
 wire n_11589;
 wire n_11590;
 wire n_11591;
 wire n_11592;
 wire n_11593;
 wire n_11594;
 wire n_11595;
 wire n_11596;
 wire n_11597;
 wire n_11598;
 wire n_11599;
 wire n_116;
 wire n_11600;
 wire n_11601;
 wire n_11602;
 wire n_11603;
 wire n_11604;
 wire n_11605;
 wire n_11606;
 wire n_11607;
 wire n_11608;
 wire n_11609;
 wire n_11610;
 wire n_11611;
 wire n_11612;
 wire n_11613;
 wire n_11614;
 wire n_11615;
 wire n_11618;
 wire n_11619;
 wire n_11620;
 wire n_11621;
 wire n_11622;
 wire n_11623;
 wire n_11624;
 wire n_11625;
 wire n_11626;
 wire n_11627;
 wire n_11628;
 wire n_11629;
 wire n_11630;
 wire n_11631;
 wire n_11632;
 wire n_11633;
 wire n_11634;
 wire n_11635;
 wire n_11636;
 wire n_11637;
 wire n_11638;
 wire n_11639;
 wire n_11640;
 wire n_11641;
 wire n_11642;
 wire n_11643;
 wire n_11644;
 wire n_11645;
 wire n_11646;
 wire n_11647;
 wire n_11648;
 wire n_11649;
 wire n_11650;
 wire n_1167;
 wire n_11693;
 wire n_11697;
 wire n_11699;
 wire n_117;
 wire n_1171;
 wire n_1175;
 wire n_1177;
 wire n_118;
 wire n_1186;
 wire n_11874;
 wire n_119;
 wire n_1192;
 wire n_1193;
 wire n_1194;
 wire n_12;
 wire n_1201;
 wire n_12053;
 wire n_12061;
 wire n_12062;
 wire n_12066;
 wire n_12067;
 wire n_12070;
 wire n_1208;
 wire n_1209;
 wire n_12097;
 wire n_12098;
 wire n_12099;
 wire n_12100;
 wire n_12106;
 wire n_12116;
 wire n_12117;
 wire n_12119;
 wire n_1214;
 wire n_12142;
 wire n_12143;
 wire n_12219;
 wire n_12225;
 wire n_12226;
 wire n_12227;
 wire n_12275;
 wire n_1228;
 wire n_1229;
 wire n_123;
 wire n_1231;
 wire n_12403;
 wire n_12404;
 wire n_12405;
 wire n_12406;
 wire n_12407;
 wire n_12408;
 wire n_12409;
 wire n_1241;
 wire n_12410;
 wire n_12411;
 wire n_12412;
 wire n_12413;
 wire n_12414;
 wire n_12415;
 wire n_12417;
 wire n_12418;
 wire n_12419;
 wire n_12420;
 wire n_12421;
 wire n_12422;
 wire n_12423;
 wire n_12424;
 wire n_12425;
 wire n_12427;
 wire n_12428;
 wire n_12429;
 wire n_12431;
 wire n_12432;
 wire n_12433;
 wire n_12434;
 wire n_12435;
 wire n_12438;
 wire n_1244;
 wire n_12440;
 wire n_12441;
 wire n_12442;
 wire n_12444;
 wire n_12445;
 wire n_12447;
 wire n_12448;
 wire n_12450;
 wire n_12452;
 wire n_12453;
 wire n_12454;
 wire n_12455;
 wire n_12456;
 wire n_12457;
 wire n_12458;
 wire n_12459;
 wire n_12461;
 wire n_12463;
 wire n_12466;
 wire n_12468;
 wire n_12469;
 wire n_12470;
 wire n_12482;
 wire n_12519;
 wire n_1259;
 wire n_1261;
 wire n_128;
 wire n_12837;
 wire n_12838;
 wire n_12839;
 wire n_1284;
 wire n_12842;
 wire n_12843;
 wire n_12845;
 wire n_12846;
 wire n_12847;
 wire n_12848;
 wire n_12849;
 wire n_1285;
 wire n_12851;
 wire n_12854;
 wire n_12855;
 wire n_12856;
 wire n_12857;
 wire n_12858;
 wire n_12859;
 wire n_1286;
 wire n_12861;
 wire n_12863;
 wire n_12865;
 wire n_12867;
 wire n_12868;
 wire n_12869;
 wire n_1287;
 wire n_12870;
 wire n_12871;
 wire n_12872;
 wire n_12873;
 wire n_12874;
 wire n_12875;
 wire n_12876;
 wire n_12877;
 wire n_12878;
 wire n_12879;
 wire n_1288;
 wire n_12880;
 wire n_12881;
 wire n_12882;
 wire n_12883;
 wire n_12884;
 wire n_12885;
 wire n_12886;
 wire n_12887;
 wire n_12888;
 wire n_12889;
 wire n_1289;
 wire n_12890;
 wire n_12891;
 wire n_12892;
 wire n_12893;
 wire n_12895;
 wire n_12896;
 wire n_12897;
 wire n_12898;
 wire n_12899;
 wire n_1290;
 wire n_12900;
 wire n_12901;
 wire n_12902;
 wire n_12908;
 wire n_1292;
 wire n_1296;
 wire n_1297;
 wire n_130;
 wire n_13027;
 wire n_13035;
 wire n_1306;
 wire n_13063;
 wire n_13064;
 wire n_13065;
 wire n_13066;
 wire n_13067;
 wire n_13068;
 wire n_13069;
 wire n_13070;
 wire n_13071;
 wire n_13072;
 wire n_13075;
 wire n_13076;
 wire n_13077;
 wire n_13079;
 wire n_13080;
 wire n_13081;
 wire n_13082;
 wire n_13083;
 wire n_13084;
 wire n_13085;
 wire n_13086;
 wire n_13087;
 wire n_13088;
 wire n_13089;
 wire n_13090;
 wire n_13092;
 wire n_13093;
 wire n_13094;
 wire n_13095;
 wire n_131;
 wire n_1310;
 wire n_13176;
 wire n_1319;
 wire n_132;
 wire n_1322;
 wire n_13236;
 wire n_13237;
 wire n_13244;
 wire n_13246;
 wire n_13247;
 wire n_13249;
 wire n_1325;
 wire n_13266;
 wire n_13269;
 wire n_1329;
 wire n_13295;
 wire n_133;
 wire n_1330;
 wire n_13304;
 wire n_13312;
 wire n_13325;
 wire n_13333;
 wire n_13347;
 wire n_1336;
 wire n_1337;
 wire n_1338;
 wire n_134;
 wire n_13405;
 wire n_13413;
 wire n_13420;
 wire n_1343;
 wire n_1346;
 wire n_13500;
 wire n_13508;
 wire n_13546;
 wire n_13547;
 wire n_13557;
 wire n_1358;
 wire n_13594;
 wire n_13595;
 wire n_13597;
 wire n_13598;
 wire n_13599;
 wire n_136;
 wire n_1361;
 wire n_1362;
 wire n_1365;
 wire n_137;
 wire n_1372;
 wire n_13734;
 wire n_13736;
 wire n_13737;
 wire n_13738;
 wire n_13742;
 wire n_13749;
 wire n_13751;
 wire n_13755;
 wire n_13758;
 wire n_1376;
 wire n_13761;
 wire n_13764;
 wire n_13777;
 wire n_13787;
 wire n_1379;
 wire n_13792;
 wire n_13794;
 wire n_13796;
 wire n_1381;
 wire n_13820;
 wire n_13821;
 wire n_13822;
 wire n_13824;
 wire n_13825;
 wire n_13827;
 wire n_13829;
 wire n_13855;
 wire n_13857;
 wire n_1386;
 wire n_1387;
 wire n_1389;
 wire n_13898;
 wire n_13899;
 wire n_139;
 wire n_1390;
 wire n_1391;
 wire n_13955;
 wire n_13968;
 wire n_13974;
 wire n_13976;
 wire n_13978;
 wire n_13980;
 wire n_13982;
 wire n_13983;
 wire n_13988;
 wire n_13989;
 wire n_13990;
 wire n_13995;
 wire n_13999;
 wire n_14;
 wire n_140;
 wire n_1400;
 wire n_14001;
 wire n_14003;
 wire n_14004;
 wire n_14006;
 wire n_14008;
 wire n_14009;
 wire n_1401;
 wire n_14010;
 wire n_14012;
 wire n_14013;
 wire n_14017;
 wire n_1403;
 wire n_14030;
 wire n_14054;
 wire n_1406;
 wire n_14098;
 wire n_14099;
 wire n_14108;
 wire n_1411;
 wire n_1418;
 wire n_1420;
 wire n_1421;
 wire n_1422;
 wire n_14226;
 wire n_14227;
 wire n_1426;
 wire n_14280;
 wire n_14288;
 wire n_14292;
 wire n_143;
 wire n_1430;
 wire n_14301;
 wire n_14309;
 wire n_14313;
 wire n_14319;
 wire n_1432;
 wire n_14324;
 wire n_14325;
 wire n_14326;
 wire n_14328;
 wire n_1433;
 wire n_14333;
 wire n_1434;
 wire n_14343;
 wire n_14345;
 wire n_1435;
 wire n_14350;
 wire n_1436;
 wire n_1437;
 wire n_14385;
 wire n_14386;
 wire n_1439;
 wire n_14390;
 wire n_14391;
 wire n_14392;
 wire n_14393;
 wire n_14394;
 wire n_14395;
 wire n_14396;
 wire n_14398;
 wire n_14399;
 wire n_144;
 wire n_1440;
 wire n_14400;
 wire n_14401;
 wire n_14402;
 wire n_14403;
 wire n_14405;
 wire n_14418;
 wire n_14424;
 wire n_14425;
 wire n_14431;
 wire n_14432;
 wire n_1444;
 wire n_14448;
 wire n_1452;
 wire n_14546;
 wire n_1455;
 wire n_1456;
 wire n_1457;
 wire n_14570;
 wire n_1459;
 wire n_146;
 wire n_1460;
 wire n_1461;
 wire n_14680;
 wire n_147;
 wire n_1470;
 wire n_1475;
 wire n_14763;
 wire n_14765;
 wire n_14788;
 wire n_14789;
 wire n_14791;
 wire n_14792;
 wire n_14794;
 wire n_148;
 wire n_14816;
 wire n_14820;
 wire n_14821;
 wire n_14825;
 wire n_1483;
 wire n_1484;
 wire n_14859;
 wire n_14864;
 wire n_1488;
 wire n_149;
 wire n_1490;
 wire n_14902;
 wire n_14904;
 wire n_14906;
 wire n_14907;
 wire n_14908;
 wire n_14909;
 wire n_14912;
 wire n_14913;
 wire n_14914;
 wire n_14917;
 wire n_14918;
 wire n_14924;
 wire n_14925;
 wire n_14926;
 wire n_14933;
 wire n_14935;
 wire n_1494;
 wire n_14944;
 wire n_14945;
 wire n_14947;
 wire n_14959;
 wire n_1496;
 wire n_14961;
 wire n_14963;
 wire n_14966;
 wire n_14969;
 wire n_14976;
 wire n_14982;
 wire n_14983;
 wire n_14985;
 wire n_15;
 wire n_15005;
 wire n_15007;
 wire n_1501;
 wire n_15020;
 wire n_15023;
 wire n_15024;
 wire n_15025;
 wire n_15026;
 wire n_1503;
 wire n_15031;
 wire n_15032;
 wire n_15034;
 wire n_15037;
 wire n_15040;
 wire n_15054;
 wire n_15056;
 wire n_15079;
 wire n_15080;
 wire n_15082;
 wire n_15084;
 wire n_15085;
 wire n_15087;
 wire n_15090;
 wire n_15092;
 wire n_15093;
 wire n_15094;
 wire n_1510;
 wire n_15100;
 wire n_15101;
 wire n_15134;
 wire n_15135;
 wire n_15136;
 wire n_15137;
 wire n_15138;
 wire n_15139;
 wire n_15141;
 wire n_15143;
 wire n_15145;
 wire n_1516;
 wire n_15166;
 wire n_1519;
 wire n_152;
 wire n_1523;
 wire n_15269;
 wire n_1527;
 wire n_15271;
 wire n_15272;
 wire n_15274;
 wire n_1528;
 wire n_153;
 wire n_1530;
 wire n_15300;
 wire n_1531;
 wire n_1534;
 wire n_1535;
 wire n_154;
 wire n_1540;
 wire n_15426;
 wire n_1544;
 wire n_1545;
 wire n_1546;
 wire n_15469;
 wire n_1547;
 wire n_15473;
 wire n_15475;
 wire n_1548;
 wire n_15481;
 wire n_15483;
 wire n_15487;
 wire n_1549;
 wire n_15491;
 wire n_15495;
 wire n_15496;
 wire n_155;
 wire n_1550;
 wire n_15506;
 wire n_1551;
 wire n_15515;
 wire n_1552;
 wire n_15521;
 wire n_1553;
 wire n_15534;
 wire n_1554;
 wire n_1555;
 wire n_1558;
 wire n_1559;
 wire n_156;
 wire n_1560;
 wire n_1561;
 wire n_1563;
 wire n_1564;
 wire n_1565;
 wire n_1566;
 wire n_1567;
 wire n_1568;
 wire n_1569;
 wire n_15693;
 wire n_15694;
 wire n_157;
 wire n_1570;
 wire n_1571;
 wire n_1572;
 wire n_1573;
 wire n_1574;
 wire n_1575;
 wire n_1576;
 wire n_1577;
 wire n_15771;
 wire n_15773;
 wire n_15775;
 wire n_1578;
 wire n_1579;
 wire n_158;
 wire n_1580;
 wire n_1581;
 wire n_1582;
 wire n_1583;
 wire n_1584;
 wire n_1585;
 wire n_15854;
 wire n_1586;
 wire n_15867;
 wire n_15869;
 wire n_1587;
 wire n_1588;
 wire n_1589;
 wire n_1590;
 wire n_1591;
 wire n_15915;
 wire n_1592;
 wire n_15920;
 wire n_15923;
 wire n_15927;
 wire n_1593;
 wire n_15931;
 wire n_1594;
 wire n_1595;
 wire n_15952;
 wire n_15954;
 wire n_1596;
 wire n_1597;
 wire n_1598;
 wire n_1599;
 wire n_16;
 wire n_160;
 wire n_1600;
 wire n_16009;
 wire n_1601;
 wire n_1602;
 wire n_1603;
 wire n_16031;
 wire n_1604;
 wire n_1605;
 wire n_1606;
 wire n_1607;
 wire n_1608;
 wire n_1609;
 wire n_161;
 wire n_1610;
 wire n_1611;
 wire n_1612;
 wire n_1613;
 wire n_1614;
 wire n_1615;
 wire n_1616;
 wire n_1617;
 wire n_1618;
 wire n_1619;
 wire n_162;
 wire n_1620;
 wire n_1621;
 wire n_1622;
 wire n_1623;
 wire n_1624;
 wire n_1625;
 wire n_1626;
 wire n_1627;
 wire n_1628;
 wire n_1629;
 wire n_1630;
 wire n_16304;
 wire n_1631;
 wire n_16314;
 wire n_1632;
 wire n_1633;
 wire n_1634;
 wire n_1635;
 wire n_1637;
 wire n_16416;
 wire n_16427;
 wire n_1643;
 wire n_16436;
 wire n_16439;
 wire n_1645;
 wire n_16458;
 wire n_1646;
 wire n_1647;
 wire n_1648;
 wire n_1649;
 wire n_1651;
 wire n_16593;
 wire n_166;
 wire n_1660;
 wire n_1661;
 wire n_1666;
 wire n_16664;
 wire n_1667;
 wire n_16671;
 wire n_16672;
 wire n_16680;
 wire n_16684;
 wire n_16720;
 wire n_16721;
 wire n_16722;
 wire n_16723;
 wire n_16724;
 wire n_16725;
 wire n_16726;
 wire n_16727;
 wire n_16728;
 wire n_16730;
 wire n_16731;
 wire n_16732;
 wire n_16733;
 wire n_16736;
 wire n_16737;
 wire n_16738;
 wire n_16739;
 wire n_16741;
 wire n_16742;
 wire n_16743;
 wire n_16749;
 wire n_16750;
 wire n_16751;
 wire n_1677;
 wire n_1678;
 wire n_16781;
 wire n_16788;
 wire n_1679;
 wire n_16797;
 wire n_16798;
 wire n_1680;
 wire n_16805;
 wire n_16807;
 wire n_1681;
 wire n_16816;
 wire n_16819;
 wire n_16828;
 wire n_16853;
 wire n_16857;
 wire n_16858;
 wire n_16880;
 wire n_16895;
 wire n_16899;
 wire n_169;
 wire n_16900;
 wire n_16908;
 wire n_1692;
 wire n_1699;
 wire n_1701;
 wire n_1704;
 wire n_1705;
 wire n_1707;
 wire n_17079;
 wire n_171;
 wire n_17108;
 wire n_17110;
 wire n_1714;
 wire n_17184;
 wire n_172;
 wire n_1723;
 wire n_17252;
 wire n_17254;
 wire n_17304;
 wire n_1734;
 wire n_1736;
 wire n_17388;
 wire n_1739;
 wire n_17399;
 wire n_17400;
 wire n_17401;
 wire n_17402;
 wire n_17403;
 wire n_1742;
 wire n_1744;
 wire n_17440;
 wire n_17441;
 wire n_1745;
 wire n_1747;
 wire n_17489;
 wire n_1749;
 wire n_17490;
 wire n_17492;
 wire n_1751;
 wire n_17513;
 wire n_1752;
 wire n_17525;
 wire n_17528;
 wire n_1753;
 wire n_17530;
 wire n_17532;
 wire n_17534;
 wire n_1754;
 wire n_17542;
 wire n_17545;
 wire n_1755;
 wire n_17563;
 wire n_17565;
 wire n_17567;
 wire n_17569;
 wire n_1757;
 wire n_17573;
 wire n_17575;
 wire n_17577;
 wire n_17578;
 wire n_17579;
 wire n_17583;
 wire n_17584;
 wire n_17591;
 wire n_17594;
 wire n_17595;
 wire n_17596;
 wire n_17597;
 wire n_17599;
 wire n_176;
 wire n_1760;
 wire n_17600;
 wire n_17606;
 wire n_17608;
 wire n_17609;
 wire n_17613;
 wire n_17614;
 wire n_17615;
 wire n_17616;
 wire n_17617;
 wire n_17618;
 wire n_1762;
 wire n_17623;
 wire n_17624;
 wire n_17625;
 wire n_17626;
 wire n_1764;
 wire n_1765;
 wire n_1766;
 wire n_1767;
 wire n_17672;
 wire n_1768;
 wire n_17686;
 wire n_17687;
 wire n_17688;
 wire n_1769;
 wire n_17690;
 wire n_1770;
 wire n_17704;
 wire n_17705;
 wire n_17706;
 wire n_17711;
 wire n_17712;
 wire n_1775;
 wire n_1777;
 wire n_17778;
 wire n_17785;
 wire n_17787;
 wire n_1779;
 wire n_178;
 wire n_1780;
 wire n_17801;
 wire n_17809;
 wire n_1781;
 wire n_1782;
 wire n_1783;
 wire n_1784;
 wire n_1785;
 wire n_1788;
 wire n_1789;
 wire n_179;
 wire n_17924;
 wire n_17925;
 wire n_17927;
 wire n_1793;
 wire n_17938;
 wire n_1794;
 wire n_1797;
 wire n_17979;
 wire n_1801;
 wire n_18018;
 wire n_1802;
 wire n_1803;
 wire n_1805;
 wire n_18058;
 wire n_18060;
 wire n_18066;
 wire n_18068;
 wire n_1807;
 wire n_1808;
 wire n_18089;
 wire n_1809;
 wire n_18092;
 wire n_181;
 wire n_1812;
 wire n_1816;
 wire n_18195;
 wire n_1820;
 wire n_1828;
 wire n_18289;
 wire n_183;
 wire n_1831;
 wire n_1836;
 wire n_1838;
 wire n_184;
 wire n_1840;
 wire n_1841;
 wire n_1842;
 wire n_1844;
 wire n_18448;
 wire n_1845;
 wire n_1846;
 wire n_1847;
 wire n_18480;
 wire n_18483;
 wire n_1849;
 wire n_18491;
 wire n_185;
 wire n_1850;
 wire n_1852;
 wire n_18524;
 wire n_1853;
 wire n_1857;
 wire n_18591;
 wire n_186;
 wire n_1861;
 wire n_1863;
 wire n_18652;
 wire n_18653;
 wire n_18654;
 wire n_18655;
 wire n_18658;
 wire n_18660;
 wire n_18666;
 wire n_18667;
 wire n_18668;
 wire n_18679;
 wire n_18683;
 wire n_18684;
 wire n_1869;
 wire n_18704;
 wire n_18706;
 wire n_18707;
 wire n_18709;
 wire n_18710;
 wire n_18711;
 wire n_1872;
 wire n_18739;
 wire n_18742;
 wire n_18743;
 wire n_18745;
 wire n_18841;
 wire n_1885;
 wire n_18857;
 wire n_1887;
 wire n_18871;
 wire n_18872;
 wire n_18873;
 wire n_18875;
 wire n_1888;
 wire n_18885;
 wire n_18886;
 wire n_18887;
 wire n_18888;
 wire n_18889;
 wire n_18894;
 wire n_18895;
 wire n_18896;
 wire n_18897;
 wire n_18899;
 wire n_18900;
 wire n_18902;
 wire n_18903;
 wire n_1892;
 wire n_18928;
 wire n_18931;
 wire n_18933;
 wire n_1894;
 wire n_1895;
 wire n_1896;
 wire n_18964;
 wire n_18966;
 wire n_19;
 wire n_190;
 wire n_19002;
 wire n_19004;
 wire n_19005;
 wire n_19006;
 wire n_19007;
 wire n_19008;
 wire n_19009;
 wire n_19010;
 wire n_19013;
 wire n_1903;
 wire n_1904;
 wire n_19045;
 wire n_19046;
 wire n_19047;
 wire n_19067;
 wire n_19068;
 wire n_19069;
 wire n_1913;
 wire n_19132;
 wire n_19133;
 wire n_1914;
 wire n_1915;
 wire n_1917;
 wire n_1919;
 wire n_1920;
 wire n_19234;
 wire n_19235;
 wire n_19237;
 wire n_19241;
 wire n_1932;
 wire n_19378;
 wire n_19383;
 wire n_19495;
 wire n_19496;
 wire n_19497;
 wire n_195;
 wire n_19501;
 wire n_19502;
 wire n_19503;
 wire n_19504;
 wire n_19505;
 wire n_19506;
 wire n_19509;
 wire n_19510;
 wire n_1955;
 wire n_1957;
 wire n_19576;
 wire n_19577;
 wire n_19578;
 wire n_1959;
 wire n_19593;
 wire n_19594;
 wire n_19615;
 wire n_19616;
 wire n_19617;
 wire n_19619;
 wire n_19620;
 wire n_19621;
 wire n_19622;
 wire n_19623;
 wire n_1965;
 wire n_19669;
 wire n_19672;
 wire n_1968;
 wire n_19687;
 wire n_19688;
 wire n_1972;
 wire n_198;
 wire n_1990;
 wire n_1992;
 wire n_1999;
 wire n_2;
 wire n_20;
 wire n_2002;
 wire n_2009;
 wire n_201;
 wire n_2013;
 wire n_2014;
 wire n_2016;
 wire n_2020;
 wire n_2021;
 wire n_2024;
 wire n_20245;
 wire n_20246;
 wire n_20247;
 wire n_2029;
 wire n_203;
 wire n_2031;
 wire n_20316;
 wire n_20317;
 wire n_20319;
 wire n_2034;
 wire n_2036;
 wire n_2038;
 wire n_20426;
 wire n_2048;
 wire n_2052;
 wire n_2053;
 wire n_2057;
 wire n_2059;
 wire n_20593;
 wire n_20594;
 wire n_20595;
 wire n_20597;
 wire n_206;
 wire n_2063;
 wire n_2065;
 wire n_20669;
 wire n_20671;
 wire n_20673;
 wire n_2073;
 wire n_2074;
 wire n_20756;
 wire n_20759;
 wire n_20760;
 wire n_20783;
 wire n_2079;
 wire n_20821;
 wire n_20824;
 wire n_2092;
 wire n_2095;
 wire n_20972;
 wire n_20973;
 wire n_2098;
 wire n_21;
 wire n_21015;
 wire n_21024;
 wire n_21026;
 wire n_21027;
 wire n_2106;
 wire n_21076;
 wire n_2108;
 wire n_21092;
 wire n_21093;
 wire n_21094;
 wire n_21095;
 wire n_21096;
 wire n_21097;
 wire n_21098;
 wire n_21099;
 wire n_211;
 wire n_21100;
 wire n_21101;
 wire n_21102;
 wire n_21103;
 wire n_21104;
 wire n_21105;
 wire n_21106;
 wire n_21107;
 wire n_21108;
 wire n_21109;
 wire n_21110;
 wire n_21111;
 wire n_21112;
 wire n_21113;
 wire n_21114;
 wire n_21115;
 wire n_21116;
 wire n_21117;
 wire n_21118;
 wire n_21119;
 wire n_21120;
 wire n_21121;
 wire n_21122;
 wire n_21123;
 wire n_21124;
 wire n_2113;
 wire n_21141;
 wire n_21147;
 wire n_21148;
 wire n_2118;
 wire n_2119;
 wire n_21190;
 wire n_212;
 wire n_2120;
 wire n_21225;
 wire n_21226;
 wire n_21231;
 wire n_21234;
 wire n_2124;
 wire n_21261;
 wire n_21263;
 wire n_21264;
 wire n_2129;
 wire n_2130;
 wire n_21311;
 wire n_21312;
 wire n_21317;
 wire n_21320;
 wire n_21321;
 wire n_21324;
 wire n_21325;
 wire n_21328;
 wire n_21331;
 wire n_21332;
 wire n_21335;
 wire n_21341;
 wire n_21342;
 wire n_21343;
 wire n_2136;
 wire n_2138;
 wire n_2143;
 wire n_2149;
 wire n_21507;
 wire n_21513;
 wire n_21514;
 wire n_21515;
 wire n_21516;
 wire n_21517;
 wire n_21518;
 wire n_21520;
 wire n_21521;
 wire n_21527;
 wire n_21530;
 wire n_21532;
 wire n_21534;
 wire n_21536;
 wire n_21538;
 wire n_21539;
 wire n_21540;
 wire n_21541;
 wire n_21543;
 wire n_21546;
 wire n_21549;
 wire n_2155;
 wire n_21550;
 wire n_21552;
 wire n_21553;
 wire n_21554;
 wire n_21599;
 wire n_21600;
 wire n_2162;
 wire n_21631;
 wire n_21638;
 wire n_2164;
 wire n_21646;
 wire n_21665;
 wire n_21669;
 wire n_21673;
 wire n_2168;
 wire n_21695;
 wire n_21696;
 wire n_21697;
 wire n_217;
 wire n_21705;
 wire n_21709;
 wire n_2174;
 wire n_2176;
 wire n_21776;
 wire n_21777;
 wire n_21778;
 wire n_21780;
 wire n_21784;
 wire n_2179;
 wire n_21793;
 wire n_21794;
 wire n_21795;
 wire n_218;
 wire n_2180;
 wire n_2183;
 wire n_2185;
 wire n_21865;
 wire n_21867;
 wire n_21871;
 wire n_21872;
 wire n_21874;
 wire n_21876;
 wire n_21878;
 wire n_2188;
 wire n_219;
 wire n_2190;
 wire n_2191;
 wire n_2193;
 wire n_21938;
 wire n_21947;
 wire n_2195;
 wire n_21996;
 wire n_22;
 wire n_220;
 wire n_22025;
 wire n_22027;
 wire n_22028;
 wire n_22029;
 wire n_2203;
 wire n_2205;
 wire n_22059;
 wire n_2206;
 wire n_22060;
 wire n_22062;
 wire n_22064;
 wire n_2207;
 wire n_2208;
 wire n_2216;
 wire n_22163;
 wire n_2217;
 wire n_22174;
 wire n_22175;
 wire n_22176;
 wire n_22177;
 wire n_22178;
 wire n_22179;
 wire n_22180;
 wire n_22181;
 wire n_22182;
 wire n_22183;
 wire n_22184;
 wire n_22185;
 wire n_22186;
 wire n_22187;
 wire n_22188;
 wire n_22189;
 wire n_22190;
 wire n_2222;
 wire n_2223;
 wire n_2224;
 wire n_22247;
 wire n_22248;
 wire n_22250;
 wire n_22252;
 wire n_22253;
 wire n_22254;
 wire n_22256;
 wire n_22257;
 wire n_2226;
 wire n_22267;
 wire n_22268;
 wire n_22269;
 wire n_2227;
 wire n_22270;
 wire n_22271;
 wire n_22272;
 wire n_22273;
 wire n_22274;
 wire n_22275;
 wire n_22276;
 wire n_22277;
 wire n_22278;
 wire n_22279;
 wire n_2228;
 wire n_22280;
 wire n_22281;
 wire n_22282;
 wire n_22283;
 wire n_223;
 wire n_2230;
 wire n_22311;
 wire n_22315;
 wire n_2232;
 wire n_2234;
 wire n_2235;
 wire n_2236;
 wire n_2237;
 wire n_22371;
 wire n_2238;
 wire n_22396;
 wire n_22407;
 wire n_22413;
 wire n_22415;
 wire n_22424;
 wire n_22430;
 wire n_22432;
 wire n_2247;
 wire n_22482;
 wire n_225;
 wire n_22505;
 wire n_22506;
 wire n_22508;
 wire n_2251;
 wire n_22530;
 wire n_22532;
 wire n_2254;
 wire n_2256;
 wire n_22577;
 wire n_22578;
 wire n_226;
 wire n_2261;
 wire n_22629;
 wire n_2263;
 wire n_22632;
 wire n_22635;
 wire n_22640;
 wire n_22642;
 wire n_2265;
 wire n_2266;
 wire n_2268;
 wire n_22694;
 wire n_227;
 wire n_2271;
 wire n_22715;
 wire n_22718;
 wire n_2273;
 wire n_2274;
 wire n_2275;
 wire n_2277;
 wire n_22774;
 wire n_22775;
 wire n_2278;
 wire n_22780;
 wire n_2281;
 wire n_2282;
 wire n_22827;
 wire n_22828;
 wire n_22829;
 wire n_22835;
 wire n_22837;
 wire n_22839;
 wire n_22841;
 wire n_22842;
 wire n_22844;
 wire n_22845;
 wire n_22846;
 wire n_22851;
 wire n_22852;
 wire n_2286;
 wire n_2288;
 wire n_2289;
 wire n_229;
 wire n_2290;
 wire n_2291;
 wire n_22919;
 wire n_2292;
 wire n_22922;
 wire n_22923;
 wire n_22924;
 wire n_22927;
 wire n_22928;
 wire n_22932;
 wire n_22933;
 wire n_22938;
 wire n_22964;
 wire n_2298;
 wire n_23;
 wire n_230;
 wire n_2302;
 wire n_2304;
 wire n_2306;
 wire n_23079;
 wire n_23099;
 wire n_231;
 wire n_23100;
 wire n_23101;
 wire n_23110;
 wire n_23129;
 wire n_23130;
 wire n_23131;
 wire n_23150;
 wire n_23154;
 wire n_232;
 wire n_23285;
 wire n_23286;
 wire n_23287;
 wire n_23289;
 wire n_23296;
 wire n_2330;
 wire n_2331;
 wire n_2332;
 wire n_2337;
 wire n_23393;
 wire n_23394;
 wire n_234;
 wire n_2345;
 wire n_2348;
 wire n_2350;
 wire n_23504;
 wire n_23508;
 wire n_23524;
 wire n_23526;
 wire n_23529;
 wire n_23530;
 wire n_23531;
 wire n_2362;
 wire n_2363;
 wire n_23655;
 wire n_23656;
 wire n_23659;
 wire n_23660;
 wire n_23661;
 wire n_23671;
 wire n_2369;
 wire n_2371;
 wire n_2373;
 wire n_2375;
 wire n_2384;
 wire n_2385;
 wire n_2393;
 wire n_23971;
 wire n_24;
 wire n_2401;
 wire n_2403;
 wire n_2413;
 wire n_2416;
 wire n_2418;
 wire n_2419;
 wire n_2420;
 wire n_2424;
 wire n_2427;
 wire n_2428;
 wire n_2429;
 wire n_24316;
 wire n_2432;
 wire n_2433;
 wire n_24336;
 wire n_24337;
 wire n_2434;
 wire n_24341;
 wire n_2435;
 wire n_24350;
 wire n_24351;
 wire n_24367;
 wire n_24373;
 wire n_24374;
 wire n_24375;
 wire n_2440;
 wire n_2442;
 wire n_2444;
 wire n_2446;
 wire n_2447;
 wire n_245;
 wire n_24509;
 wire n_24510;
 wire n_24511;
 wire n_24512;
 wire n_24513;
 wire n_24516;
 wire n_2452;
 wire n_24523;
 wire n_24524;
 wire n_2453;
 wire n_24532;
 wire n_24536;
 wire n_2454;
 wire n_24553;
 wire n_2458;
 wire n_24580;
 wire n_24586;
 wire n_24587;
 wire n_24588;
 wire n_24594;
 wire n_24595;
 wire n_24596;
 wire n_2462;
 wire n_24622;
 wire n_24623;
 wire n_24624;
 wire n_24625;
 wire n_24626;
 wire n_24627;
 wire n_24628;
 wire n_24632;
 wire n_24633;
 wire n_24635;
 wire n_24637;
 wire n_2464;
 wire n_24641;
 wire n_2465;
 wire n_2466;
 wire n_24669;
 wire n_2467;
 wire n_24670;
 wire n_24672;
 wire n_2468;
 wire n_247;
 wire n_2470;
 wire n_2471;
 wire n_24725;
 wire n_24726;
 wire n_2473;
 wire n_24730;
 wire n_24732;
 wire n_24733;
 wire n_24734;
 wire n_24735;
 wire n_24736;
 wire n_24737;
 wire n_24738;
 wire n_24739;
 wire n_24741;
 wire n_24742;
 wire n_24745;
 wire n_2475;
 wire n_24750;
 wire n_24753;
 wire n_24759;
 wire n_24761;
 wire n_24762;
 wire n_24763;
 wire n_24764;
 wire n_2477;
 wire n_2478;
 wire n_2479;
 wire n_24801;
 wire n_24803;
 wire n_24804;
 wire n_24805;
 wire n_24806;
 wire n_24807;
 wire n_24808;
 wire n_24809;
 wire n_24810;
 wire n_24811;
 wire n_24812;
 wire n_24813;
 wire n_24814;
 wire n_24815;
 wire n_24816;
 wire n_24817;
 wire n_24818;
 wire n_24819;
 wire n_24820;
 wire n_24821;
 wire n_24822;
 wire n_24823;
 wire n_24824;
 wire n_24825;
 wire n_24826;
 wire n_24827;
 wire n_24828;
 wire n_24829;
 wire n_24830;
 wire n_24831;
 wire n_24832;
 wire n_24833;
 wire n_24835;
 wire n_24837;
 wire n_24838;
 wire n_2486;
 wire n_24883;
 wire n_24886;
 wire n_24888;
 wire n_24889;
 wire n_24890;
 wire n_24891;
 wire n_24892;
 wire n_2490;
 wire n_2491;
 wire n_2492;
 wire n_2496;
 wire n_24975;
 wire n_24978;
 wire n_24979;
 wire n_2498;
 wire n_24980;
 wire n_24981;
 wire n_24982;
 wire n_24984;
 wire n_24985;
 wire n_24986;
 wire n_24987;
 wire n_24988;
 wire n_24989;
 wire n_24990;
 wire n_24991;
 wire n_24992;
 wire n_24993;
 wire n_24995;
 wire n_24997;
 wire n_24998;
 wire n_24999;
 wire n_25;
 wire n_2500;
 wire n_25001;
 wire n_25002;
 wire n_25004;
 wire n_25005;
 wire n_25006;
 wire n_25007;
 wire n_25008;
 wire n_25009;
 wire n_25010;
 wire n_2503;
 wire n_2508;
 wire n_2509;
 wire n_2511;
 wire n_2513;
 wire n_2516;
 wire n_2517;
 wire n_2518;
 wire n_2519;
 wire n_2520;
 wire n_2522;
 wire n_2523;
 wire n_2524;
 wire n_25293;
 wire n_25294;
 wire n_253;
 wire n_25330;
 wire n_25331;
 wire n_25332;
 wire n_25333;
 wire n_25378;
 wire n_25379;
 wire n_25380;
 wire n_25381;
 wire n_25382;
 wire n_25383;
 wire n_25384;
 wire n_25385;
 wire n_25386;
 wire n_25387;
 wire n_25388;
 wire n_25389;
 wire n_2539;
 wire n_25390;
 wire n_25391;
 wire n_25392;
 wire n_25393;
 wire n_25394;
 wire n_25395;
 wire n_25398;
 wire n_2540;
 wire n_25405;
 wire n_2541;
 wire n_25438;
 wire n_25439;
 wire n_2544;
 wire n_25440;
 wire n_2546;
 wire n_25528;
 wire n_25529;
 wire n_25530;
 wire n_2557;
 wire n_256;
 wire n_2560;
 wire n_2564;
 wire n_2565;
 wire n_2566;
 wire n_2567;
 wire n_25673;
 wire n_25674;
 wire n_25675;
 wire n_25677;
 wire n_25678;
 wire n_25679;
 wire n_25680;
 wire n_25681;
 wire n_25682;
 wire n_257;
 wire n_2571;
 wire n_2573;
 wire n_2574;
 wire n_2575;
 wire n_2576;
 wire n_2578;
 wire n_2579;
 wire n_258;
 wire n_2584;
 wire n_259;
 wire n_25928;
 wire n_2594;
 wire n_2595;
 wire n_25953;
 wire n_25954;
 wire n_25955;
 wire n_25956;
 wire n_2596;
 wire n_25961;
 wire n_25964;
 wire n_25965;
 wire n_25967;
 wire n_2598;
 wire n_2603;
 wire n_26050;
 wire n_26054;
 wire n_26055;
 wire n_26057;
 wire n_2608;
 wire n_2609;
 wire n_26098;
 wire n_2610;
 wire n_26103;
 wire n_2611;
 wire n_2612;
 wire n_26182;
 wire n_26183;
 wire n_2619;
 wire n_262;
 wire n_2620;
 wire n_2623;
 wire n_2624;
 wire n_26250;
 wire n_26254;
 wire n_26255;
 wire n_263;
 wire n_26376;
 wire n_26379;
 wire n_26382;
 wire n_26383;
 wire n_26384;
 wire n_26385;
 wire n_26386;
 wire n_26387;
 wire n_26388;
 wire n_26389;
 wire n_2639;
 wire n_26390;
 wire n_26391;
 wire n_26392;
 wire n_26393;
 wire n_26394;
 wire n_26395;
 wire n_26396;
 wire n_26398;
 wire n_26399;
 wire n_264;
 wire n_2640;
 wire n_26400;
 wire n_26401;
 wire n_26402;
 wire n_26403;
 wire n_26404;
 wire n_26405;
 wire n_26406;
 wire n_26407;
 wire n_26408;
 wire n_26409;
 wire n_2641;
 wire n_26410;
 wire n_26411;
 wire n_26412;
 wire n_26413;
 wire n_26414;
 wire n_26415;
 wire n_26416;
 wire n_26417;
 wire n_26418;
 wire n_26419;
 wire n_2642;
 wire n_26427;
 wire n_26428;
 wire n_2643;
 wire n_2644;
 wire n_2645;
 wire n_2646;
 wire n_2647;
 wire n_26497;
 wire n_26498;
 wire n_26499;
 wire n_265;
 wire n_2650;
 wire n_26501;
 wire n_2651;
 wire n_2652;
 wire n_2653;
 wire n_26539;
 wire n_26540;
 wire n_26541;
 wire n_2655;
 wire n_26553;
 wire n_26556;
 wire n_2657;
 wire n_26577;
 wire n_26579;
 wire n_26581;
 wire n_2660;
 wire n_2663;
 wire n_2664;
 wire n_26645;
 wire n_26646;
 wire n_2669;
 wire n_267;
 wire n_26710;
 wire n_26711;
 wire n_26712;
 wire n_26713;
 wire n_26714;
 wire n_26733;
 wire n_2678;
 wire n_26801;
 wire n_26802;
 wire n_26803;
 wire n_26806;
 wire n_26807;
 wire n_26811;
 wire n_26815;
 wire n_26819;
 wire n_26823;
 wire n_26827;
 wire n_2683;
 wire n_26831;
 wire n_2684;
 wire n_2685;
 wire n_26859;
 wire n_2686;
 wire n_2687;
 wire n_2688;
 wire n_2689;
 wire n_269;
 wire n_26904;
 wire n_2691;
 wire n_2692;
 wire n_2693;
 wire n_2694;
 wire n_2695;
 wire n_2696;
 wire n_27003;
 wire n_27004;
 wire n_27013;
 wire n_2702;
 wire n_27038;
 wire n_27057;
 wire n_27058;
 wire n_27059;
 wire n_2706;
 wire n_27060;
 wire n_27061;
 wire n_2708;
 wire n_2712;
 wire n_27128;
 wire n_27129;
 wire n_2713;
 wire n_27131;
 wire n_27132;
 wire n_27133;
 wire n_27134;
 wire n_27135;
 wire n_27136;
 wire n_2715;
 wire n_2716;
 wire n_2719;
 wire n_2721;
 wire n_27219;
 wire n_27223;
 wire n_27224;
 wire n_27225;
 wire n_27227;
 wire n_27234;
 wire n_27235;
 wire n_27236;
 wire n_27237;
 wire n_2724;
 wire n_27257;
 wire n_2727;
 wire n_273;
 wire n_27305;
 wire n_27315;
 wire n_27316;
 wire n_27317;
 wire n_27320;
 wire n_27321;
 wire n_2733;
 wire n_2734;
 wire n_27341;
 wire n_2735;
 wire n_27368;
 wire n_27369;
 wire n_2737;
 wire n_27370;
 wire n_27372;
 wire n_27373;
 wire n_27381;
 wire n_27382;
 wire n_27383;
 wire n_274;
 wire n_2741;
 wire n_2743;
 wire n_2744;
 wire n_2746;
 wire n_2748;
 wire n_275;
 wire n_2752;
 wire n_27521;
 wire n_2753;
 wire n_2767;
 wire n_2773;
 wire n_2775;
 wire n_278;
 wire n_27878;
 wire n_2788;
 wire n_27880;
 wire n_280;
 wire n_281;
 wire n_28102;
 wire n_28103;
 wire n_28110;
 wire n_28111;
 wire n_28121;
 wire n_28122;
 wire n_2817;
 wire n_28235;
 wire n_28239;
 wire n_28240;
 wire n_28246;
 wire n_28251;
 wire n_28276;
 wire n_28294;
 wire n_28316;
 wire n_28327;
 wire n_28330;
 wire n_2836;
 wire n_28364;
 wire n_28367;
 wire n_28368;
 wire n_28370;
 wire n_28371;
 wire n_28381;
 wire n_28391;
 wire n_28412;
 wire n_28413;
 wire n_28424;
 wire n_28441;
 wire n_28443;
 wire n_285;
 wire n_28520;
 wire n_28521;
 wire n_28528;
 wire n_28529;
 wire n_28594;
 wire n_28595;
 wire n_286;
 wire n_28662;
 wire n_28663;
 wire n_28664;
 wire n_28669;
 wire n_28671;
 wire n_28672;
 wire n_28673;
 wire n_28674;
 wire n_28689;
 wire n_28690;
 wire n_28691;
 wire n_28692;
 wire n_28696;
 wire n_28745;
 wire n_28746;
 wire n_28747;
 wire n_28774;
 wire n_28808;
 wire n_28810;
 wire n_28811;
 wire n_28814;
 wire n_28848;
 wire n_28849;
 wire n_28850;
 wire n_28852;
 wire n_28879;
 wire n_28880;
 wire n_28881;
 wire n_28884;
 wire n_28885;
 wire n_28893;
 wire n_28895;
 wire n_289;
 wire n_28901;
 wire n_28913;
 wire n_28926;
 wire n_28948;
 wire n_28950;
 wire n_28951;
 wire n_28952;
 wire n_28953;
 wire n_28954;
 wire n_28955;
 wire n_290;
 wire n_29003;
 wire n_29004;
 wire n_29005;
 wire n_29006;
 wire n_29007;
 wire n_29008;
 wire n_29009;
 wire n_29010;
 wire n_29011;
 wire n_29012;
 wire n_29013;
 wire n_29014;
 wire n_29015;
 wire n_29016;
 wire n_29017;
 wire n_29018;
 wire n_29019;
 wire n_29020;
 wire n_29021;
 wire n_29022;
 wire n_29023;
 wire n_29024;
 wire n_29025;
 wire n_29026;
 wire n_29027;
 wire n_29028;
 wire n_29029;
 wire n_29030;
 wire n_29031;
 wire n_29032;
 wire n_29033;
 wire n_29034;
 wire n_29035;
 wire n_29036;
 wire n_29037;
 wire n_29038;
 wire n_29039;
 wire n_29040;
 wire n_29041;
 wire n_29073;
 wire n_29074;
 wire n_29076;
 wire n_29077;
 wire n_29078;
 wire n_29079;
 wire n_29080;
 wire n_29081;
 wire n_29082;
 wire n_29083;
 wire n_29088;
 wire n_29089;
 wire n_29092;
 wire n_29093;
 wire n_29094;
 wire n_29095;
 wire n_29096;
 wire n_29097;
 wire n_29098;
 wire n_29099;
 wire n_291;
 wire n_29100;
 wire n_29101;
 wire n_29102;
 wire n_29103;
 wire n_29104;
 wire n_29105;
 wire n_29106;
 wire n_29107;
 wire n_293;
 wire n_2931;
 wire n_29310;
 wire n_29312;
 wire n_29313;
 wire n_29314;
 wire n_2932;
 wire n_2933;
 wire n_2934;
 wire n_2935;
 wire n_29352;
 wire n_29355;
 wire n_29356;
 wire n_29358;
 wire n_29361;
 wire n_29362;
 wire n_29364;
 wire n_29365;
 wire n_29366;
 wire n_294;
 wire n_2940;
 wire n_2941;
 wire n_2947;
 wire n_2948;
 wire n_29495;
 wire n_295;
 wire n_2950;
 wire n_2951;
 wire n_2952;
 wire n_29527;
 wire n_29528;
 wire n_29529;
 wire n_2953;
 wire n_29530;
 wire n_29531;
 wire n_29532;
 wire n_29533;
 wire n_29534;
 wire n_29543;
 wire n_29544;
 wire n_29545;
 wire n_29546;
 wire n_29547;
 wire n_29548;
 wire n_29549;
 wire n_2955;
 wire n_29550;
 wire n_29553;
 wire n_29554;
 wire n_29555;
 wire n_29556;
 wire n_29557;
 wire n_29558;
 wire n_2956;
 wire n_2957;
 wire n_29618;
 wire n_29619;
 wire n_29621;
 wire n_29630;
 wire n_2964;
 wire n_2965;
 wire n_29657;
 wire n_29658;
 wire n_29659;
 wire n_29661;
 wire n_29662;
 wire n_2967;
 wire n_29687;
 wire n_29688;
 wire n_2974;
 wire n_2976;
 wire n_2977;
 wire n_29787;
 wire n_29790;
 wire n_2980;
 wire n_2983;
 wire n_2984;
 wire n_2985;
 wire n_29874;
 wire n_29881;
 wire n_29883;
 wire n_29884;
 wire n_29885;
 wire n_29888;
 wire n_29889;
 wire n_29890;
 wire n_29891;
 wire n_29896;
 wire n_29897;
 wire n_29898;
 wire n_29899;
 wire n_2990;
 wire n_29902;
 wire n_29903;
 wire n_29904;
 wire n_29905;
 wire n_29906;
 wire n_29907;
 wire n_29908;
 wire n_29909;
 wire n_29910;
 wire n_29911;
 wire n_29914;
 wire n_29915;
 wire n_29934;
 wire n_29938;
 wire n_29939;
 wire n_29940;
 wire n_29948;
 wire n_29949;
 wire n_29953;
 wire n_29970;
 wire n_3;
 wire n_30059;
 wire n_30060;
 wire n_30061;
 wire n_30062;
 wire n_30078;
 wire n_301;
 wire n_30235;
 wire n_30247;
 wire n_30253;
 wire n_30254;
 wire n_303;
 wire n_30330;
 wire n_30331;
 wire n_30332;
 wire n_30357;
 wire n_30452;
 wire n_30453;
 wire n_30469;
 wire n_30471;
 wire n_30472;
 wire n_30483;
 wire n_306;
 wire n_30616;
 wire n_3063;
 wire n_307;
 wire n_3077;
 wire n_3081;
 wire n_310;
 wire n_31056;
 wire n_31057;
 wire n_31058;
 wire n_31078;
 wire n_31107;
 wire n_31127;
 wire n_31128;
 wire n_31129;
 wire n_31190;
 wire n_31191;
 wire n_312;
 wire n_31227;
 wire n_31228;
 wire n_31272;
 wire n_31273;
 wire n_31311;
 wire n_31396;
 wire n_31397;
 wire n_31445;
 wire n_31455;
 wire n_31460;
 wire n_31464;
 wire n_31534;
 wire n_31535;
 wire n_31538;
 wire n_31561;
 wire n_31579;
 wire n_31581;
 wire n_316;
 wire n_317;
 wire n_31720;
 wire n_31724;
 wire n_31726;
 wire n_31732;
 wire n_31733;
 wire n_31740;
 wire n_31741;
 wire n_31742;
 wire n_31743;
 wire n_31747;
 wire n_31748;
 wire n_31750;
 wire n_31754;
 wire n_31770;
 wire n_31777;
 wire n_31779;
 wire n_31781;
 wire n_31786;
 wire n_31795;
 wire n_31801;
 wire n_31821;
 wire n_31834;
 wire n_31844;
 wire n_31849;
 wire n_31850;
 wire n_31863;
 wire n_31864;
 wire n_31865;
 wire n_31866;
 wire n_31867;
 wire n_31869;
 wire n_31870;
 wire n_31871;
 wire n_31872;
 wire n_3188;
 wire n_31886;
 wire n_31888;
 wire n_31890;
 wire n_31891;
 wire n_31892;
 wire n_31895;
 wire n_319;
 wire n_31900;
 wire n_31907;
 wire n_321;
 wire n_32162;
 wire n_32163;
 wire n_32164;
 wire n_32299;
 wire n_32300;
 wire n_32302;
 wire n_32317;
 wire n_32318;
 wire n_32319;
 wire n_32320;
 wire n_32321;
 wire n_32322;
 wire n_32323;
 wire n_32324;
 wire n_32325;
 wire n_32326;
 wire n_32327;
 wire n_32328;
 wire n_32330;
 wire n_32331;
 wire n_32332;
 wire n_32333;
 wire n_32334;
 wire n_32335;
 wire n_32336;
 wire n_32337;
 wire n_32338;
 wire n_32339;
 wire n_32341;
 wire n_32343;
 wire n_32344;
 wire n_32345;
 wire n_32346;
 wire n_32348;
 wire n_32349;
 wire n_32381;
 wire n_32382;
 wire n_32383;
 wire n_32384;
 wire n_32385;
 wire n_32386;
 wire n_32387;
 wire n_32388;
 wire n_32389;
 wire n_32390;
 wire n_32391;
 wire n_32392;
 wire n_32393;
 wire n_32394;
 wire n_32395;
 wire n_32396;
 wire n_32398;
 wire n_32399;
 wire n_32400;
 wire n_32401;
 wire n_32402;
 wire n_32403;
 wire n_32404;
 wire n_32405;
 wire n_32406;
 wire n_32407;
 wire n_32408;
 wire n_32409;
 wire n_32410;
 wire n_32411;
 wire n_32582;
 wire n_32583;
 wire n_32584;
 wire n_32585;
 wire n_32587;
 wire n_32588;
 wire n_32589;
 wire n_32590;
 wire n_32591;
 wire n_32592;
 wire n_32593;
 wire n_32595;
 wire n_32597;
 wire n_32599;
 wire n_32600;
 wire n_32601;
 wire n_32644;
 wire n_32650;
 wire n_3285;
 wire n_329;
 wire n_32916;
 wire n_33;
 wire n_330;
 wire n_33024;
 wire n_331;
 wire n_33100;
 wire n_33112;
 wire n_332;
 wire n_3320;
 wire n_33203;
 wire n_336;
 wire n_33603;
 wire n_33604;
 wire n_33644;
 wire n_3365;
 wire n_33654;
 wire n_33655;
 wire n_33656;
 wire n_33657;
 wire n_33658;
 wire n_33659;
 wire n_33660;
 wire n_33661;
 wire n_33662;
 wire n_33663;
 wire n_33664;
 wire n_33665;
 wire n_33666;
 wire n_33667;
 wire n_33668;
 wire n_33670;
 wire n_33671;
 wire n_33672;
 wire n_33673;
 wire n_33674;
 wire n_33675;
 wire n_33676;
 wire n_33677;
 wire n_33678;
 wire n_33679;
 wire n_33681;
 wire n_33682;
 wire n_33683;
 wire n_33684;
 wire n_33685;
 wire n_33686;
 wire n_33687;
 wire n_33771;
 wire n_33772;
 wire n_33774;
 wire n_33777;
 wire n_33784;
 wire n_33786;
 wire n_33787;
 wire n_33788;
 wire n_33789;
 wire n_33790;
 wire n_33791;
 wire n_33792;
 wire n_33793;
 wire n_33795;
 wire n_33796;
 wire n_3386;
 wire n_339;
 wire n_34;
 wire n_340;
 wire n_34081;
 wire n_34082;
 wire n_34098;
 wire n_34099;
 wire n_34102;
 wire n_3415;
 wire n_34190;
 wire n_3420;
 wire n_34203;
 wire n_34234;
 wire n_34235;
 wire n_3425;
 wire n_34362;
 wire n_34363;
 wire n_34377;
 wire n_34378;
 wire n_34412;
 wire n_34413;
 wire n_34420;
 wire n_34421;
 wire n_34422;
 wire n_34433;
 wire n_34434;
 wire n_34472;
 wire n_34473;
 wire n_34475;
 wire n_34479;
 wire n_34480;
 wire n_34482;
 wire n_34483;
 wire n_34484;
 wire n_34486;
 wire n_34487;
 wire n_34488;
 wire n_34490;
 wire n_34491;
 wire n_34492;
 wire n_34494;
 wire n_34495;
 wire n_34498;
 wire n_34499;
 wire n_34500;
 wire n_34502;
 wire n_34503;
 wire n_34504;
 wire n_34505;
 wire n_34506;
 wire n_34507;
 wire n_34524;
 wire n_34525;
 wire n_34526;
 wire n_3453;
 wire n_34532;
 wire n_34533;
 wire n_34534;
 wire n_34535;
 wire n_34536;
 wire n_34537;
 wire n_34538;
 wire n_34539;
 wire n_3454;
 wire n_34540;
 wire n_34541;
 wire n_3460;
 wire n_3461;
 wire n_34613;
 wire n_34614;
 wire n_34633;
 wire n_34634;
 wire n_34644;
 wire n_34645;
 wire n_34648;
 wire n_34649;
 wire n_3468;
 wire n_347;
 wire n_34837;
 wire n_34841;
 wire n_35041;
 wire n_35120;
 wire n_35121;
 wire n_35122;
 wire n_35215;
 wire n_35390;
 wire n_35391;
 wire n_35392;
 wire n_35393;
 wire n_35398;
 wire n_35399;
 wire n_35407;
 wire n_35437;
 wire n_35457;
 wire n_35458;
 wire n_35459;
 wire n_35460;
 wire n_35461;
 wire n_35462;
 wire n_35463;
 wire n_35466;
 wire n_35467;
 wire n_35468;
 wire n_35469;
 wire n_35474;
 wire n_35476;
 wire n_35550;
 wire n_35577;
 wire n_35578;
 wire n_356;
 wire n_35632;
 wire n_35633;
 wire n_35634;
 wire n_35636;
 wire n_35637;
 wire n_35638;
 wire n_35645;
 wire n_35653;
 wire n_35654;
 wire n_35655;
 wire n_35656;
 wire n_357;
 wire n_35902;
 wire n_35904;
 wire n_35908;
 wire n_35909;
 wire n_35910;
 wire n_35911;
 wire n_360;
 wire n_36007;
 wire n_36008;
 wire n_36010;
 wire n_36011;
 wire n_36012;
 wire n_36013;
 wire n_36014;
 wire n_36068;
 wire n_36071;
 wire n_36072;
 wire n_36073;
 wire n_36076;
 wire n_36077;
 wire n_36078;
 wire n_36079;
 wire n_36080;
 wire n_36081;
 wire n_36082;
 wire n_36083;
 wire n_36084;
 wire n_36085;
 wire n_36086;
 wire n_36089;
 wire n_36090;
 wire n_36091;
 wire n_36092;
 wire n_36094;
 wire n_36095;
 wire n_36097;
 wire n_36098;
 wire n_36099;
 wire n_36100;
 wire n_36101;
 wire n_36102;
 wire n_36103;
 wire n_36107;
 wire n_362;
 wire n_3621;
 wire n_36224;
 wire n_36256;
 wire n_36288;
 wire n_36289;
 wire n_36290;
 wire n_36291;
 wire n_363;
 wire n_3635;
 wire n_36361;
 wire n_36363;
 wire n_36364;
 wire n_36366;
 wire n_36367;
 wire n_3638;
 wire n_36382;
 wire n_36383;
 wire n_36385;
 wire n_36405;
 wire n_36478;
 wire n_36525;
 wire n_36528;
 wire n_36530;
 wire n_36531;
 wire n_36580;
 wire n_36581;
 wire n_36582;
 wire n_36583;
 wire n_366;
 wire n_36613;
 wire n_36628;
 wire n_36635;
 wire n_36662;
 wire n_36769;
 wire n_36770;
 wire n_36771;
 wire n_368;
 wire n_36843;
 wire n_369;
 wire n_36968;
 wire n_36969;
 wire n_3697;
 wire n_36971;
 wire n_36975;
 wire n_3698;
 wire n_3699;
 wire n_37;
 wire n_370;
 wire n_3700;
 wire n_3701;
 wire n_3702;
 wire n_3703;
 wire n_37051;
 wire n_37052;
 wire n_3709;
 wire n_3710;
 wire n_37110;
 wire n_37111;
 wire n_3712;
 wire n_3713;
 wire n_37136;
 wire n_37137;
 wire n_37138;
 wire n_37139;
 wire n_3714;
 wire n_37140;
 wire n_37141;
 wire n_37142;
 wire n_3716;
 wire n_3717;
 wire n_3718;
 wire n_3719;
 wire n_3720;
 wire n_37200;
 wire n_3721;
 wire n_3722;
 wire n_37311;
 wire n_37335;
 wire n_37336;
 wire n_37337;
 wire n_37338;
 wire n_37339;
 wire n_37340;
 wire n_37341;
 wire n_37342;
 wire n_37344;
 wire n_37350;
 wire n_37355;
 wire n_37367;
 wire n_37368;
 wire n_37381;
 wire n_37383;
 wire n_37384;
 wire n_37386;
 wire n_37387;
 wire n_374;
 wire n_37456;
 wire n_37457;
 wire n_37458;
 wire n_37459;
 wire n_37460;
 wire n_375;
 wire n_37521;
 wire n_37601;
 wire n_37606;
 wire n_37611;
 wire n_37616;
 wire n_37621;
 wire n_37626;
 wire n_379;
 wire n_37935;
 wire n_38;
 wire n_3815;
 wire n_38363;
 wire n_38364;
 wire n_38365;
 wire n_38366;
 wire n_38367;
 wire n_38368;
 wire n_38369;
 wire n_38370;
 wire n_38371;
 wire n_38373;
 wire n_38374;
 wire n_38375;
 wire n_38376;
 wire n_38377;
 wire n_38378;
 wire n_38379;
 wire n_38380;
 wire n_38381;
 wire n_38382;
 wire n_3858;
 wire n_3862;
 wire n_387;
 wire n_38705;
 wire n_38758;
 wire n_38759;
 wire n_38760;
 wire n_38761;
 wire n_38792;
 wire n_38797;
 wire n_388;
 wire n_38802;
 wire n_389;
 wire n_39;
 wire n_390;
 wire n_3900;
 wire n_3906;
 wire n_3907;
 wire n_3908;
 wire n_3909;
 wire n_391;
 wire n_3913;
 wire n_3933;
 wire n_3934;
 wire n_3935;
 wire n_3937;
 wire n_3941;
 wire n_3947;
 wire n_3948;
 wire n_3955;
 wire n_3956;
 wire n_3959;
 wire n_396;
 wire n_3985;
 wire n_399;
 wire n_3991;
 wire n_3993;
 wire n_3996;
 wire n_3999;
 wire n_4;
 wire n_40;
 wire n_4003;
 wire n_401;
 wire n_402;
 wire n_4024;
 wire n_4027;
 wire n_4028;
 wire n_40286;
 wire n_40287;
 wire n_40371;
 wire n_40372;
 wire n_40379;
 wire n_4040;
 wire n_40416;
 wire n_40417;
 wire n_40418;
 wire n_40419;
 wire n_4042;
 wire n_40420;
 wire n_40421;
 wire n_4048;
 wire n_4070;
 wire n_40712;
 wire n_4075;
 wire n_4077;
 wire n_4078;
 wire n_4081;
 wire n_4082;
 wire n_40824;
 wire n_4083;
 wire n_4084;
 wire n_4086;
 wire n_4087;
 wire n_40900;
 wire n_40902;
 wire n_40904;
 wire n_40905;
 wire n_4092;
 wire n_40954;
 wire n_40955;
 wire n_40956;
 wire n_40978;
 wire n_4098;
 wire n_40982;
 wire n_40983;
 wire n_40985;
 wire n_40986;
 wire n_40987;
 wire n_40988;
 wire n_40989;
 wire n_40990;
 wire n_40992;
 wire n_40993;
 wire n_40994;
 wire n_41;
 wire n_41034;
 wire n_4114;
 wire n_41152;
 wire n_41154;
 wire n_4116;
 wire n_4117;
 wire n_4119;
 wire n_41248;
 wire n_41323;
 wire n_41375;
 wire n_41376;
 wire n_41377;
 wire n_41378;
 wire n_41379;
 wire n_41434;
 wire n_41435;
 wire n_4146;
 wire n_41491;
 wire n_41492;
 wire n_415;
 wire n_4155;
 wire n_4156;
 wire n_41606;
 wire n_41608;
 wire n_41609;
 wire n_4161;
 wire n_41610;
 wire n_41611;
 wire n_41612;
 wire n_4162;
 wire n_41636;
 wire n_41637;
 wire n_417;
 wire n_41758;
 wire n_41759;
 wire n_41761;
 wire n_41767;
 wire n_41768;
 wire n_41769;
 wire n_4177;
 wire n_4179;
 wire n_4180;
 wire n_4186;
 wire n_419;
 wire n_41910;
 wire n_42;
 wire n_4202;
 wire n_42030;
 wire n_42031;
 wire n_4207;
 wire n_4208;
 wire n_4224;
 wire n_42248;
 wire n_42249;
 wire n_4225;
 wire n_42251;
 wire n_42252;
 wire n_42253;
 wire n_42254;
 wire n_42255;
 wire n_42256;
 wire n_42257;
 wire n_42258;
 wire n_42260;
 wire n_42261;
 wire n_42262;
 wire n_42263;
 wire n_42264;
 wire n_423;
 wire n_4230;
 wire n_4232;
 wire n_425;
 wire n_4253;
 wire n_4254;
 wire n_4258;
 wire n_4261;
 wire n_42613;
 wire n_42615;
 wire n_42616;
 wire n_42617;
 wire n_42618;
 wire n_42619;
 wire n_42620;
 wire n_42621;
 wire n_427;
 wire n_42722;
 wire n_42723;
 wire n_42724;
 wire n_42725;
 wire n_42726;
 wire n_42727;
 wire n_42728;
 wire n_42729;
 wire n_42730;
 wire n_42731;
 wire n_42732;
 wire n_42733;
 wire n_42734;
 wire n_42735;
 wire n_42736;
 wire n_42737;
 wire n_42738;
 wire n_42739;
 wire n_42740;
 wire n_4276;
 wire n_42779;
 wire n_42799;
 wire n_4280;
 wire n_42801;
 wire n_43;
 wire n_43020;
 wire n_43028;
 wire n_43075;
 wire n_43077;
 wire n_43078;
 wire n_43082;
 wire n_43083;
 wire n_43084;
 wire n_43085;
 wire n_43086;
 wire n_43087;
 wire n_43088;
 wire n_43089;
 wire n_43090;
 wire n_43091;
 wire n_43092;
 wire n_43094;
 wire n_43095;
 wire n_43096;
 wire n_43097;
 wire n_43098;
 wire n_43099;
 wire n_431;
 wire n_43100;
 wire n_4312;
 wire n_4316;
 wire n_43169;
 wire n_43170;
 wire n_43171;
 wire n_43172;
 wire n_4318;
 wire n_432;
 wire n_4320;
 wire n_43201;
 wire n_43202;
 wire n_43203;
 wire n_43204;
 wire n_43205;
 wire n_43206;
 wire n_4324;
 wire n_43281;
 wire n_43282;
 wire n_43290;
 wire n_43291;
 wire n_43305;
 wire n_43306;
 wire n_43317;
 wire n_43318;
 wire n_43319;
 wire n_4332;
 wire n_43320;
 wire n_4339;
 wire n_43394;
 wire n_43395;
 wire n_434;
 wire n_4340;
 wire n_4341;
 wire n_4342;
 wire n_4343;
 wire n_4345;
 wire n_4346;
 wire n_43467;
 wire n_43468;
 wire n_43469;
 wire n_4347;
 wire n_435;
 wire n_4350;
 wire n_4353;
 wire n_43530;
 wire n_43531;
 wire n_43533;
 wire n_43534;
 wire n_43535;
 wire n_43536;
 wire n_43537;
 wire n_4355;
 wire n_4356;
 wire n_4357;
 wire n_4359;
 wire n_43604;
 wire n_43605;
 wire n_43606;
 wire n_43607;
 wire n_4361;
 wire n_4362;
 wire n_4363;
 wire n_4364;
 wire n_4366;
 wire n_43665;
 wire n_43666;
 wire n_43667;
 wire n_4369;
 wire n_4371;
 wire n_4372;
 wire n_43720;
 wire n_43721;
 wire n_4373;
 wire n_4374;
 wire n_4375;
 wire n_43760;
 wire n_43761;
 wire n_4377;
 wire n_4379;
 wire n_4381;
 wire n_4383;
 wire n_4384;
 wire n_4390;
 wire n_4392;
 wire n_44;
 wire n_4401;
 wire n_4404;
 wire n_4405;
 wire n_4407;
 wire n_4408;
 wire n_4409;
 wire n_4410;
 wire n_4413;
 wire n_4415;
 wire n_4416;
 wire n_4418;
 wire n_442;
 wire n_4422;
 wire n_4423;
 wire n_4424;
 wire n_4425;
 wire n_4426;
 wire n_4427;
 wire n_4428;
 wire n_443;
 wire n_4430;
 wire n_4434;
 wire n_4438;
 wire n_4439;
 wire n_4441;
 wire n_4443;
 wire n_44440;
 wire n_44447;
 wire n_4445;
 wire n_44452;
 wire n_44456;
 wire n_4448;
 wire n_445;
 wire n_4450;
 wire n_4451;
 wire n_4453;
 wire n_44556;
 wire n_4456;
 wire n_4457;
 wire n_4460;
 wire n_4461;
 wire n_4462;
 wire n_4464;
 wire n_4470;
 wire n_4471;
 wire n_4472;
 wire n_4473;
 wire n_4474;
 wire n_4475;
 wire n_4481;
 wire n_4483;
 wire n_4484;
 wire n_4485;
 wire n_4486;
 wire n_44864;
 wire n_4487;
 wire n_4488;
 wire n_4489;
 wire n_4495;
 wire n_4496;
 wire n_4498;
 wire n_450;
 wire n_4500;
 wire n_4502;
 wire n_4505;
 wire n_451;
 wire n_4513;
 wire n_4514;
 wire n_4515;
 wire n_4516;
 wire n_452;
 wire n_4524;
 wire n_4525;
 wire n_4527;
 wire n_4533;
 wire n_45330;
 wire n_4534;
 wire n_4535;
 wire n_4536;
 wire n_4537;
 wire n_45388;
 wire n_454;
 wire n_4540;
 wire n_4541;
 wire n_4542;
 wire n_4544;
 wire n_4546;
 wire n_4548;
 wire n_4549;
 wire n_455;
 wire n_45569;
 wire n_4557;
 wire n_456;
 wire n_45607;
 wire n_4562;
 wire n_45624;
 wire n_45625;
 wire n_45627;
 wire n_4568;
 wire n_4572;
 wire n_4573;
 wire n_4574;
 wire n_4578;
 wire n_4579;
 wire n_4588;
 wire n_459;
 wire n_4591;
 wire n_4592;
 wire n_4593;
 wire n_4594;
 wire n_4595;
 wire n_4596;
 wire n_4597;
 wire n_4598;
 wire n_4599;
 wire n_46;
 wire n_460;
 wire n_4600;
 wire n_4603;
 wire n_4604;
 wire n_461;
 wire n_46110;
 wire n_46111;
 wire n_4614;
 wire n_46163;
 wire n_4617;
 wire n_46182;
 wire n_46183;
 wire n_46184;
 wire n_46185;
 wire n_46186;
 wire n_46187;
 wire n_46188;
 wire n_46189;
 wire n_46190;
 wire n_46191;
 wire n_46192;
 wire n_462;
 wire n_46227;
 wire n_46228;
 wire n_46229;
 wire n_46230;
 wire n_46231;
 wire n_46232;
 wire n_46233;
 wire n_46234;
 wire n_46235;
 wire n_46236;
 wire n_46237;
 wire n_46238;
 wire n_46239;
 wire n_4624;
 wire n_46240;
 wire n_46241;
 wire n_46242;
 wire n_46243;
 wire n_46244;
 wire n_46245;
 wire n_46246;
 wire n_46247;
 wire n_46248;
 wire n_46249;
 wire n_46250;
 wire n_46251;
 wire n_46252;
 wire n_46253;
 wire n_46254;
 wire n_46255;
 wire n_46256;
 wire n_46257;
 wire n_46258;
 wire n_46259;
 wire n_46260;
 wire n_46261;
 wire n_46262;
 wire n_46263;
 wire n_46289;
 wire n_463;
 wire n_46334;
 wire n_46335;
 wire n_46336;
 wire n_464;
 wire n_4641;
 wire n_46422;
 wire n_4644;
 wire n_4645;
 wire n_4646;
 wire n_46477;
 wire n_46478;
 wire n_46479;
 wire n_46480;
 wire n_46485;
 wire n_46486;
 wire n_46558;
 wire n_46559;
 wire n_4656;
 wire n_46562;
 wire n_46563;
 wire n_46564;
 wire n_46566;
 wire n_46567;
 wire n_4657;
 wire n_4658;
 wire n_46587;
 wire n_46588;
 wire n_4661;
 wire n_4662;
 wire n_4663;
 wire n_46638;
 wire n_46639;
 wire n_4664;
 wire n_46640;
 wire n_46642;
 wire n_46643;
 wire n_46644;
 wire n_4665;
 wire n_4667;
 wire n_46697;
 wire n_46698;
 wire n_467;
 wire n_4670;
 wire n_46700;
 wire n_46701;
 wire n_4671;
 wire n_4673;
 wire n_4674;
 wire n_4675;
 wire n_46750;
 wire n_468;
 wire n_4689;
 wire n_469;
 wire n_4691;
 wire n_4693;
 wire n_4695;
 wire n_47;
 wire n_4707;
 wire n_4710;
 wire n_4711;
 wire n_4712;
 wire n_47121;
 wire n_47127;
 wire n_4713;
 wire n_4715;
 wire n_47157;
 wire n_47164;
 wire n_4717;
 wire n_47184;
 wire n_4719;
 wire n_47192;
 wire n_4721;
 wire n_47217;
 wire n_47255;
 wire n_47261;
 wire n_47266;
 wire n_47287;
 wire n_47306;
 wire n_47322;
 wire n_47334;
 wire n_47340;
 wire n_47348;
 wire n_47357;
 wire n_47373;
 wire n_47390;
 wire n_47391;
 wire n_47403;
 wire n_47415;
 wire n_47498;
 wire n_47500;
 wire n_47538;
 wire n_47539;
 wire n_47540;
 wire n_47541;
 wire n_47551;
 wire n_47552;
 wire n_47553;
 wire n_47554;
 wire n_47613;
 wire n_47616;
 wire n_47631;
 wire n_47632;
 wire n_47682;
 wire n_47683;
 wire n_477;
 wire n_47706;
 wire n_47707;
 wire n_47739;
 wire n_47740;
 wire n_47767;
 wire n_47768;
 wire n_47769;
 wire n_47770;
 wire n_47771;
 wire n_47772;
 wire n_47778;
 wire n_47780;
 wire n_47786;
 wire n_47787;
 wire n_47791;
 wire n_47792;
 wire n_47793;
 wire n_47794;
 wire n_4784;
 wire n_4787;
 wire n_4788;
 wire n_4792;
 wire n_4794;
 wire n_4795;
 wire n_4798;
 wire n_48;
 wire n_48052;
 wire n_48053;
 wire n_48055;
 wire n_48056;
 wire n_48057;
 wire n_48058;
 wire n_48060;
 wire n_4807;
 wire n_48105;
 wire n_48106;
 wire n_48107;
 wire n_48109;
 wire n_48110;
 wire n_48145;
 wire n_48146;
 wire n_48147;
 wire n_48148;
 wire n_48149;
 wire n_48150;
 wire n_48151;
 wire n_48152;
 wire n_48153;
 wire n_48154;
 wire n_48155;
 wire n_48156;
 wire n_48157;
 wire n_48158;
 wire n_48159;
 wire n_48160;
 wire n_48161;
 wire n_48162;
 wire n_48163;
 wire n_48164;
 wire n_48165;
 wire n_48166;
 wire n_48167;
 wire n_48168;
 wire n_48169;
 wire n_4817;
 wire n_48170;
 wire n_48171;
 wire n_48172;
 wire n_48173;
 wire n_48174;
 wire n_48175;
 wire n_48176;
 wire n_48177;
 wire n_4818;
 wire n_4819;
 wire n_48223;
 wire n_48224;
 wire n_48225;
 wire n_4823;
 wire n_4824;
 wire n_4825;
 wire n_4826;
 wire n_4827;
 wire n_4829;
 wire n_4831;
 wire n_4832;
 wire n_4833;
 wire n_4834;
 wire n_4835;
 wire n_4840;
 wire n_48404;
 wire n_48405;
 wire n_48407;
 wire n_48412;
 wire n_48413;
 wire n_48415;
 wire n_4842;
 wire n_48423;
 wire n_48425;
 wire n_48426;
 wire n_48427;
 wire n_48428;
 wire n_48429;
 wire n_48430;
 wire n_48431;
 wire n_48432;
 wire n_48433;
 wire n_48434;
 wire n_48436;
 wire n_48437;
 wire n_4844;
 wire n_48454;
 wire n_48455;
 wire n_48456;
 wire n_4846;
 wire n_4848;
 wire n_4849;
 wire n_4850;
 wire n_4851;
 wire n_4852;
 wire n_4856;
 wire n_4858;
 wire n_4859;
 wire n_4860;
 wire n_4861;
 wire n_4862;
 wire n_48624;
 wire n_48625;
 wire n_48626;
 wire n_48627;
 wire n_48628;
 wire n_48629;
 wire n_4863;
 wire n_48630;
 wire n_48631;
 wire n_48632;
 wire n_48633;
 wire n_48634;
 wire n_48635;
 wire n_48636;
 wire n_48637;
 wire n_48638;
 wire n_48639;
 wire n_4864;
 wire n_48640;
 wire n_48642;
 wire n_48643;
 wire n_48644;
 wire n_48645;
 wire n_48646;
 wire n_48647;
 wire n_48648;
 wire n_4865;
 wire n_4867;
 wire n_48675;
 wire n_48676;
 wire n_4868;
 wire n_4869;
 wire n_487;
 wire n_4870;
 wire n_4871;
 wire n_4872;
 wire n_48729;
 wire n_4873;
 wire n_4875;
 wire n_4876;
 wire n_4877;
 wire n_4878;
 wire n_488;
 wire n_4881;
 wire n_4882;
 wire n_4883;
 wire n_4884;
 wire n_4886;
 wire n_48972;
 wire n_48974;
 wire n_4899;
 wire n_49;
 wire n_490;
 wire n_4900;
 wire n_4901;
 wire n_4902;
 wire n_4903;
 wire n_4904;
 wire n_4905;
 wire n_4906;
 wire n_4907;
 wire n_4908;
 wire n_4909;
 wire n_491;
 wire n_4910;
 wire n_4911;
 wire n_4912;
 wire n_49129;
 wire n_4913;
 wire n_49131;
 wire n_4914;
 wire n_49143;
 wire n_4915;
 wire n_4916;
 wire n_4917;
 wire n_49172;
 wire n_49173;
 wire n_49175;
 wire n_49177;
 wire n_49178;
 wire n_49179;
 wire n_4918;
 wire n_49180;
 wire n_49181;
 wire n_49182;
 wire n_4919;
 wire n_4920;
 wire n_49203;
 wire n_4922;
 wire n_4927;
 wire n_4928;
 wire n_4929;
 wire n_49309;
 wire n_49319;
 wire n_4932;
 wire n_49320;
 wire n_4933;
 wire n_4936;
 wire n_4937;
 wire n_4938;
 wire n_49387;
 wire n_4939;
 wire n_4940;
 wire n_4942;
 wire n_4945;
 wire n_49499;
 wire n_4950;
 wire n_49500;
 wire n_4952;
 wire n_4956;
 wire n_49617;
 wire n_49618;
 wire n_49619;
 wire n_49620;
 wire n_49625;
 wire n_49626;
 wire n_49641;
 wire n_497;
 wire n_49719;
 wire n_4976;
 wire n_4988;
 wire n_4990;
 wire n_4992;
 wire n_4998;
 wire n_4999;
 wire n_5;
 wire n_5000;
 wire n_5002;
 wire n_5003;
 wire n_5004;
 wire n_5005;
 wire n_5007;
 wire n_5008;
 wire n_50088;
 wire n_5009;
 wire n_50090;
 wire n_50091;
 wire n_5010;
 wire n_50109;
 wire n_5011;
 wire n_5012;
 wire n_5014;
 wire n_5015;
 wire n_5016;
 wire n_5020;
 wire n_5021;
 wire n_50217;
 wire n_50218;
 wire n_50219;
 wire n_5022;
 wire n_50220;
 wire n_50221;
 wire n_50222;
 wire n_50223;
 wire n_50224;
 wire n_50225;
 wire n_50226;
 wire n_50227;
 wire n_50228;
 wire n_50229;
 wire n_5023;
 wire n_50230;
 wire n_50231;
 wire n_50232;
 wire n_50233;
 wire n_50234;
 wire n_50235;
 wire n_50236;
 wire n_50237;
 wire n_50238;
 wire n_50239;
 wire n_5024;
 wire n_50240;
 wire n_50241;
 wire n_50242;
 wire n_50243;
 wire n_50245;
 wire n_50246;
 wire n_50247;
 wire n_50250;
 wire n_50251;
 wire n_5028;
 wire n_50287;
 wire n_50289;
 wire n_50290;
 wire n_50291;
 wire n_50292;
 wire n_50293;
 wire n_50295;
 wire n_503;
 wire n_50319;
 wire n_50341;
 wire n_50342;
 wire n_50343;
 wire n_50344;
 wire n_5036;
 wire n_50388;
 wire n_50389;
 wire n_5041;
 wire n_50426;
 wire n_50427;
 wire n_50452;
 wire n_50453;
 wire n_50454;
 wire n_50455;
 wire n_50456;
 wire n_50457;
 wire n_50458;
 wire n_50459;
 wire n_50460;
 wire n_50461;
 wire n_50463;
 wire n_5054;
 wire n_50541;
 wire n_50546;
 wire n_50548;
 wire n_50549;
 wire n_50551;
 wire n_50552;
 wire n_50553;
 wire n_50554;
 wire n_50555;
 wire n_506;
 wire n_50601;
 wire n_50602;
 wire n_50619;
 wire n_5062;
 wire n_50660;
 wire n_50702;
 wire n_50703;
 wire n_50704;
 wire n_50705;
 wire n_50706;
 wire n_50707;
 wire n_50709;
 wire n_5071;
 wire n_50710;
 wire n_50711;
 wire n_50712;
 wire n_5072;
 wire n_5073;
 wire n_5074;
 wire n_5077;
 wire n_50792;
 wire n_50793;
 wire n_50794;
 wire n_50808;
 wire n_50809;
 wire n_5081;
 wire n_50810;
 wire n_50812;
 wire n_50814;
 wire n_5082;
 wire n_5087;
 wire n_5088;
 wire n_509;
 wire n_5091;
 wire n_5093;
 wire n_5094;
 wire n_5097;
 wire n_5098;
 wire n_51;
 wire n_5100;
 wire n_5101;
 wire n_5103;
 wire n_51030;
 wire n_51032;
 wire n_51033;
 wire n_51034;
 wire n_51035;
 wire n_51036;
 wire n_51037;
 wire n_51038;
 wire n_51039;
 wire n_5104;
 wire n_51040;
 wire n_51041;
 wire n_51042;
 wire n_51045;
 wire n_51046;
 wire n_51047;
 wire n_51048;
 wire n_51049;
 wire n_5105;
 wire n_51051;
 wire n_51053;
 wire n_5106;
 wire n_5111;
 wire n_5112;
 wire n_5113;
 wire n_5114;
 wire n_51158;
 wire n_51159;
 wire n_51160;
 wire n_5118;
 wire n_512;
 wire n_5121;
 wire n_5125;
 wire n_5127;
 wire n_51288;
 wire n_5129;
 wire n_51296;
 wire n_5133;
 wire n_5135;
 wire n_5139;
 wire n_5143;
 wire n_51464;
 wire n_51478;
 wire n_51479;
 wire n_51481;
 wire n_51482;
 wire n_51483;
 wire n_51484;
 wire n_51486;
 wire n_51487;
 wire n_51488;
 wire n_51489;
 wire n_5149;
 wire n_51490;
 wire n_51493;
 wire n_51495;
 wire n_51496;
 wire n_51498;
 wire n_51499;
 wire n_51500;
 wire n_5152;
 wire n_5153;
 wire n_5154;
 wire n_5156;
 wire n_5157;
 wire n_5158;
 wire n_5159;
 wire n_5160;
 wire n_5161;
 wire n_517;
 wire n_5171;
 wire n_5172;
 wire n_5173;
 wire n_5177;
 wire n_5178;
 wire n_5181;
 wire n_5185;
 wire n_519;
 wire n_5195;
 wire n_5196;
 wire n_5197;
 wire n_5198;
 wire n_5199;
 wire n_52;
 wire n_5200;
 wire n_5201;
 wire n_5202;
 wire n_5203;
 wire n_5204;
 wire n_5207;
 wire n_5208;
 wire n_521;
 wire n_5211;
 wire n_5212;
 wire n_522;
 wire n_5221;
 wire n_5222;
 wire n_5223;
 wire n_5224;
 wire n_5225;
 wire n_523;
 wire n_5258;
 wire n_5263;
 wire n_5266;
 wire n_5267;
 wire n_5268;
 wire n_5269;
 wire n_5271;
 wire n_5272;
 wire n_5273;
 wire n_5274;
 wire n_5275;
 wire n_5276;
 wire n_52768;
 wire n_52769;
 wire n_5277;
 wire n_52770;
 wire n_5278;
 wire n_5279;
 wire n_528;
 wire n_5280;
 wire n_5281;
 wire n_5282;
 wire n_5283;
 wire n_5284;
 wire n_5285;
 wire n_5286;
 wire n_5287;
 wire n_5288;
 wire n_52880;
 wire n_5289;
 wire n_52892;
 wire n_52893;
 wire n_52895;
 wire n_52896;
 wire n_52897;
 wire n_52898;
 wire n_52899;
 wire n_529;
 wire n_5290;
 wire n_52900;
 wire n_52901;
 wire n_52902;
 wire n_52903;
 wire n_52905;
 wire n_52906;
 wire n_52907;
 wire n_52908;
 wire n_52909;
 wire n_5291;
 wire n_52910;
 wire n_52911;
 wire n_52912;
 wire n_52913;
 wire n_52914;
 wire n_52915;
 wire n_52916;
 wire n_52917;
 wire n_52918;
 wire n_52919;
 wire n_5292;
 wire n_52920;
 wire n_52921;
 wire n_52922;
 wire n_52923;
 wire n_52924;
 wire n_52926;
 wire n_5293;
 wire n_52932;
 wire n_52933;
 wire n_52934;
 wire n_52935;
 wire n_52936;
 wire n_52937;
 wire n_52938;
 wire n_52939;
 wire n_5294;
 wire n_52940;
 wire n_52948;
 wire n_52949;
 wire n_5295;
 wire n_52950;
 wire n_52951;
 wire n_5296;
 wire n_5297;
 wire n_52978;
 wire n_52979;
 wire n_5298;
 wire n_5299;
 wire n_53;
 wire n_5300;
 wire n_53002;
 wire n_53003;
 wire n_5301;
 wire n_5302;
 wire n_5303;
 wire n_5304;
 wire n_5305;
 wire n_5306;
 wire n_5307;
 wire n_5308;
 wire n_5309;
 wire n_5310;
 wire n_53101;
 wire n_53102;
 wire n_5311;
 wire n_5312;
 wire n_5313;
 wire n_5314;
 wire n_5315;
 wire n_5316;
 wire n_5317;
 wire n_5318;
 wire n_5319;
 wire n_532;
 wire n_5320;
 wire n_5321;
 wire n_5322;
 wire n_5323;
 wire n_5324;
 wire n_5325;
 wire n_5326;
 wire n_53263;
 wire n_53264;
 wire n_5327;
 wire n_5328;
 wire n_5329;
 wire n_5330;
 wire n_5331;
 wire n_5332;
 wire n_5333;
 wire n_5335;
 wire n_5336;
 wire n_53365;
 wire n_53366;
 wire n_53367;
 wire n_53368;
 wire n_53369;
 wire n_5337;
 wire n_53370;
 wire n_53371;
 wire n_53372;
 wire n_5338;
 wire n_534;
 wire n_5340;
 wire n_5341;
 wire n_5343;
 wire n_5344;
 wire n_5345;
 wire n_5346;
 wire n_5347;
 wire n_5348;
 wire n_5349;
 wire n_5350;
 wire n_5351;
 wire n_5352;
 wire n_5353;
 wire n_5354;
 wire n_5355;
 wire n_5356;
 wire n_5357;
 wire n_5358;
 wire n_5359;
 wire n_5360;
 wire n_5361;
 wire n_5362;
 wire n_5363;
 wire n_5364;
 wire n_5365;
 wire n_5366;
 wire n_5367;
 wire n_5368;
 wire n_5369;
 wire n_5370;
 wire n_5371;
 wire n_5372;
 wire n_5373;
 wire n_5374;
 wire n_5375;
 wire n_5376;
 wire n_5377;
 wire n_5378;
 wire n_5379;
 wire n_5380;
 wire n_5381;
 wire n_5382;
 wire n_5383;
 wire n_5384;
 wire n_5385;
 wire n_5386;
 wire n_5387;
 wire n_5388;
 wire n_5389;
 wire n_5390;
 wire n_5391;
 wire n_5392;
 wire n_5393;
 wire n_5394;
 wire n_5395;
 wire n_5396;
 wire n_5397;
 wire n_5398;
 wire n_5399;
 wire n_5400;
 wire n_5401;
 wire n_5402;
 wire n_5403;
 wire n_5404;
 wire n_5405;
 wire n_5406;
 wire n_5407;
 wire n_5408;
 wire n_5409;
 wire n_5410;
 wire n_5411;
 wire n_5412;
 wire n_5413;
 wire n_5414;
 wire n_5415;
 wire n_5416;
 wire n_5417;
 wire n_5418;
 wire n_5419;
 wire n_5420;
 wire n_5421;
 wire n_5422;
 wire n_5423;
 wire n_5424;
 wire n_5425;
 wire n_5426;
 wire n_5427;
 wire n_5428;
 wire n_5429;
 wire n_543;
 wire n_5430;
 wire n_5431;
 wire n_5432;
 wire n_5433;
 wire n_5434;
 wire n_5435;
 wire n_5436;
 wire n_5437;
 wire n_5438;
 wire n_5439;
 wire n_5440;
 wire n_5441;
 wire n_5442;
 wire n_5443;
 wire n_5444;
 wire n_5445;
 wire n_5446;
 wire n_5447;
 wire n_5448;
 wire n_5449;
 wire n_5450;
 wire n_5451;
 wire n_5452;
 wire n_5453;
 wire n_5454;
 wire n_5455;
 wire n_5456;
 wire n_54564;
 wire n_54566;
 wire n_5457;
 wire n_5458;
 wire n_5459;
 wire n_5460;
 wire n_5461;
 wire n_5462;
 wire n_5463;
 wire n_5464;
 wire n_5465;
 wire n_5466;
 wire n_5467;
 wire n_5468;
 wire n_5469;
 wire n_5470;
 wire n_5471;
 wire n_5472;
 wire n_5473;
 wire n_5474;
 wire n_5475;
 wire n_5476;
 wire n_5477;
 wire n_5478;
 wire n_5479;
 wire n_5480;
 wire n_5481;
 wire n_5482;
 wire n_5483;
 wire n_5484;
 wire n_5485;
 wire n_5486;
 wire n_5487;
 wire n_5488;
 wire n_5489;
 wire n_549;
 wire n_5490;
 wire n_5491;
 wire n_5492;
 wire n_5493;
 wire n_5494;
 wire n_5495;
 wire n_5496;
 wire n_5497;
 wire n_5498;
 wire n_5499;
 wire n_55;
 wire n_550;
 wire n_5500;
 wire n_5501;
 wire n_5502;
 wire n_5503;
 wire n_5504;
 wire n_5505;
 wire n_5506;
 wire n_5507;
 wire n_5508;
 wire n_5509;
 wire n_5510;
 wire n_5511;
 wire n_5512;
 wire n_5513;
 wire n_5514;
 wire n_5515;
 wire n_5516;
 wire n_5517;
 wire n_5518;
 wire n_5519;
 wire n_552;
 wire n_5520;
 wire n_5521;
 wire n_5522;
 wire n_5523;
 wire n_5524;
 wire n_5525;
 wire n_5526;
 wire n_5527;
 wire n_5528;
 wire n_5529;
 wire n_5530;
 wire n_5532;
 wire n_5533;
 wire n_5534;
 wire n_5536;
 wire n_5537;
 wire n_556;
 wire n_557;
 wire n_56;
 wire n_560;
 wire n_56056;
 wire n_56057;
 wire n_56059;
 wire n_56060;
 wire n_56062;
 wire n_5674;
 wire n_56842;
 wire n_56844;
 wire n_56845;
 wire n_56846;
 wire n_56847;
 wire n_56848;
 wire n_56849;
 wire n_56850;
 wire n_56851;
 wire n_56852;
 wire n_56853;
 wire n_56854;
 wire n_56855;
 wire n_56856;
 wire n_56857;
 wire n_56858;
 wire n_56859;
 wire n_56860;
 wire n_56861;
 wire n_56863;
 wire n_56864;
 wire n_56865;
 wire n_56866;
 wire n_56867;
 wire n_56868;
 wire n_56869;
 wire n_5687;
 wire n_56870;
 wire n_56871;
 wire n_56879;
 wire n_56881;
 wire n_5691;
 wire n_57;
 wire n_57041;
 wire n_5706;
 wire n_57084;
 wire n_57289;
 wire n_573;
 wire n_5741;
 wire n_5748;
 wire n_57733;
 wire n_57758;
 wire n_57759;
 wire n_57760;
 wire n_5789;
 wire n_57963;
 wire n_57964;
 wire n_57965;
 wire n_57966;
 wire n_58;
 wire n_58150;
 wire n_5845;
 wire n_5846;
 wire n_5847;
 wire n_5848;
 wire n_5849;
 wire n_58646;
 wire n_58647;
 wire n_58648;
 wire n_58649;
 wire n_58650;
 wire n_58710;
 wire n_58734;
 wire n_58735;
 wire n_588;
 wire n_589;
 wire n_58959;
 wire n_58960;
 wire n_59;
 wire n_59252;
 wire n_59256;
 wire n_59338;
 wire n_59339;
 wire n_59340;
 wire n_59341;
 wire n_59474;
 wire n_59476;
 wire n_59477;
 wire n_59639;
 wire n_59640;
 wire n_59641;
 wire n_59642;
 wire n_59643;
 wire n_59644;
 wire n_597;
 wire n_59759;
 wire n_59763;
 wire n_59764;
 wire n_6;
 wire n_603;
 wire n_6044;
 wire n_60456;
 wire n_6051;
 wire n_60588;
 wire n_6065;
 wire n_607;
 wire n_6071;
 wire n_608;
 wire n_60873;
 wire n_60874;
 wire n_6115;
 wire n_6122;
 wire n_61228;
 wire n_61229;
 wire n_61242;
 wire n_61243;
 wire n_61244;
 wire n_61245;
 wire n_6136;
 wire n_6138;
 wire n_6141;
 wire n_6144;
 wire n_6146;
 wire n_616;
 wire n_61773;
 wire n_61785;
 wire n_61786;
 wire n_61883;
 wire n_61885;
 wire n_61887;
 wire n_61889;
 wire n_61895;
 wire n_61901;
 wire n_61957;
 wire n_61963;
 wire n_62;
 wire n_62124;
 wire n_6232;
 wire n_624;
 wire n_6242;
 wire n_6248;
 wire n_6249;
 wire n_625;
 wire n_62612;
 wire n_62613;
 wire n_62614;
 wire n_62615;
 wire n_62634;
 wire n_62657;
 wire n_62717;
 wire n_62718;
 wire n_62918;
 wire n_62919;
 wire n_62920;
 wire n_62940;
 wire n_6295;
 wire n_6297;
 wire n_6299;
 wire n_63;
 wire n_6301;
 wire n_633;
 wire n_634;
 wire n_635;
 wire n_636;
 wire n_63778;
 wire n_63785;
 wire n_63786;
 wire n_63999;
 wire n_64;
 wire n_640;
 wire n_64000;
 wire n_64014;
 wire n_64102;
 wire n_64103;
 wire n_64133;
 wire n_64191;
 wire n_64192;
 wire n_64296;
 wire n_64297;
 wire n_643;
 wire n_644;
 wire n_64672;
 wire n_64696;
 wire n_64697;
 wire n_64708;
 wire n_64709;
 wire n_64710;
 wire n_64711;
 wire n_64713;
 wire n_64714;
 wire n_64715;
 wire n_64716;
 wire n_64744;
 wire n_64745;
 wire n_64793;
 wire n_64794;
 wire n_64812;
 wire n_64813;
 wire n_64814;
 wire n_64816;
 wire n_64817;
 wire n_64818;
 wire n_64819;
 wire n_64833;
 wire n_64834;
 wire n_64847;
 wire n_64848;
 wire n_64849;
 wire n_64851;
 wire n_64852;
 wire n_64853;
 wire n_64854;
 wire n_64855;
 wire n_64856;
 wire n_64861;
 wire n_64862;
 wire n_64974;
 wire n_64993;
 wire n_64994;
 wire n_64995;
 wire n_64996;
 wire n_64997;
 wire n_64998;
 wire n_65;
 wire n_65000;
 wire n_65001;
 wire n_65029;
 wire n_65030;
 wire n_65053;
 wire n_65054;
 wire n_65055;
 wire n_65056;
 wire n_65057;
 wire n_65058;
 wire n_65236;
 wire n_65238;
 wire n_65239;
 wire n_65240;
 wire n_65241;
 wire n_65242;
 wire n_65243;
 wire n_65244;
 wire n_65245;
 wire n_65246;
 wire n_65247;
 wire n_65248;
 wire n_65249;
 wire n_65250;
 wire n_65251;
 wire n_65252;
 wire n_65253;
 wire n_65254;
 wire n_65255;
 wire n_65256;
 wire n_65257;
 wire n_65258;
 wire n_65260;
 wire n_65261;
 wire n_65262;
 wire n_65263;
 wire n_65265;
 wire n_65266;
 wire n_65267;
 wire n_65268;
 wire n_65269;
 wire n_65270;
 wire n_65292;
 wire n_65293;
 wire n_65297;
 wire n_65298;
 wire n_65325;
 wire n_65326;
 wire n_65327;
 wire n_65328;
 wire n_65329;
 wire n_65395;
 wire n_655;
 wire n_6552;
 wire n_65577;
 wire n_65578;
 wire n_65642;
 wire n_65643;
 wire n_65644;
 wire n_65645;
 wire n_65646;
 wire n_65763;
 wire n_65764;
 wire n_6583;
 wire n_65879;
 wire n_65895;
 wire n_65896;
 wire n_65897;
 wire n_65898;
 wire n_65899;
 wire n_659;
 wire n_65900;
 wire n_65902;
 wire n_65905;
 wire n_65906;
 wire n_65908;
 wire n_65910;
 wire n_65911;
 wire n_65912;
 wire n_65914;
 wire n_65915;
 wire n_65917;
 wire n_65918;
 wire n_65919;
 wire n_65920;
 wire n_65921;
 wire n_65922;
 wire n_65924;
 wire n_65925;
 wire n_65927;
 wire n_65928;
 wire n_65929;
 wire n_65930;
 wire n_65931;
 wire n_65932;
 wire n_65933;
 wire n_65934;
 wire n_65936;
 wire n_65937;
 wire n_65941;
 wire n_65947;
 wire n_65948;
 wire n_65949;
 wire n_65950;
 wire n_65951;
 wire n_65952;
 wire n_65953;
 wire n_65954;
 wire n_65955;
 wire n_65958;
 wire n_65959;
 wire n_65961;
 wire n_65962;
 wire n_65964;
 wire n_65965;
 wire n_65967;
 wire n_65968;
 wire n_65969;
 wire n_65970;
 wire n_65971;
 wire n_65972;
 wire n_65975;
 wire n_65977;
 wire n_65978;
 wire n_65980;
 wire n_65983;
 wire n_65984;
 wire n_65989;
 wire n_65990;
 wire n_65992;
 wire n_65993;
 wire n_65995;
 wire n_65996;
 wire n_65997;
 wire n_65998;
 wire n_65999;
 wire n_66;
 wire n_660;
 wire n_66000;
 wire n_66001;
 wire n_66002;
 wire n_66003;
 wire n_66004;
 wire n_66005;
 wire n_66007;
 wire n_66008;
 wire n_66010;
 wire n_66011;
 wire n_66014;
 wire n_66015;
 wire n_66016;
 wire n_66017;
 wire n_66023;
 wire n_66024;
 wire n_66025;
 wire n_66026;
 wire n_66030;
 wire n_66031;
 wire n_66032;
 wire n_66054;
 wire n_66076;
 wire n_6615;
 wire n_6616;
 wire n_66198;
 wire n_66199;
 wire n_666;
 wire n_66658;
 wire n_66659;
 wire n_66660;
 wire n_66661;
 wire n_66662;
 wire n_66663;
 wire n_66664;
 wire n_66665;
 wire n_66666;
 wire n_66667;
 wire n_66668;
 wire n_66669;
 wire n_66670;
 wire n_66671;
 wire n_66672;
 wire n_66673;
 wire n_66674;
 wire n_66675;
 wire n_66676;
 wire n_66677;
 wire n_66678;
 wire n_66679;
 wire n_66680;
 wire n_66681;
 wire n_66682;
 wire n_66683;
 wire n_66799;
 wire n_66801;
 wire n_66802;
 wire n_66803;
 wire n_66804;
 wire n_66805;
 wire n_66806;
 wire n_66807;
 wire n_66808;
 wire n_66809;
 wire n_66810;
 wire n_66812;
 wire n_66813;
 wire n_66814;
 wire n_66815;
 wire n_66816;
 wire n_66817;
 wire n_66818;
 wire n_66819;
 wire n_66820;
 wire n_66821;
 wire n_66822;
 wire n_66824;
 wire n_66825;
 wire n_66826;
 wire n_66827;
 wire n_66828;
 wire n_66829;
 wire n_66830;
 wire n_66831;
 wire n_66832;
 wire n_66833;
 wire n_66834;
 wire n_66835;
 wire n_66842;
 wire n_66843;
 wire n_66855;
 wire n_66856;
 wire n_66868;
 wire n_66869;
 wire n_66881;
 wire n_67;
 wire n_670;
 wire n_672;
 wire n_6721;
 wire n_67246;
 wire n_67247;
 wire n_67248;
 wire n_67249;
 wire n_6732;
 wire n_67328;
 wire n_67329;
 wire n_6748;
 wire n_67490;
 wire n_675;
 wire n_67546;
 wire n_67568;
 wire n_678;
 wire n_68;
 wire n_68207;
 wire n_68211;
 wire n_68212;
 wire n_68215;
 wire n_68217;
 wire n_68219;
 wire n_68221;
 wire n_68223;
 wire n_68227;
 wire n_68229;
 wire n_68231;
 wire n_684;
 wire n_69;
 wire n_69010;
 wire n_69011;
 wire n_69012;
 wire n_69013;
 wire n_69014;
 wire n_69015;
 wire n_69016;
 wire n_69017;
 wire n_69018;
 wire n_69019;
 wire n_69020;
 wire n_69021;
 wire n_69022;
 wire n_69023;
 wire n_69024;
 wire n_69025;
 wire n_69026;
 wire n_69027;
 wire n_69028;
 wire n_69029;
 wire n_695;
 wire n_6956;
 wire n_696;
 wire n_6960;
 wire n_6961;
 wire n_6972;
 wire n_69795;
 wire n_69796;
 wire n_698;
 wire n_7;
 wire n_70;
 wire n_700;
 wire n_70038;
 wire n_70039;
 wire n_70040;
 wire n_70042;
 wire n_70043;
 wire n_70044;
 wire n_70045;
 wire n_70046;
 wire n_70047;
 wire n_70048;
 wire n_70050;
 wire n_70051;
 wire n_70052;
 wire n_70053;
 wire n_70054;
 wire n_70055;
 wire n_70056;
 wire n_70057;
 wire n_70058;
 wire n_70059;
 wire n_70060;
 wire n_70061;
 wire n_70062;
 wire n_70063;
 wire n_70064;
 wire n_70065;
 wire n_70066;
 wire n_70067;
 wire n_70068;
 wire n_70069;
 wire n_70070;
 wire n_70071;
 wire n_70072;
 wire n_70198;
 wire n_70199;
 wire n_70200;
 wire n_70201;
 wire n_70240;
 wire n_70241;
 wire n_703;
 wire n_70322;
 wire n_70323;
 wire n_70324;
 wire n_70325;
 wire n_70326;
 wire n_70411;
 wire n_70413;
 wire n_70414;
 wire n_70415;
 wire n_705;
 wire n_706;
 wire n_70621;
 wire n_70622;
 wire n_70648;
 wire n_70649;
 wire n_707;
 wire n_7082;
 wire n_7083;
 wire n_7084;
 wire n_7086;
 wire n_7087;
 wire n_70885;
 wire n_70886;
 wire n_70887;
 wire n_7089;
 wire n_709;
 wire n_71;
 wire n_710;
 wire n_713;
 wire n_7132;
 wire n_71350;
 wire n_71351;
 wire n_71352;
 wire n_71390;
 wire n_71391;
 wire n_71392;
 wire n_71393;
 wire n_71394;
 wire n_71395;
 wire n_714;
 wire n_7152;
 wire n_7167;
 wire n_7168;
 wire n_7169;
 wire n_7170;
 wire n_7171;
 wire n_7172;
 wire n_7173;
 wire n_7174;
 wire n_7175;
 wire n_7176;
 wire n_719;
 wire n_7195;
 wire n_7196;
 wire n_71971;
 wire n_71972;
 wire n_71973;
 wire n_71974;
 wire n_72;
 wire n_720;
 wire n_7202;
 wire n_7204;
 wire n_72057;
 wire n_72058;
 wire n_72059;
 wire n_7206;
 wire n_72060;
 wire n_72061;
 wire n_72062;
 wire n_72063;
 wire n_72064;
 wire n_72065;
 wire n_7207;
 wire n_7208;
 wire n_72081;
 wire n_72082;
 wire n_72083;
 wire n_72084;
 wire n_72087;
 wire n_7209;
 wire n_7212;
 wire n_7215;
 wire n_7216;
 wire n_7218;
 wire n_7219;
 wire n_7221;
 wire n_7222;
 wire n_7225;
 wire n_7226;
 wire n_7227;
 wire n_72307;
 wire n_72308;
 wire n_7231;
 wire n_7249;
 wire n_725;
 wire n_7251;
 wire n_7270;
 wire n_728;
 wire n_7285;
 wire n_7288;
 wire n_729;
 wire n_72908;
 wire n_72909;
 wire n_73;
 wire n_7308;
 wire n_73154;
 wire n_73169;
 wire n_73170;
 wire n_73171;
 wire n_73172;
 wire n_73173;
 wire n_73174;
 wire n_73175;
 wire n_73176;
 wire n_73177;
 wire n_7319;
 wire n_73300;
 wire n_73301;
 wire n_73302;
 wire n_73303;
 wire n_73304;
 wire n_73305;
 wire n_73306;
 wire n_73307;
 wire n_73308;
 wire n_73309;
 wire n_73310;
 wire n_73311;
 wire n_73312;
 wire n_73313;
 wire n_73314;
 wire n_7335;
 wire n_73388;
 wire n_73399;
 wire n_73400;
 wire n_736;
 wire n_737;
 wire n_73996;
 wire n_73997;
 wire n_73999;
 wire n_74;
 wire n_7408;
 wire n_7410;
 wire n_7411;
 wire n_7414;
 wire n_7417;
 wire n_7418;
 wire n_742;
 wire n_7426;
 wire n_7430;
 wire n_744;
 wire n_7442;
 wire n_7486;
 wire n_7491;
 wire n_75;
 wire n_7500;
 wire n_7501;
 wire n_7502;
 wire n_7510;
 wire n_7511;
 wire n_7514;
 wire n_752;
 wire n_7522;
 wire n_7523;
 wire n_7524;
 wire n_7526;
 wire n_7527;
 wire n_7538;
 wire n_7541;
 wire n_7542;
 wire n_7543;
 wire n_7544;
 wire n_7562;
 wire n_7563;
 wire n_7564;
 wire n_7567;
 wire n_7569;
 wire n_7570;
 wire n_7571;
 wire n_7572;
 wire n_75733;
 wire n_75734;
 wire n_75735;
 wire n_75736;
 wire n_75792;
 wire n_75793;
 wire n_75794;
 wire n_75795;
 wire n_7582;
 wire n_7586;
 wire n_7588;
 wire n_7589;
 wire n_759;
 wire n_7597;
 wire n_76;
 wire n_76054;
 wire n_76055;
 wire n_76056;
 wire n_761;
 wire n_7641;
 wire n_7653;
 wire n_7656;
 wire n_7665;
 wire n_7667;
 wire n_7668;
 wire n_7671;
 wire n_7672;
 wire n_7673;
 wire n_7676;
 wire n_76763;
 wire n_76764;
 wire n_76778;
 wire n_7689;
 wire n_769;
 wire n_7691;
 wire n_7692;
 wire n_7693;
 wire n_7694;
 wire n_7695;
 wire n_76986;
 wire n_7712;
 wire n_77233;
 wire n_77234;
 wire n_7725;
 wire n_7735;
 wire n_77396;
 wire n_77397;
 wire n_77398;
 wire n_7743;
 wire n_7744;
 wire n_775;
 wire n_7753;
 wire n_7754;
 wire n_7755;
 wire n_7756;
 wire n_7766;
 wire n_7772;
 wire n_77796;
 wire n_77797;
 wire n_778;
 wire n_7781;
 wire n_77853;
 wire n_77855;
 wire n_7788;
 wire n_77964;
 wire n_7800;
 wire n_78002;
 wire n_7803;
 wire n_78040;
 wire n_78041;
 wire n_78042;
 wire n_78043;
 wire n_78044;
 wire n_78045;
 wire n_7806;
 wire n_78094;
 wire n_78134;
 wire n_78135;
 wire n_78137;
 wire n_78138;
 wire n_78139;
 wire n_78140;
 wire n_78141;
 wire n_78164;
 wire n_78166;
 wire n_78167;
 wire n_782;
 wire n_78273;
 wire n_78274;
 wire n_78275;
 wire n_78276;
 wire n_78410;
 wire n_78411;
 wire n_7859;
 wire n_786;
 wire n_78621;
 wire n_78622;
 wire n_7863;
 wire n_78683;
 wire n_78684;
 wire n_78685;
 wire n_78686;
 wire n_7869;
 wire n_7872;
 wire n_7881;
 wire n_78810;
 wire n_78813;
 wire n_7883;
 wire n_7888;
 wire n_78930;
 wire n_78931;
 wire n_78932;
 wire n_78933;
 wire n_78934;
 wire n_78935;
 wire n_78936;
 wire n_78937;
 wire n_78938;
 wire n_78939;
 wire n_78940;
 wire n_78941;
 wire n_78942;
 wire n_78943;
 wire n_78944;
 wire n_78945;
 wire n_78946;
 wire n_78947;
 wire n_78948;
 wire n_78949;
 wire n_78950;
 wire n_78951;
 wire n_78952;
 wire n_78953;
 wire n_78954;
 wire n_78955;
 wire n_78956;
 wire n_78957;
 wire n_78958;
 wire n_78959;
 wire n_79;
 wire n_79016;
 wire n_79017;
 wire n_79019;
 wire n_79103;
 wire n_79104;
 wire n_79167;
 wire n_79168;
 wire n_79175;
 wire n_79176;
 wire n_79177;
 wire n_79178;
 wire n_79179;
 wire n_79192;
 wire n_79193;
 wire n_79194;
 wire n_79195;
 wire n_79196;
 wire n_79197;
 wire n_79198;
 wire n_79199;
 wire n_79200;
 wire n_79201;
 wire n_79202;
 wire n_79203;
 wire n_79204;
 wire n_79205;
 wire n_79206;
 wire n_79207;
 wire n_79208;
 wire n_7927;
 wire n_79305;
 wire n_79306;
 wire n_79307;
 wire n_79308;
 wire n_79326;
 wire n_79327;
 wire n_7939;
 wire n_7941;
 wire n_7942;
 wire n_798;
 wire n_7990;
 wire n_7994;
 wire n_7995;
 wire n_7997;
 wire n_79971;
 wire n_79972;
 wire n_79973;
 wire n_7999;
 wire n_8;
 wire n_80;
 wire n_8005;
 wire n_8006;
 wire n_8007;
 wire n_8008;
 wire n_801;
 wire n_8012;
 wire n_8013;
 wire n_805;
 wire n_806;
 wire n_81;
 wire n_811;
 wire n_8111;
 wire n_8112;
 wire n_8113;
 wire n_8117;
 wire n_8118;
 wire n_8119;
 wire n_8123;
 wire n_8124;
 wire n_8128;
 wire n_8173;
 wire n_8174;
 wire n_8175;
 wire n_8177;
 wire n_8183;
 wire n_8186;
 wire n_8189;
 wire n_8191;
 wire n_8192;
 wire n_8212;
 wire n_8220;
 wire n_8228;
 wire n_8232;
 wire n_8234;
 wire n_8235;
 wire n_8236;
 wire n_8238;
 wire n_8242;
 wire n_8246;
 wire n_8247;
 wire n_8248;
 wire n_8251;
 wire n_8252;
 wire n_8255;
 wire n_8256;
 wire n_8262;
 wire n_8278;
 wire n_8279;
 wire n_8280;
 wire n_8296;
 wire n_8299;
 wire n_83;
 wire n_8301;
 wire n_8306;
 wire n_8307;
 wire n_8308;
 wire n_8309;
 wire n_8311;
 wire n_8313;
 wire n_8314;
 wire n_8315;
 wire n_8319;
 wire n_8320;
 wire n_8321;
 wire n_8332;
 wire n_8333;
 wire n_8334;
 wire n_8336;
 wire n_8337;
 wire n_8338;
 wire n_8339;
 wire n_8340;
 wire n_8341;
 wire n_8351;
 wire n_8354;
 wire n_8357;
 wire n_8360;
 wire n_8363;
 wire n_8366;
 wire n_8369;
 wire n_8372;
 wire n_8375;
 wire n_8378;
 wire n_84;
 wire n_842;
 wire n_8443;
 wire n_8446;
 wire n_8449;
 wire n_8452;
 wire n_8464;
 wire n_8469;
 wire n_8474;
 wire n_8479;
 wire n_8484;
 wire n_8489;
 wire n_8494;
 wire n_8499;
 wire n_8504;
 wire n_8509;
 wire n_8514;
 wire n_8519;
 wire n_8524;
 wire n_8529;
 wire n_8534;
 wire n_8539;
 wire n_8544;
 wire n_8549;
 wire n_8554;
 wire n_8559;
 wire n_8564;
 wire n_8569;
 wire n_8574;
 wire n_8579;
 wire n_8584;
 wire n_8589;
 wire n_8594;
 wire n_8599;
 wire n_86;
 wire n_8604;
 wire n_8609;
 wire n_8614;
 wire n_8619;
 wire n_8624;
 wire n_8634;
 wire n_8638;
 wire n_8643;
 wire n_8648;
 wire n_8653;
 wire n_8658;
 wire n_8664;
 wire n_8668;
 wire n_8674;
 wire n_8678;
 wire n_8683;
 wire n_8688;
 wire n_88;
 wire n_89;
 wire n_9;
 wire n_90;
 wire n_908;
 wire n_9294;
 wire n_9295;
 wire n_9296;
 wire n_9297;
 wire n_9298;
 wire n_9299;
 wire n_93;
 wire n_9300;
 wire n_9301;
 wire n_933;
 wire n_9344;
 wire n_9345;
 wire n_9346;
 wire n_9347;
 wire n_9348;
 wire n_9349;
 wire n_9350;
 wire n_9351;
 wire n_9394;
 wire n_9395;
 wire n_9396;
 wire n_9397;
 wire n_9398;
 wire n_94;
 wire n_9466;
 wire n_9467;
 wire n_9468;
 wire n_9476;
 wire n_95;
 wire n_9555;
 wire n_9629;
 wire n_9630;
 wire n_9650;
 wire n_9654;
 wire n_9663;
 wire n_9665;
 wire n_9682;
 wire n_9686;
 wire n_97;
 wire n_9701;
 wire n_9703;
 wire n_9711;
 wire n_9713;
 wire n_9717;
 wire n_9721;
 wire n_9722;
 wire n_9723;
 wire n_9726;
 wire n_9727;
 wire n_9731;
 wire n_9735;
 wire n_9738;
 wire n_9742;
 wire n_9745;
 wire n_9747;
 wire n_9751;
 wire n_9752;
 wire n_9755;
 wire n_9756;
 wire n_9757;
 wire n_9760;
 wire n_9767;
 wire n_9772;
 wire n_9774;
 wire n_9776;
 wire n_9780;
 wire n_9781;
 wire n_9784;
 wire n_9785;
 wire n_9786;
 wire n_9790;
 wire n_9793;
 wire n_9800;
 wire n_9802;
 wire n_9804;
 wire n_9808;
 wire n_9810;
 wire n_9811;
 wire n_9814;
 wire n_9815;
 wire n_9817;
 wire n_9822;
 wire n_9828;
 wire n_9832;
 wire n_9834;
 wire n_9838;
 wire n_9840;
 wire n_9841;
 wire n_9843;
 wire n_9844;
 wire n_9849;
 wire n_9851;
 wire n_9857;
 wire n_9860;
 wire n_9863;
 wire n_9867;
 wire n_9869;
 wire n_9870;
 wire n_9873;
 wire n_9874;
 wire n_9877;
 wire n_9880;
 wire n_9886;
 wire n_9889;
 wire n_9892;
 wire n_9896;
 wire n_9898;
 wire n_9899;
 wire n_99;
 wire n_9902;
 wire n_9903;
 wire n_9907;
 wire n_9909;
 wire n_9914;
 wire n_9922;
 wire n_9926;
 wire n_9930;
 wire n_9936;
 wire n_9938;
 wire n_9941;
 wire n_9942;
 wire n_9944;
 wire n_9949;
 wire n_9954;
 wire n_9957;
 wire n_9958;
 wire n_9959;
 wire n_9960;
 wire n_9963;
 wire n_9967;
 wire n_9996;
 wire o3_empty;
 wire o3_we;
 wire o4_empty;
 wire o4_we;
 wire o6_empty;
 wire o6_we;
 wire o7_empty;
 wire o7_we;
 wire o8_empty;
 wire o8_we;
 wire o9_empty;
 wire o9_we;
 wire resume_req;
 wire rf_we;
 wire u12_re1;
 wire u12_re2;
 wire u12_wb_ack_o_745;
 wire \u12_wb_data_o[0]_713 ;
 wire \u12_wb_data_o[10]_723 ;
 wire \u12_wb_data_o[11]_724 ;
 wire \u12_wb_data_o[12]_725 ;
 wire \u12_wb_data_o[13]_726 ;
 wire \u12_wb_data_o[14]_727 ;
 wire \u12_wb_data_o[15]_728 ;
 wire \u12_wb_data_o[16]_729 ;
 wire \u12_wb_data_o[17]_730 ;
 wire \u12_wb_data_o[18]_731 ;
 wire \u12_wb_data_o[19]_732 ;
 wire \u12_wb_data_o[1]_714 ;
 wire \u12_wb_data_o[20]_733 ;
 wire \u12_wb_data_o[21]_734 ;
 wire \u12_wb_data_o[22]_735 ;
 wire \u12_wb_data_o[23]_736 ;
 wire \u12_wb_data_o[24]_737 ;
 wire \u12_wb_data_o[25]_738 ;
 wire \u12_wb_data_o[26]_739 ;
 wire \u12_wb_data_o[27]_740 ;
 wire \u12_wb_data_o[28]_741 ;
 wire \u12_wb_data_o[29]_742 ;
 wire \u12_wb_data_o[2]_715 ;
 wire \u12_wb_data_o[30]_743 ;
 wire \u12_wb_data_o[31]_744 ;
 wire \u12_wb_data_o[3]_716 ;
 wire \u12_wb_data_o[4]_717 ;
 wire \u12_wb_data_o[5]_718 ;
 wire \u12_wb_data_o[6]_719 ;
 wire \u12_wb_data_o[7]_720 ;
 wire \u12_wb_data_o[8]_721 ;
 wire \u12_wb_data_o[9]_722 ;
 wire u12_we1;
 wire u12_we2;
 wire u13_int_1643;
 wire u14_u0_en_out_l2;
 wire u14_u0_full_empty_r;
 wire u14_u1_en_out_l2;
 wire u14_u1_full_empty_r;
 wire u14_u2_en_out_l2;
 wire u14_u2_full_empty_r;
 wire u14_u3_en_out_l2;
 wire u14_u3_full_empty_r;
 wire u14_u4_en_out_l2;
 wire u14_u4_full_empty_r;
 wire u14_u5_en_out_l2;
 wire u14_u5_full_empty_r;
 wire u14_u6_en_out_l2;
 wire u14_u6_en_out_l_44;
 wire u14_u6_full_empty_r;
 wire u14_u7_en_out_l2;
 wire u14_u7_en_out_l_44;
 wire u14_u7_full_empty_r;
 wire u14_u8_en_out_l2;
 wire u14_u8_en_out_l_44;
 wire u14_u8_full_empty_r;
 wire u15_crac_rd;
 wire u15_crac_we_r;
 wire u15_rdd1;
 wire u15_rdd2;
 wire u15_rdd3;
 wire u15_valid_r;
 wire u16_u0_dma_req_52;
 wire u16_u0_dma_req_r1;
 wire u16_u1_dma_req_52;
 wire u16_u1_dma_req_r1;
 wire u16_u2_dma_req_52;
 wire u16_u2_dma_req_r1;
 wire u16_u3_dma_req_52;
 wire u16_u3_dma_req_r1;
 wire u16_u4_dma_req_52;
 wire u16_u4_dma_req_r1;
 wire u16_u5_dma_req_52;
 wire u16_u5_dma_req_r1;
 wire u16_u6_dma_req_52;
 wire u16_u6_dma_req_r1;
 wire u16_u7_dma_req_52;
 wire u16_u7_dma_req_r1;
 wire u16_u8_dma_req_52;
 wire u16_u8_dma_req_r1;
 wire u1_sdata_in_r;
 wire u26_ac97_rst_104;
 wire u2_bit_clk_e;
 wire u2_bit_clk_r;
 wire u2_bit_clk_r1;
 wire u2_sync_beat;
 wire u2_sync_resume;
 wire valid;
 wire valid_s;
 wire valid_s1;
 wire [15:0] crac_din;
 wire [31:0] crac_out;
 wire [31:0] i3_dout;
 wire [1:0] i3_status;
 wire [31:0] i4_dout;
 wire [1:0] i4_status;
 wire [31:0] i6_dout;
 wire [1:0] i6_status;
 wire [6:0] ic0_cfg;
 wire [2:0] ic0_int_set;
 wire [6:0] ic1_cfg;
 wire [2:0] ic1_int_set;
 wire [6:0] ic2_cfg;
 wire [2:0] ic2_int_set;
 wire [15:0] in_slt0;
 wire [11:0] in_slt1;
 wire [19:0] in_slt2;
 wire [19:0] in_slt3;
 wire [19:0] in_slt4;
 wire [19:0] in_slt6;
 wire [2:0] in_valid;
 wire [2:0] in_valid_s;
 wire [2:0] in_valid_s1;
 wire [1:0] o3_status;
 wire [1:0] o4_status;
 wire [1:0] o6_status;
 wire [1:0] o7_status;
 wire [1:0] o8_status;
 wire [1:0] o9_status;
 wire [6:0] oc0_cfg;
 wire [2:0] oc0_int_set;
 wire [6:0] oc1_cfg;
 wire [2:0] oc1_int_set;
 wire [6:0] oc2_cfg;
 wire [2:0] oc2_int_set;
 wire [6:0] oc3_cfg;
 wire [2:0] oc3_int_set;
 wire [6:0] oc4_cfg;
 wire [2:0] oc4_int_set;
 wire [6:0] oc5_cfg;
 wire [2:0] oc5_int_set;
 wire [5:0] out_le;
 wire [14:0] out_slt0;
 wire [19:0] out_slt3;
 wire [19:0] out_slt4;
 wire [19:0] out_slt6;
 wire [19:0] out_slt7;
 wire [19:0] out_slt8;
 wire [19:0] out_slt9;
 wire [15:0] u0_slt0_r;
 wire [19:0] u0_slt1_r;
 wire [19:0] u0_slt2_r;
 wire [19:0] u0_slt3_r;
 wire [19:0] u0_slt4_r;
 wire [19:0] u0_slt5_r;
 wire [19:0] u0_slt6_r;
 wire [19:0] u0_slt7_r;
 wire [19:0] u0_slt8_r;
 wire [19:0] u0_slt9_r;
 wire [15:0] u10_din_tmp1;
 wire [31:0] \u10_mem[0] ;
 wire [31:0] \u10_mem[1] ;
 wire [31:0] \u10_mem[2] ;
 wire [31:0] \u10_mem[3] ;
 wire [2:0] u10_rp;
 wire [3:0] u10_wp;
 wire [15:0] u11_din_tmp1;
 wire [31:0] \u11_mem[0] ;
 wire [31:0] \u11_mem[1] ;
 wire [31:0] \u11_mem[2] ;
 wire [31:0] \u11_mem[3] ;
 wire [2:0] u11_rp;
 wire [3:0] u11_wp;
 wire [1:0] u13_csr;
 wire [23:0] u13_icc_r;
 wire [28:0] u13_intm_r;
 wire [28:0] u13_ints_r;
 wire [31:0] u13_occ0_r;
 wire [15:0] u13_occ1_r;
 wire [19:0] u1_sr;
 wire [2:0] u26_cnt;
 wire [5:0] u26_ps_cnt;
 wire [7:0] u2_cnt;
 wire [3:0] u2_res_cnt;
 wire [5:0] u2_to_cnt;
 wire [31:0] \u3_mem[0] ;
 wire [31:0] \u3_mem[1] ;
 wire [31:0] \u3_mem[2] ;
 wire [31:0] \u3_mem[3] ;
 wire [3:0] u3_rp;
 wire [2:0] u3_wp;
 wire [31:0] \u4_mem[0] ;
 wire [31:0] \u4_mem[1] ;
 wire [31:0] \u4_mem[2] ;
 wire [31:0] \u4_mem[3] ;
 wire [3:0] u4_rp;
 wire [2:0] u4_wp;
 wire [31:0] \u5_mem[0] ;
 wire [31:0] \u5_mem[1] ;
 wire [31:0] \u5_mem[2] ;
 wire [31:0] \u5_mem[3] ;
 wire [3:0] u5_rp;
 wire [2:0] u5_wp;
 wire [31:0] \u6_mem[0] ;
 wire [31:0] \u6_mem[1] ;
 wire [31:0] \u6_mem[2] ;
 wire [31:0] \u6_mem[3] ;
 wire [3:0] u6_rp;
 wire [2:0] u6_wp;
 wire [31:0] \u7_mem[0] ;
 wire [31:0] \u7_mem[1] ;
 wire [31:0] \u7_mem[2] ;
 wire [31:0] \u7_mem[3] ;
 wire [3:0] u7_rp;
 wire [2:0] u7_wp;
 wire [31:0] \u8_mem[0] ;
 wire [31:0] \u8_mem[1] ;
 wire [31:0] \u8_mem[2] ;
 wire [31:0] \u8_mem[3] ;
 wire [3:0] u8_rp;
 wire [2:0] u8_wp;
 wire [15:0] u9_din_tmp1;
 wire [31:0] \u9_mem[0] ;
 wire [31:0] \u9_mem[1] ;
 wire [31:0] \u9_mem[2] ;
 wire [31:0] \u9_mem[3] ;
 wire [2:0] u9_rp;
 wire [3:0] u9_wp;
 wire [30:0] wb_din;

 HB1xp67_ASAP7_75t_R drc_buf_sp164977 (.A(n_5529),
    .Y(n_9294));
 HB1xp67_ASAP7_75t_R drc_buf_sp164978 (.A(n_5529),
    .Y(n_9295));
 HB1xp67_ASAP7_75t_R drc_buf_sp164979 (.A(n_5529),
    .Y(n_9296));
 HB1xp67_ASAP7_75t_R drc_buf_sp164980 (.A(n_5529),
    .Y(n_9297));
 HB1xp67_ASAP7_75t_R drc_buf_sp164981 (.A(n_5529),
    .Y(n_9298));
 HB1xp67_ASAP7_75t_R drc_buf_sp164982 (.A(n_5529),
    .Y(n_9299));
 HB1xp67_ASAP7_75t_R drc_buf_sp164983 (.A(n_5529),
    .Y(n_9300));
 HB1xp67_ASAP7_75t_R drc_buf_sp164984 (.A(n_5529),
    .Y(n_9301));
 HB1xp67_ASAP7_75t_R drc_buf_sp165026 (.A(ld),
    .Y(n_9344));
 HB1xp67_ASAP7_75t_R drc_buf_sp165027 (.A(ld),
    .Y(n_9345));
 HB1xp67_ASAP7_75t_R drc_buf_sp165028 (.A(ld),
    .Y(n_9346));
 HB1xp67_ASAP7_75t_R drc_buf_sp165029 (.A(ld),
    .Y(n_9347));
 HB1xp67_ASAP7_75t_R drc_buf_sp165030 (.A(ld),
    .Y(n_9348));
 HB1xp67_ASAP7_75t_R drc_buf_sp165031 (.A(ld),
    .Y(n_9349));
 HB1xp67_ASAP7_75t_R drc_buf_sp165032 (.A(ld),
    .Y(n_9350));
 HB1xp67_ASAP7_75t_R drc_buf_sp165033 (.A(ld),
    .Y(n_9351));
 HB1xp67_ASAP7_75t_R drc_buf_sp165077 (.A(n_9394),
    .Y(n_9396));
 HB1xp67_ASAP7_75t_R drc_buf_sp165078 (.A(n_9394),
    .Y(n_9397));
 HB1xp67_ASAP7_75t_R drc_buf_sp165079 (.A(n_9394),
    .Y(n_9398));
 HB1xp67_ASAP7_75t_R drc_buf_sp165082 (.A(n_9394),
    .Y(n_9395));
 HB1xp67_ASAP7_75t_R drc_buf_sp165083 (.A(ld),
    .Y(n_9394));
 HB1xp67_ASAP7_75t_R drc_buf_sp165146 (.A(n_5522),
    .Y(n_9466));
 HB1xp67_ASAP7_75t_R drc_buf_sp165147 (.A(n_5522),
    .Y(n_9467));
 HB1xp67_ASAP7_75t_R drc_buf_sp165148 (.A(n_5522),
    .Y(n_9468));
 HB1xp67_ASAP7_75t_R drc_buf_sp165270 (.A(n_5532),
    .Y(n_9629));
 HB1xp67_ASAP7_75t_R drc_buf_sp165271 (.A(n_5532),
    .Y(n_9630));
 INVx1_ASAP7_75t_L drc_buf_sp165370 (.A(n_66031),
    .Y(n_9735));
 INVx1_ASAP7_75t_SL drc_buf_sp165428 (.A(n_65968),
    .Y(n_9793));
 INVx1_ASAP7_75t_SL drc_buf_sp165457 (.A(n_65999),
    .Y(n_9822));
 INVx1_ASAP7_75t_SL drc_buf_sp165486 (.A(n_65962),
    .Y(n_9851));
 INVx1_ASAP7_75t_L drc_buf_sp165573 (.A(n_65993),
    .Y(n_9938));
 INVx2_ASAP7_75t_SL drc_buf_sp165576 (.A(n_9938),
    .Y(n_9942));
 INVx1_ASAP7_75t_SL drc_buf_sp165631 (.A(n_65965),
    .Y(n_9996));
 INVx2_ASAP7_75t_SL drc_buf_sp165634 (.A(n_9996),
    .Y(n_10000));
 INVx2_ASAP7_75t_SL drc_buf_sp165659 (.A(n_10025),
    .Y(n_10026));
 INVx1_ASAP7_75t_SL drc_buf_sp165660 (.A(n_65996),
    .Y(n_10025));
 INVx1_ASAP7_75t_L drc_buf_sp165689 (.A(n_65959),
    .Y(n_10054));
 INVx2_ASAP7_75t_SL drc_buf_sp165692 (.A(n_10054),
    .Y(n_10058));
 INVx1_ASAP7_75t_SL drc_buf_sp165718 (.A(n_65954),
    .Y(n_10083));
 INVx1_ASAP7_75t_SL drc_buf_sp165747 (.A(n_65948),
    .Y(n_10112));
 INVx1_ASAP7_75t_SL drc_buf_sp165775 (.A(n_65951),
    .Y(n_10140));
 INVx2_ASAP7_75t_SL drc_buf_sp165777 (.A(n_10140),
    .Y(n_10143));
 INVx2_ASAP7_75t_SL drc_buf_sp165826 (.A(n_10195),
    .Y(n_10196));
 INVx1_ASAP7_75t_SL drc_buf_sp165827 (.A(n_65932),
    .Y(n_10195));
 INVx2_ASAP7_75t_SL drc_buf_sp165829 (.A(n_10195),
    .Y(n_10198));
 INVx1_ASAP7_75t_SL drc_buf_sp165935 (.A(n_65929),
    .Y(n_10303));
 INVx2_ASAP7_75t_SL drc_buf_sp165962 (.A(n_65899),
    .Y(n_10330));
 INVx1_ASAP7_75t_SL drc_buf_sp165988 (.A(n_65919),
    .Y(n_10356));
 INVxp67_ASAP7_75t_SL drc_buf_sp166284 (.A(wb_din[29]),
    .Y(n_10661));
 HB1xp67_ASAP7_75t_R drc_buf_sp166329 (.A(out_le[4]),
    .Y(n_10709));
 HB1xp67_ASAP7_75t_R drc_buf_sp166354 (.A(out_le[3]),
    .Y(n_10735));
 HB1xp67_ASAP7_75t_R drc_buf_sp166379 (.A(n_5338),
    .Y(n_10761));
 HB1xp67_ASAP7_75t_R drc_buf_sp166404 (.A(n_5341),
    .Y(n_10787));
 HB1xp67_ASAP7_75t_R drc_buf_sp166429 (.A(n_5333),
    .Y(n_10813));
 HB1xp67_ASAP7_75t_R drc_buf_sp166454 (.A(out_le[5]),
    .Y(n_10839));
 HB1xp67_ASAP7_75t_R drc_buf_sp166649 (.A(out_le[2]),
    .Y(n_11046));
 INVx2_ASAP7_75t_SL drc_buf_sp170772 (.A(n_10661),
    .Y(n_15952));
 BUFx3_ASAP7_75t_SL drc_buf_sp213876 (.A(n_66842),
    .Y(n_66843));
 BUFx3_ASAP7_75t_SL drc_buf_sp213877 (.A(n_65965),
    .Y(n_66842));
 BUFx3_ASAP7_75t_SL drc_buf_sp213888 (.A(n_66855),
    .Y(n_66856));
 BUFx3_ASAP7_75t_SL drc_buf_sp213889 (.A(n_65962),
    .Y(n_66855));
 BUFx3_ASAP7_75t_SL drc_buf_sp213900 (.A(n_66868),
    .Y(n_66869));
 BUFx3_ASAP7_75t_SL drc_buf_sp213901 (.A(n_65959),
    .Y(n_66868));
 BUFx3_ASAP7_75t_SL drc_buf_sp213913 (.A(n_65993),
    .Y(n_66881));
 INVx5_ASAP7_75t_SL drc_buf_sp215496 (.A(n_9967),
    .Y(n_69010));
 BUFx3_ASAP7_75t_SL drc_buf_sp225155 (.A(n_79973),
    .Y(n_79971));
 BUFx3_ASAP7_75t_SL drc_buf_sp225156 (.A(n_79973),
    .Y(n_79972));
 HB1xp67_ASAP7_75t_SL drc_buf_sp225157 (.A(n_66881),
    .Y(n_79973));
 INVx2_ASAP7_75t_L drc_buf_sp40 (.A(n_10168),
    .Y(n_10171));
 INVx1_ASAP7_75t_SL drc_buf_sp41 (.A(n_65934),
    .Y(n_10168));
 INVx2_ASAP7_75t_L drc_buf_sp45 (.A(n_10890),
    .Y(n_10891));
 INVx1_ASAP7_75t_SL drc_buf_sp46 (.A(wb_din[1]),
    .Y(n_10890));
 INVx2_ASAP7_75t_L drc_buf_sp47 (.A(n_10637),
    .Y(n_10638));
 INVx2_ASAP7_75t_SL drc_buf_sp48 (.A(n_10637),
    .Y(n_10640));
 INVxp67_ASAP7_75t_SL drc_buf_sp49 (.A(wb_din[30]),
    .Y(n_10637));
 HB1xp67_ASAP7_75t_SL drc_bufs12 (.A(n_69010),
    .Y(n_69025));
 HB1xp67_ASAP7_75t_SL drc_bufs15 (.A(n_32582),
    .Y(n_32585));
 INVx1_ASAP7_75t_R drc_bufs164353 (.A(n_80),
    .Y(wb_ack_o));
 INVx1_ASAP7_75t_R drc_bufs164354 (.A(u12_wb_ack_o_745),
    .Y(n_80));
 HB1xp67_ASAP7_75t_SL drc_bufs164361 (.A(u26_ac97_rst_104),
    .Y(n_8351));
 HB1xp67_ASAP7_75t_SL drc_bufs164364 (.A(\u12_wb_data_o[29]_742 ),
    .Y(n_8354));
 HB1xp67_ASAP7_75t_SL drc_bufs164367 (.A(\u12_wb_data_o[30]_743 ),
    .Y(n_8357));
 HB1xp67_ASAP7_75t_SL drc_bufs164370 (.A(u13_int_1643),
    .Y(n_8360));
 HB1xp67_ASAP7_75t_SL drc_bufs164373 (.A(\u12_wb_data_o[16]_729 ),
    .Y(n_8363));
 HB1xp67_ASAP7_75t_SL drc_bufs164376 (.A(\u12_wb_data_o[20]_733 ),
    .Y(n_8366));
 HB1xp67_ASAP7_75t_SL drc_bufs164379 (.A(\u12_wb_data_o[21]_734 ),
    .Y(n_8369));
 HB1xp67_ASAP7_75t_SL drc_bufs164382 (.A(\u12_wb_data_o[22]_735 ),
    .Y(n_8372));
 HB1xp67_ASAP7_75t_SL drc_bufs164385 (.A(\u12_wb_data_o[25]_738 ),
    .Y(n_8375));
 HB1xp67_ASAP7_75t_SL drc_bufs164388 (.A(\u12_wb_data_o[27]_740 ),
    .Y(n_8378));
 INVxp67_ASAP7_75t_R drc_bufs164393 (.A(u16_u0_dma_req_52),
    .Y(n_46));
 INVxp67_ASAP7_75t_R drc_bufs164399 (.A(u16_u1_dma_req_52),
    .Y(n_131));
 INVxp67_ASAP7_75t_R drc_bufs164405 (.A(u16_u2_dma_req_52),
    .Y(n_33));
 INVxp67_ASAP7_75t_R drc_bufs164411 (.A(u16_u3_dma_req_52),
    .Y(n_25));
 INVxp67_ASAP7_75t_R drc_bufs164417 (.A(u16_u7_dma_req_52),
    .Y(n_15));
 INVxp67_ASAP7_75t_R drc_bufs164423 (.A(u16_u4_dma_req_52),
    .Y(n_83));
 INVxp67_ASAP7_75t_R drc_bufs164429 (.A(u16_u5_dma_req_52),
    .Y(n_119));
 INVxp67_ASAP7_75t_R drc_bufs164435 (.A(u16_u6_dma_req_52),
    .Y(n_86));
 INVxp67_ASAP7_75t_R drc_bufs164441 (.A(u16_u8_dma_req_52),
    .Y(n_108));
 HB1xp67_ASAP7_75t_SL drc_bufs164453 (.A(n_2467),
    .Y(n_8443));
 HB1xp67_ASAP7_75t_SL drc_bufs164456 (.A(u0_slt0_r[15]),
    .Y(n_8446));
 HB1xp67_ASAP7_75t_SL drc_bufs164459 (.A(\u12_wb_data_o[26]_739 ),
    .Y(n_8449));
 HB1xp67_ASAP7_75t_SL drc_bufs164462 (.A(\u12_wb_data_o[28]_741 ),
    .Y(n_8452));
 INVxp33_ASAP7_75t_R drc_bufs164466 (.A(n_31724),
    .Y(sync_pad_o));
 INVxp67_ASAP7_75t_R drc_bufs164469 (.A(n_8464),
    .Y(wb_data_o[17]));
 INVxp67_ASAP7_75t_R drc_bufs164470 (.A(\u12_wb_data_o[17]_730 ),
    .Y(n_8464));
 INVxp67_ASAP7_75t_R drc_bufs164472 (.A(n_8469),
    .Y(wb_data_o[19]));
 INVxp67_ASAP7_75t_R drc_bufs164473 (.A(\u12_wb_data_o[19]_732 ),
    .Y(n_8469));
 INVxp67_ASAP7_75t_R drc_bufs164475 (.A(n_8474),
    .Y(wb_data_o[5]));
 INVxp67_ASAP7_75t_R drc_bufs164476 (.A(\u12_wb_data_o[5]_718 ),
    .Y(n_8474));
 INVxp67_ASAP7_75t_R drc_bufs164478 (.A(n_8479),
    .Y(wb_data_o[31]));
 INVxp67_ASAP7_75t_R drc_bufs164479 (.A(\u12_wb_data_o[31]_744 ),
    .Y(n_8479));
 INVxp67_ASAP7_75t_R drc_bufs164481 (.A(n_8484),
    .Y(wb_data_o[1]));
 INVxp67_ASAP7_75t_R drc_bufs164482 (.A(\u12_wb_data_o[1]_714 ),
    .Y(n_8484));
 INVxp67_ASAP7_75t_R drc_bufs164484 (.A(n_8489),
    .Y(wb_data_o[2]));
 INVxp67_ASAP7_75t_R drc_bufs164485 (.A(\u12_wb_data_o[2]_715 ),
    .Y(n_8489));
 INVxp67_ASAP7_75t_R drc_bufs164487 (.A(n_8494),
    .Y(wb_data_o[14]));
 INVxp67_ASAP7_75t_R drc_bufs164488 (.A(\u12_wb_data_o[14]_727 ),
    .Y(n_8494));
 INVxp67_ASAP7_75t_R drc_bufs164490 (.A(n_8499),
    .Y(wb_data_o[8]));
 INVxp67_ASAP7_75t_R drc_bufs164491 (.A(\u12_wb_data_o[8]_721 ),
    .Y(n_8499));
 INVxp67_ASAP7_75t_R drc_bufs164493 (.A(n_8504),
    .Y(wb_data_o[6]));
 INVxp67_ASAP7_75t_R drc_bufs164494 (.A(\u12_wb_data_o[6]_719 ),
    .Y(n_8504));
 INVxp67_ASAP7_75t_R drc_bufs164496 (.A(n_8509),
    .Y(wb_data_o[18]));
 INVxp67_ASAP7_75t_R drc_bufs164497 (.A(\u12_wb_data_o[18]_731 ),
    .Y(n_8509));
 INVxp67_ASAP7_75t_R drc_bufs164499 (.A(n_8514),
    .Y(wb_data_o[10]));
 INVxp67_ASAP7_75t_R drc_bufs164500 (.A(\u12_wb_data_o[10]_723 ),
    .Y(n_8514));
 INVxp67_ASAP7_75t_R drc_bufs164502 (.A(n_8519),
    .Y(wb_data_o[0]));
 INVxp67_ASAP7_75t_R drc_bufs164503 (.A(\u12_wb_data_o[0]_713 ),
    .Y(n_8519));
 INVxp67_ASAP7_75t_R drc_bufs164505 (.A(n_8524),
    .Y(wb_data_o[12]));
 INVxp67_ASAP7_75t_R drc_bufs164506 (.A(\u12_wb_data_o[12]_725 ),
    .Y(n_8524));
 INVxp67_ASAP7_75t_R drc_bufs164508 (.A(n_8529),
    .Y(wb_data_o[13]));
 INVxp67_ASAP7_75t_R drc_bufs164509 (.A(\u12_wb_data_o[13]_726 ),
    .Y(n_8529));
 INVxp67_ASAP7_75t_R drc_bufs164511 (.A(n_8534),
    .Y(wb_data_o[15]));
 INVxp67_ASAP7_75t_R drc_bufs164512 (.A(\u12_wb_data_o[15]_728 ),
    .Y(n_8534));
 INVxp67_ASAP7_75t_R drc_bufs164514 (.A(n_8539),
    .Y(wb_data_o[11]));
 INVxp67_ASAP7_75t_R drc_bufs164515 (.A(\u12_wb_data_o[11]_724 ),
    .Y(n_8539));
 INVxp67_ASAP7_75t_R drc_bufs164517 (.A(n_8544),
    .Y(wb_data_o[23]));
 INVxp67_ASAP7_75t_R drc_bufs164518 (.A(\u12_wb_data_o[23]_736 ),
    .Y(n_8544));
 INVxp67_ASAP7_75t_R drc_bufs164520 (.A(n_8549),
    .Y(wb_data_o[7]));
 INVxp67_ASAP7_75t_R drc_bufs164521 (.A(\u12_wb_data_o[7]_720 ),
    .Y(n_8549));
 INVxp67_ASAP7_75t_R drc_bufs164523 (.A(n_8554),
    .Y(wb_data_o[4]));
 INVxp67_ASAP7_75t_R drc_bufs164524 (.A(\u12_wb_data_o[4]_717 ),
    .Y(n_8554));
 INVxp67_ASAP7_75t_R drc_bufs164526 (.A(n_8559),
    .Y(wb_data_o[24]));
 INVxp67_ASAP7_75t_R drc_bufs164527 (.A(\u12_wb_data_o[24]_737 ),
    .Y(n_8559));
 INVxp67_ASAP7_75t_R drc_bufs164529 (.A(n_8564),
    .Y(wb_data_o[3]));
 INVxp67_ASAP7_75t_R drc_bufs164530 (.A(\u12_wb_data_o[3]_716 ),
    .Y(n_8564));
 INVxp67_ASAP7_75t_R drc_bufs164532 (.A(n_8569),
    .Y(wb_data_o[9]));
 INVxp67_ASAP7_75t_R drc_bufs164533 (.A(\u12_wb_data_o[9]_722 ),
    .Y(n_8569));
 INVxp67_ASAP7_75t_R drc_bufs164535 (.A(n_8574),
    .Y(ac97_reset_pad_o_));
 INVxp67_ASAP7_75t_R drc_bufs164536 (.A(n_8351),
    .Y(n_8574));
 INVxp67_ASAP7_75t_R drc_bufs164538 (.A(n_8579),
    .Y(wb_data_o[30]));
 INVxp67_ASAP7_75t_R drc_bufs164539 (.A(n_8357),
    .Y(n_8579));
 INVxp67_ASAP7_75t_R drc_bufs164541 (.A(n_8584),
    .Y(wb_data_o[21]));
 INVxp67_ASAP7_75t_R drc_bufs164542 (.A(n_8369),
    .Y(n_8584));
 INVxp67_ASAP7_75t_R drc_bufs164544 (.A(n_8589),
    .Y(wb_data_o[22]));
 INVxp67_ASAP7_75t_R drc_bufs164545 (.A(n_8372),
    .Y(n_8589));
 INVxp67_ASAP7_75t_R drc_bufs164547 (.A(n_8594),
    .Y(int_o));
 INVxp67_ASAP7_75t_R drc_bufs164548 (.A(n_8360),
    .Y(n_8594));
 INVxp67_ASAP7_75t_R drc_bufs164550 (.A(n_8599),
    .Y(wb_data_o[25]));
 INVxp67_ASAP7_75t_R drc_bufs164551 (.A(n_8375),
    .Y(n_8599));
 INVxp67_ASAP7_75t_R drc_bufs164553 (.A(n_8604),
    .Y(wb_data_o[27]));
 INVxp67_ASAP7_75t_R drc_bufs164554 (.A(n_8378),
    .Y(n_8604));
 INVxp67_ASAP7_75t_R drc_bufs164556 (.A(n_8609),
    .Y(sdata_pad_o));
 INVxp67_ASAP7_75t_R drc_bufs164557 (.A(n_8446),
    .Y(n_8609));
 INVxp67_ASAP7_75t_R drc_bufs164559 (.A(n_8614),
    .Y(wb_data_o[29]));
 INVxp67_ASAP7_75t_R drc_bufs164560 (.A(n_8354),
    .Y(n_8614));
 INVxp67_ASAP7_75t_R drc_bufs164562 (.A(n_8619),
    .Y(wb_data_o[16]));
 INVxp67_ASAP7_75t_R drc_bufs164563 (.A(n_8363),
    .Y(n_8619));
 INVxp67_ASAP7_75t_R drc_bufs164565 (.A(n_8624),
    .Y(wb_data_o[20]));
 INVxp67_ASAP7_75t_R drc_bufs164566 (.A(n_8366),
    .Y(n_8624));
 INVxp33_ASAP7_75t_SL drc_bufs164571 (.A(n_8634),
    .Y(suspended_o));
 INVxp67_ASAP7_75t_R drc_bufs164572 (.A(n_8443),
    .Y(n_8634));
 INVxp33_ASAP7_75t_R drc_bufs164574 (.A(n_15),
    .Y(n_8638));
 INVxp33_ASAP7_75t_R drc_bufs164577 (.A(n_83),
    .Y(n_8643));
 INVxp33_ASAP7_75t_R drc_bufs164580 (.A(n_119),
    .Y(n_8648));
 INVxp33_ASAP7_75t_R drc_bufs164583 (.A(n_86),
    .Y(n_8653));
 INVxp33_ASAP7_75t_R drc_bufs164586 (.A(n_108),
    .Y(n_8658));
 INVxp67_ASAP7_75t_R drc_bufs164589 (.A(n_8664),
    .Y(wb_data_o[26]));
 INVxp67_ASAP7_75t_R drc_bufs164590 (.A(n_8449),
    .Y(n_8664));
 INVxp33_ASAP7_75t_R drc_bufs164592 (.A(n_46),
    .Y(n_8668));
 INVxp67_ASAP7_75t_R drc_bufs164595 (.A(n_8674),
    .Y(wb_data_o[28]));
 INVxp67_ASAP7_75t_R drc_bufs164596 (.A(n_8452),
    .Y(n_8674));
 INVxp33_ASAP7_75t_R drc_bufs164598 (.A(n_131),
    .Y(n_8678));
 INVxp33_ASAP7_75t_R drc_bufs164601 (.A(n_33),
    .Y(n_8683));
 INVxp33_ASAP7_75t_R drc_bufs164604 (.A(n_25),
    .Y(n_8688));
 INVxp33_ASAP7_75t_L drc_bufs189334 (.A(n_37601),
    .Y(dma_req_o[7]));
 INVxp67_ASAP7_75t_R drc_bufs189335 (.A(n_8638),
    .Y(n_37601));
 INVxp33_ASAP7_75t_L drc_bufs189336 (.A(n_37606),
    .Y(dma_req_o[4]));
 INVxp67_ASAP7_75t_R drc_bufs189337 (.A(n_8643),
    .Y(n_37606));
 INVxp33_ASAP7_75t_L drc_bufs189338 (.A(n_37611),
    .Y(dma_req_o[5]));
 INVxp67_ASAP7_75t_R drc_bufs189339 (.A(n_8648),
    .Y(n_37611));
 INVxp33_ASAP7_75t_L drc_bufs189340 (.A(n_37616),
    .Y(dma_req_o[0]));
 INVxp67_ASAP7_75t_R drc_bufs189341 (.A(n_8668),
    .Y(n_37616));
 INVxp33_ASAP7_75t_L drc_bufs189342 (.A(n_37621),
    .Y(dma_req_o[2]));
 INVxp67_ASAP7_75t_R drc_bufs189343 (.A(n_8683),
    .Y(n_37621));
 INVxp33_ASAP7_75t_L drc_bufs189344 (.A(n_37626),
    .Y(dma_req_o[1]));
 INVxp67_ASAP7_75t_R drc_bufs189345 (.A(n_8678),
    .Y(n_37626));
 INVxp33_ASAP7_75t_L drc_bufs190211 (.A(n_38792),
    .Y(dma_req_o[6]));
 INVxp67_ASAP7_75t_R drc_bufs190212 (.A(n_8653),
    .Y(n_38792));
 INVxp33_ASAP7_75t_L drc_bufs190213 (.A(n_38797),
    .Y(dma_req_o[8]));
 INVxp67_ASAP7_75t_R drc_bufs190214 (.A(n_8658),
    .Y(n_38797));
 INVxp33_ASAP7_75t_L drc_bufs190215 (.A(n_38802),
    .Y(dma_req_o[3]));
 INVxp67_ASAP7_75t_R drc_bufs190216 (.A(n_8688),
    .Y(n_38802));
 HB1xp67_ASAP7_75t_SL drc_bufs213859 (.A(n_66817),
    .Y(n_66824));
 HB1xp67_ASAP7_75t_R drc_bufs6 (.A(n_67246),
    .Y(n_66801));
 BUFx2_ASAP7_75t_R fopt (.A(n_5024),
    .Y(n_31863));
 INVx1_ASAP7_75t_SL fopt1 (.A(oc0_cfg[4]),
    .Y(n_18900));
 INVx1_ASAP7_75t_SL fopt1322 (.A(n_43090),
    .Y(n_7781));
 INVx1_ASAP7_75t_L fopt1377 (.A(n_7671),
    .Y(n_7672));
 INVx1_ASAP7_75t_SL fopt1378 (.A(oc2_cfg[3]),
    .Y(n_7671));
 BUFx2_ASAP7_75t_SL fopt1385 (.A(n_7668),
    .Y(n_698));
 INVx1_ASAP7_75t_SL fopt162394 (.A(n_1968),
    .Y(n_5674));
 INVx1_ASAP7_75t_SL fopt162402 (.A(n_5691),
    .Y(n_5687));
 INVx1_ASAP7_75t_SL fopt162413 (.A(n_41637),
    .Y(n_5706));
 HB1xp67_ASAP7_75t_SL fopt162431 (.A(n_26376),
    .Y(n_5741));
 BUFx3_ASAP7_75t_SL fopt162437 (.A(n_79019),
    .Y(n_5748));
 INVx2_ASAP7_75t_SL fopt162699 (.A(n_64993),
    .Y(n_6071));
 HB1xp67_ASAP7_75t_R fopt162739 (.A(n_18895),
    .Y(n_6115));
 INVxp67_ASAP7_75t_R fopt162752 (.A(n_12097),
    .Y(n_6136));
 HB1xp67_ASAP7_75t_SL fopt162754 (.A(n_21076),
    .Y(n_6138));
 INVx1_ASAP7_75t_SL fopt162757 (.A(oc3_cfg[3]),
    .Y(n_6141));
 INVx1_ASAP7_75t_R fopt162758 (.A(n_6146),
    .Y(n_6144));
 INVxp67_ASAP7_75t_SL fopt162760 (.A(n_64714),
    .Y(n_6146));
 HB1xp67_ASAP7_75t_R fopt162854 (.A(n_24588),
    .Y(n_6242));
 INVxp67_ASAP7_75t_SL fopt162859 (.A(u3_rp[2]),
    .Y(n_6248));
 INVx3_ASAP7_75t_SL fopt162860 (.A(u3_rp[2]),
    .Y(n_6249));
 INVxp67_ASAP7_75t_SL fopt163534 (.A(n_8212),
    .Y(n_6956));
 INVx2_ASAP7_75t_SL fopt163538 (.A(n_6960),
    .Y(n_6961));
 INVx1_ASAP7_75t_SL fopt163540 (.A(n_8212),
    .Y(n_6972));
 INVx11_ASAP7_75t_SL fopt163741_dup (.A(wb_addr_i[6]),
    .Y(n_6552));
 INVxp67_ASAP7_75t_SL fopt163801 (.A(n_1828),
    .Y(n_7319));
 INVx1_ASAP7_75t_SL fopt163956 (.A(n_17399),
    .Y(n_7582));
 INVx4_ASAP7_75t_SL fopt163967 (.A(u7_rp[2]),
    .Y(n_7653));
 INVx1_ASAP7_75t_SL fopt163968 (.A(u7_rp[2]),
    .Y(n_7656));
 INVx1_ASAP7_75t_SL fopt163976 (.A(oc2_cfg[3]),
    .Y(n_7667));
 BUFx2_ASAP7_75t_SL fopt163978 (.A(n_7671),
    .Y(n_2596));
 INVx2_ASAP7_75t_SL fopt164030 (.A(n_4339),
    .Y(n_7859));
 INVx1_ASAP7_75t_L fopt164034 (.A(n_19616),
    .Y(n_7863));
 INVx3_ASAP7_75t_SL fopt164037 (.A(u5_rp[1]),
    .Y(n_7869));
 BUFx3_ASAP7_75t_SL fopt164092 (.A(oc0_cfg[3]),
    .Y(n_573));
 INVxp67_ASAP7_75t_L fopt167964 (.A(n_31869),
    .Y(n_12519));
 INVx4_ASAP7_75t_SL fopt168634 (.A(n_2735),
    .Y(n_13295));
 INVx4_ASAP7_75t_SL fopt168635 (.A(n_27058),
    .Y(n_13304));
 INVx4_ASAP7_75t_SL fopt168636 (.A(n_27058),
    .Y(n_13312));
 INVx4_ASAP7_75t_SL fopt168641 (.A(n_2737),
    .Y(n_13325));
 INVx4_ASAP7_75t_SL fopt168642 (.A(n_2737),
    .Y(n_13333));
 HB1xp67_ASAP7_75t_R fopt168704 (.A(n_1661),
    .Y(n_13413));
 INVx4_ASAP7_75t_SL fopt168784 (.A(n_2836),
    .Y(n_13500));
 INVx4_ASAP7_75t_SL fopt168785 (.A(n_2836),
    .Y(n_13508));
 INVxp33_ASAP7_75t_SL fopt169158 (.A(n_36628),
    .Y(n_13978));
 INVxp67_ASAP7_75t_SL fopt169162 (.A(n_78273),
    .Y(n_13980));
 INVxp67_ASAP7_75t_SL fopt169190 (.A(n_14006),
    .Y(n_14009));
 INVx3_ASAP7_75t_SL fopt169192 (.A(u5_rp[2]),
    .Y(n_14010));
 INVx1_ASAP7_75t_SL fopt169193 (.A(n_26427),
    .Y(n_14012));
 INVx4_ASAP7_75t_SL fopt170775 (.A(n_2735),
    .Y(n_15954));
 INVx4_ASAP7_75t_SL fopt171563 (.A(n_2733),
    .Y(n_16900));
 INVx4_ASAP7_75t_SL fopt171564 (.A(n_2733),
    .Y(n_16908));
 INVxp67_ASAP7_75t_SL fopt172293 (.A(n_1828),
    .Y(n_17712));
 BUFx3_ASAP7_75t_SL fopt173083 (.A(n_78937),
    .Y(n_18739));
 HB1xp67_ASAP7_75t_SL fopt173087 (.A(n_77796),
    .Y(n_18743));
 INVx1_ASAP7_75t_SL fopt173234 (.A(n_18894),
    .Y(n_18895));
 INVx1_ASAP7_75t_L fopt173235 (.A(n_78938),
    .Y(n_18894));
 INVxp67_ASAP7_75t_R fopt173238 (.A(n_18894),
    .Y(n_18897));
 INVxp33_ASAP7_75t_R fopt173240 (.A(n_18900),
    .Y(n_18899));
 INVxp33_ASAP7_75t_R fopt173241 (.A(n_18903),
    .Y(n_18902));
 INVx1_ASAP7_75t_SL fopt173242 (.A(oc1_cfg[5]),
    .Y(n_18903));
 INVx2_ASAP7_75t_SL fopt173278 (.A(n_18964),
    .Y(n_18966));
 INVx2_ASAP7_75t_SL fopt173279 (.A(u6_wp[0]),
    .Y(n_18964));
 HB1xp67_ASAP7_75t_R fopt173311 (.A(u13_intm_r[1]),
    .Y(n_19002));
 INVx1_ASAP7_75t_SL fopt173318 (.A(n_19010),
    .Y(n_19009));
 BUFx3_ASAP7_75t_SL fopt173319 (.A(n_19013),
    .Y(n_19010));
 HB1xp67_ASAP7_75t_SL fopt173320 (.A(u26_ps_cnt[2]),
    .Y(n_19013));
 INVx1_ASAP7_75t_SL fopt173873 (.A(n_7869),
    .Y(n_19616));
 INVx3_ASAP7_75t_SL fopt174830 (.A(u6_wp[0]),
    .Y(n_20669));
 INVx1_ASAP7_75t_SL fopt174832 (.A(u6_wp[0]),
    .Y(n_20671));
 BUFx2_ASAP7_75t_SL fopt174833 (.A(n_20669),
    .Y(n_20673));
 INVx1_ASAP7_75t_SL fopt175575 (.A(n_4261),
    .Y(n_21507));
 INVx1_ASAP7_75t_SL fopt176458 (.A(n_7863),
    .Y(n_19593));
 BUFx6f_ASAP7_75t_SL fopt176651_dup (.A(n_32381),
    .Y(n_22780));
 INVx3_ASAP7_75t_SL fopt176671 (.A(n_78041),
    .Y(n_6122));
 INVx2_ASAP7_75t_SL fopt177154 (.A(u4_rp[2]),
    .Y(n_23524));
 BUFx3_ASAP7_75t_SL fopt177156 (.A(n_23524),
    .Y(n_23526));
 INVx2_ASAP7_75t_SL fopt178088 (.A(n_24587),
    .Y(n_24588));
 INVx1_ASAP7_75t_SL fopt178089 (.A(n_24586),
    .Y(n_24587));
 INVx1_ASAP7_75t_L fopt178090 (.A(u3_rp[2]),
    .Y(n_24586));
 HB1xp67_ASAP7_75t_R fopt178139 (.A(u13_intm_r[26]),
    .Y(n_24637));
 INVxp67_ASAP7_75t_SL fopt178188 (.A(n_24726),
    .Y(n_24725));
 HB1xp67_ASAP7_75t_SL fopt178189 (.A(u26_ps_cnt[3]),
    .Y(n_24726));
 INVx1_ASAP7_75t_L fopt178202 (.A(n_24742),
    .Y(n_24741));
 INVx1_ASAP7_75t_L fopt178203 (.A(n_24745),
    .Y(n_24742));
 INVx1_ASAP7_75t_SL fopt178204 (.A(u6_wp[1]),
    .Y(n_24745));
 BUFx3_ASAP7_75t_SL fopt178207 (.A(u6_wp[1]),
    .Y(n_24750));
 BUFx3_ASAP7_75t_L fopt178822 (.A(n_31844),
    .Y(n_25405));
 INVxp67_ASAP7_75t_SL fopt179708 (.A(n_26427),
    .Y(n_26428));
 HB1xp67_ASAP7_75t_SL fopt179709 (.A(n_14010),
    .Y(n_26427));
 INVxp67_ASAP7_75t_R fopt181935 (.A(n_28848),
    .Y(n_28850));
 INVx3_ASAP7_75t_SL fopt181975 (.A(n_176),
    .Y(n_425));
 BUFx6f_ASAP7_75t_SL fopt181996 (.A(n_65990),
    .Y(n_28913));
 BUFx6f_ASAP7_75t_SL fopt182304_dup188806 (.A(n_37387),
    .Y(n_36971));
 INVx3_ASAP7_75t_SL fopt182409 (.A(n_24750),
    .Y(n_29352));
 BUFx6f_ASAP7_75t_SL fopt182608 (.A(n_29619),
    .Y(n_29621));
 INVxp67_ASAP7_75t_SL fopt182915 (.A(n_51487),
    .Y(n_29953));
 INVx3_ASAP7_75t_SL fopt184226 (.A(n_26499),
    .Y(n_31460));
 INVx3_ASAP7_75t_SL fopt184227 (.A(n_26499),
    .Y(n_31464));
 INVxp67_ASAP7_75t_SL fopt184617 (.A(n_70241),
    .Y(n_31869));
 INVxp67_ASAP7_75t_SL fopt184619 (.A(n_31850),
    .Y(n_31872));
 BUFx6f_ASAP7_75t_SL fopt184937 (.A(n_32381),
    .Y(n_32382));
 BUFx3_ASAP7_75t_L fopt185166 (.A(n_66002),
    .Y(n_32644));
 BUFx2_ASAP7_75t_R fopt185167 (.A(n_66002),
    .Y(n_32650));
 BUFx3_ASAP7_75t_SL fopt185394 (.A(n_66015),
    .Y(n_32916));
 BUFx3_ASAP7_75t_SL fopt185483 (.A(n_66024),
    .Y(n_33024));
 BUFx3_ASAP7_75t_L fopt185622 (.A(n_75733),
    .Y(n_33203));
 INVx2_ASAP7_75t_SL fopt186117 (.A(u3_rp[2]),
    .Y(n_33784));
 BUFx2_ASAP7_75t_L fopt187722 (.A(out_slt0[7]),
    .Y(n_35645));
 BUFx6f_ASAP7_75t_SL fopt188056 (.A(valid_s),
    .Y(n_36068));
 INVx4_ASAP7_75t_SL fopt188067 (.A(n_62919),
    .Y(n_36078));
 INVx2_ASAP7_75t_SL fopt188071 (.A(n_62919),
    .Y(n_36082));
 INVxp67_ASAP7_75t_SL fopt188226 (.A(n_14054),
    .Y(n_36256));
 BUFx6f_ASAP7_75t_SL fopt188811 (.A(n_37387),
    .Y(n_36975));
 INVxp67_ASAP7_75t_SL fopt188959 (.A(n_1793),
    .Y(n_37142));
 INVx1_ASAP7_75t_SL fopt189096 (.A(oc3_cfg[3]),
    .Y(n_37335));
 INVx2_ASAP7_75t_SL fopt191528 (.A(n_40416),
    .Y(n_40417));
 INVx4_ASAP7_75t_SL fopt191529 (.A(u3_rp[1]),
    .Y(n_40416));
 INVxp67_ASAP7_75t_SL fopt191858 (.A(n_8306),
    .Y(n_40824));
 HB1xp67_ASAP7_75t_SL fopt192214 (.A(n_28952),
    .Y(n_41248));
 INVx1_ASAP7_75t_SL fopt192379 (.A(n_78276),
    .Y(n_41434));
 INVx4_ASAP7_75t_SL fopt193817 (.A(n_2734),
    .Y(n_43020));
 INVx4_ASAP7_75t_SL fopt193818 (.A(n_2734),
    .Y(n_43028));
 BUFx3_ASAP7_75t_SL fopt193864 (.A(n_43085),
    .Y(n_43088));
 HB1xp67_ASAP7_75t_SL fopt196699 (.A(n_46232),
    .Y(n_46233));
 BUFx6f_ASAP7_75t_SL fopt196702 (.A(n_46232),
    .Y(n_46234));
 INVx5_ASAP7_75t_SL fopt198341 (.A(n_48145),
    .Y(n_48146));
 INVx2_ASAP7_75t_SL fopt198349 (.A(n_48145),
    .Y(n_48153));
 BUFx6f_ASAP7_75t_SL fopt198736 (.A(n_48624),
    .Y(n_48625));
 BUFx3_ASAP7_75t_SL fopt198745 (.A(n_48624),
    .Y(n_48633));
 INVx5_ASAP7_75t_SL fopt198752 (.A(n_48625),
    .Y(n_48637));
 INVx2_ASAP7_75t_L fopt198759 (.A(n_48633),
    .Y(n_48648));
 INVxp67_ASAP7_75t_SL fopt2 (.A(n_36385),
    .Y(n_31886));
 INVx1_ASAP7_75t_SL fopt200058 (.A(o7_we),
    .Y(n_50109));
 INVx3_ASAP7_75t_SL fopt200240 (.A(n_7564),
    .Y(n_50342));
 INVx4_ASAP7_75t_SL fopt200277 (.A(n_7564),
    .Y(n_50388));
 INVx1_ASAP7_75t_SL fopt200350 (.A(n_64847),
    .Y(n_50463));
 INVxp67_ASAP7_75t_SL fopt200481 (.A(n_65030),
    .Y(n_50619));
 INVx1_ASAP7_75t_SL fopt200647 (.A(n_50810),
    .Y(n_5691));
 INVx2_ASAP7_75t_SL fopt200648 (.A(n_50809),
    .Y(n_50810));
 INVx2_ASAP7_75t_SL fopt200649 (.A(u4_rp[1]),
    .Y(n_50809));
 INVx4_ASAP7_75t_SL fopt200829 (.A(u7_rp[1]),
    .Y(n_51030));
 INVx4_ASAP7_75t_SL fopt201048 (.A(n_48436),
    .Y(n_51288));
 INVx4_ASAP7_75t_SL fopt201049 (.A(n_48436),
    .Y(n_51296));
 BUFx6f_ASAP7_75t_SL fopt202285 (.A(n_52892),
    .Y(n_52893));
 BUFx6f_ASAP7_75t_SL fopt202291 (.A(n_52892),
    .Y(n_52898));
 INVx1_ASAP7_75t_SL fopt202580 (.A(u8_rp[1]),
    .Y(n_53263));
 INVx3_ASAP7_75t_SL fopt202581 (.A(u8_rp[1]),
    .Y(n_53264));
 INVx3_ASAP7_75t_SL fopt205429 (.A(n_12219),
    .Y(n_56879));
 INVx3_ASAP7_75t_SL fopt205430 (.A(n_12219),
    .Y(n_56881));
 BUFx12f_ASAP7_75t_SL fopt212222 (.A(n_31888),
    .Y(n_64833));
 HB1xp67_ASAP7_75t_R fopt212236 (.A(n_14012),
    .Y(n_64848));
 INVx4_ASAP7_75t_SL fopt212376 (.A(n_2002),
    .Y(n_64993));
 INVx4_ASAP7_75t_SL fopt212592 (.A(n_65236),
    .Y(n_65239));
 INVx3_ASAP7_75t_SL fopt212932 (.A(n_7872),
    .Y(n_65642));
 INVxp33_ASAP7_75t_L fopt214309 (.A(n_67329),
    .Y(n_67328));
 INVx1_ASAP7_75t_SL fopt214310 (.A(u14_u5_en_out_l2),
    .Y(n_67329));
 BUFx3_ASAP7_75t_SL fopt218179 (.A(n_72057),
    .Y(n_72058));
 HB1xp67_ASAP7_75t_SL fopt223686 (.A(n_78932),
    .Y(n_78137));
 INVx2_ASAP7_75t_SL fopt224452 (.A(u8_rp[1]),
    .Y(n_78930));
 INVx2_ASAP7_75t_SL fopt224454 (.A(n_78930),
    .Y(n_78932));
 INVx4_ASAP7_75t_SL fopt224459 (.A(u6_rp[1]),
    .Y(n_78937));
 INVx4_ASAP7_75t_SL fopt224460 (.A(u6_rp[2]),
    .Y(n_78938));
 INVx2_ASAP7_75t_SL fopt2363 (.A(n_34541),
    .Y(n_5024));
 INVxp33_ASAP7_75t_R fopt3 (.A(n_65990),
    .Y(n_28926));
 INVxp33_ASAP7_75t_SL fopt60 (.A(n_7564),
    .Y(n_43394));
 INVx1_ASAP7_75t_SL fopt8 (.A(n_70322),
    .Y(n_5789));
 HB1xp67_ASAP7_75t_R g1 (.A(n_24736),
    .Y(n_21263));
 NOR2xp33_ASAP7_75t_SL g10 (.A(n_11011),
    .B(n_27061),
    .Y(n_13792));
 AND3x1_ASAP7_75t_R g100 (.A(n_12142),
    .B(n_48675),
    .C(n_75733),
    .Y(n_15495));
 OAI21xp33_ASAP7_75t_SL g102 (.A1(n_14914),
    .A2(n_15079),
    .B(n_43089),
    .Y(n_14917));
 AOI211x1_ASAP7_75t_SL g104 (.A1(n_7743),
    .A2(n_5028),
    .B(n_79202),
    .C(n_73306),
    .Y(n_7744));
 NAND3xp33_ASAP7_75t_SL g105 (.A(n_1433),
    .B(n_2254),
    .C(n_7514),
    .Y(n_7743));
 NAND2x1_ASAP7_75t_L g107 (.A(n_50456),
    .B(n_48639),
    .Y(n_12482));
 BUFx3_ASAP7_75t_SL g108 (.A(n_65954),
    .Y(n_65955));
 OAI211xp5_ASAP7_75t_SL g109 (.A1(n_59639),
    .A2(n_59640),
    .B(n_59641),
    .C(n_59642),
    .Y(n_59643));
 NOR2xp67_ASAP7_75t_SL g11 (.A(n_19615),
    .B(n_19593),
    .Y(n_19594));
 AOI221xp5_ASAP7_75t_SL g110 (.A1(n_8174),
    .A2(i4_dout[3]),
    .B1(i6_dout[3]),
    .B2(n_14933),
    .C(n_7087),
    .Y(n_16731));
 AOI21xp5_ASAP7_75t_SL g111 (.A1(n_2038),
    .A2(n_10626),
    .B(n_50289),
    .Y(n_16730));
 NAND2xp5_ASAP7_75t_SL g112 (.A(n_8341),
    .B(i3_dout[3]),
    .Y(n_16732));
 O2A1O1Ixp33_ASAP7_75t_R g113 (.A1(u8_wp[2]),
    .A2(n_2689),
    .B(n_463),
    .C(n_2743),
    .Y(n_43075));
 INVx2_ASAP7_75t_SL g114 (.A(n_37200),
    .Y(n_59639));
 INVxp33_ASAP7_75t_R g116 (.A(i3_dout[27]),
    .Y(n_65896));
 AOI22xp5_ASAP7_75t_SL g118 (.A1(n_24735),
    .A2(n_46558),
    .B1(\u9_mem[3] [2]),
    .B2(n_45330),
    .Y(n_46559));
 INVx1_ASAP7_75t_L g119 (.A(n_31058),
    .Y(n_17489));
 AND3x1_ASAP7_75t_SL g12 (.A(n_78094),
    .B(oc2_cfg[6]),
    .C(n_64296),
    .Y(n_64297));
 A2O1A1Ixp33_ASAP7_75t_SL g121 (.A1(n_47632),
    .A2(n_14966),
    .B(n_48223),
    .C(n_36363),
    .Y(n_14969));
 NAND2xp5_ASAP7_75t_SL g122 (.A(n_12097),
    .B(n_36525),
    .Y(n_14966));
 OAI222xp33_ASAP7_75t_SL g123 (.A1(n_14009),
    .A2(n_46227),
    .B1(n_2523),
    .B2(n_7571),
    .C1(n_2524),
    .C2(n_16672),
    .Y(n_7572));
 INVx1_ASAP7_75t_SL g124 (.A(n_7570),
    .Y(n_7571));
 NAND2xp5_ASAP7_75t_SL g125 (.A(n_1259),
    .B(n_6044),
    .Y(n_7570));
 AOI221xp5_ASAP7_75t_SL g126 (.A1(n_46644),
    .A2(n_25956),
    .B1(n_5062),
    .B2(out_slt7[14]),
    .C(n_4427),
    .Y(n_30357));
 AO21x1_ASAP7_75t_L g127 (.A1(u10_din_tmp1[11]),
    .A2(n_24336),
    .B(n_17609),
    .Y(n_61243));
 AND2x2_ASAP7_75t_L g128 (.A(out_slt4[14]),
    .B(n_43087),
    .Y(n_7586));
 AND2x2_ASAP7_75t_R g1282 (.A(out_slt4[11]),
    .B(n_7781),
    .Y(n_7788));
 O2A1O1Ixp33_ASAP7_75t_SL g1287 (.A1(n_35463),
    .A2(n_37051),
    .B(n_13825),
    .C(n_64852),
    .Y(n_7800));
 AOI21xp33_ASAP7_75t_SL g129 (.A1(n_2029),
    .A2(n_10626),
    .B(n_46110),
    .Y(n_46111));
 NAND2xp5_ASAP7_75t_SL g1292 (.A(n_20973),
    .B(n_1932),
    .Y(n_7806));
 NAND2x1p5_ASAP7_75t_SL g13 (.A(o6_we),
    .B(u5_wp[0]),
    .Y(n_24367));
 AOI221xp5_ASAP7_75t_SL g130 (.A1(n_14424),
    .A2(n_5091),
    .B1(n_4988),
    .B2(out_slt9[13]),
    .C(n_4356),
    .Y(n_14425));
 AOI21xp5_ASAP7_75t_SL g1300 (.A1(n_7766),
    .A2(n_35462),
    .B(n_26376),
    .Y(n_7803));
 AND2x2_ASAP7_75t_SL g1306 (.A(n_26379),
    .B(n_396),
    .Y(n_7772));
 NAND4xp25_ASAP7_75t_SL g131 (.A(n_1386),
    .B(n_2052),
    .C(n_2016),
    .D(n_1437),
    .Y(n_14424));
 NAND4xp25_ASAP7_75t_SL g132 (.A(n_2195),
    .B(n_2183),
    .C(n_1992),
    .D(n_1460),
    .Y(n_23393));
 AND2x4_ASAP7_75t_SL g1359 (.A(u5_rp[0]),
    .B(n_7667),
    .Y(n_7668));
 OAI211xp5_ASAP7_75t_SL g136 (.A1(n_46227),
    .A2(n_46228),
    .B(n_46229),
    .C(n_46230),
    .Y(n_46231));
 NOR2xp33_ASAP7_75t_SL g1360 (.A(n_65645),
    .B(n_29495),
    .Y(n_7689));
 AND2x2_ASAP7_75t_SL g1365 (.A(n_31907),
    .B(n_56864),
    .Y(n_7665));
 INVxp67_ASAP7_75t_L g1368 (.A(n_56864),
    .Y(n_7676));
 INVxp67_ASAP7_75t_L g1369 (.A(n_31907),
    .Y(n_7673));
 AOI211xp5_ASAP7_75t_SL g137 (.A1(n_7249),
    .A2(n_79104),
    .B(n_38377),
    .C(n_66671),
    .Y(n_7251));
 OAI211xp5_ASAP7_75t_SL g138 (.A1(n_2596),
    .A2(n_4320),
    .B(n_1457),
    .C(n_64998),
    .Y(n_7249));
 NAND2xp5_ASAP7_75t_SL g139 (.A(n_425),
    .B(n_48729),
    .Y(n_46230));
 AND2x2_ASAP7_75t_SL g14 (.A(u8_wp[0]),
    .B(o9_we),
    .Y(n_64191));
 AOI22xp5_ASAP7_75t_SL g140 (.A1(n_24735),
    .A2(n_15693),
    .B1(\u9_mem[3] [11]),
    .B2(n_45330),
    .Y(n_15694));
 NAND2x1_ASAP7_75t_SL g141 (.A(n_48643),
    .B(n_17594),
    .Y(n_15693));
 INVxp67_ASAP7_75t_L g143 (.A(n_10884),
    .Y(n_16726));
 NAND2xp5_ASAP7_75t_SL g144 (.A(n_65292),
    .B(n_78002),
    .Y(n_65293));
 AOI22xp5_ASAP7_75t_SL g145 (.A1(n_79178),
    .A2(\u8_mem[2] [6]),
    .B1(n_70885),
    .B2(\u8_mem[0] [6]),
    .Y(n_65292));
 NAND2x1_ASAP7_75t_SL g15 (.A(o9_we),
    .B(u8_wp[0]),
    .Y(n_64192));
 AOI22xp33_ASAP7_75t_R g152426__2398 (.A1(u0_slt0_r[14]),
    .A2(n_5522),
    .B1(n_9351),
    .B2(n_1913),
    .Y(n_5537));
 AOI22xp33_ASAP7_75t_R g152428__5107 (.A1(u0_slt0_r[13]),
    .A2(n_9630),
    .B1(out_slt0[14]),
    .B2(n_9344),
    .Y(n_5536));
 AOI22xp33_ASAP7_75t_R g152430__6260 (.A1(u0_slt0_r[12]),
    .A2(n_9296),
    .B1(out_slt0[13]),
    .B2(n_9395),
    .Y(n_5534));
 AOI22xp33_ASAP7_75t_R g152432__4319 (.A1(u0_slt0_r[11]),
    .A2(n_9629),
    .B1(n_1042),
    .B2(n_9394),
    .Y(n_5533));
 AOI22xp33_ASAP7_75t_R g152434__8428 (.A1(u0_slt0_r[10]),
    .A2(n_9295),
    .B1(n_517),
    .B2(n_9396),
    .Y(n_5530));
 NAND2xp33_ASAP7_75t_R g152436__5526 (.A(u0_slt0_r[9]),
    .B(n_9295),
    .Y(n_5528));
 AOI22xp33_ASAP7_75t_R g152438__6783 (.A1(u0_slt0_r[8]),
    .A2(n_9629),
    .B1(n_62918),
    .B2(n_9398),
    .Y(n_5527));
 AOI22xp33_ASAP7_75t_R g152440__3680 (.A1(u0_slt0_r[7]),
    .A2(n_9297),
    .B1(n_181),
    .B2(n_9398),
    .Y(n_5526));
 AOI22xp33_ASAP7_75t_R g152442__1617 (.A1(u0_slt0_r[6]),
    .A2(n_9298),
    .B1(n_35645),
    .B2(n_9397),
    .Y(n_5525));
 AOI22xp33_ASAP7_75t_R g152444__2802 (.A1(u0_slt0_r[5]),
    .A2(n_9630),
    .B1(n_37457),
    .B2(n_9396),
    .Y(n_5524));
 NAND2xp33_ASAP7_75t_R g152446__1705 (.A(u0_slt0_r[4]),
    .B(n_5522),
    .Y(n_5523));
 NAND2xp33_ASAP7_75t_R g152448__5122 (.A(u0_slt0_r[3]),
    .B(n_9629),
    .Y(n_5521));
 NAND2xp33_ASAP7_75t_R g152450__8246 (.A(u0_slt0_r[2]),
    .B(n_9300),
    .Y(n_5520));
 NAND2xp33_ASAP7_75t_R g152452__7098 (.A(u0_slt0_r[1]),
    .B(n_9299),
    .Y(n_5519));
 NAND2xp33_ASAP7_75t_R g152454__6131 (.A(u0_slt0_r[0]),
    .B(n_9298),
    .Y(n_5518));
 NAND2xp33_ASAP7_75t_R g152456__1881 (.A(u0_slt1_r[19]),
    .B(n_9467),
    .Y(n_5517));
 AOI22xp33_ASAP7_75t_R g152458__5115 (.A1(u0_slt1_r[18]),
    .A2(n_9468),
    .B1(crac_out[31]),
    .B2(n_9350),
    .Y(n_5516));
 AOI22xp33_ASAP7_75t_R g152460__7482 (.A1(u0_slt1_r[17]),
    .A2(n_9299),
    .B1(crac_out[22]),
    .B2(n_9349),
    .Y(n_5515));
 AOI22xp33_ASAP7_75t_R g152462__4733 (.A1(u0_slt1_r[16]),
    .A2(n_9629),
    .B1(crac_out[21]),
    .B2(n_9395),
    .Y(n_5514));
 AOI22xp33_ASAP7_75t_R g152464__6161 (.A1(u0_slt1_r[15]),
    .A2(n_9300),
    .B1(crac_out[20]),
    .B2(n_9394),
    .Y(n_5513));
 AOI22xp33_ASAP7_75t_R g152466__9315 (.A1(u0_slt1_r[14]),
    .A2(n_9301),
    .B1(crac_out[19]),
    .B2(n_9395),
    .Y(n_5512));
 AOI22xp33_ASAP7_75t_R g152468__9945 (.A1(u0_slt1_r[13]),
    .A2(n_9294),
    .B1(crac_out[18]),
    .B2(n_9348),
    .Y(n_5511));
 AOI22xp33_ASAP7_75t_R g152470__2883 (.A1(u0_slt1_r[12]),
    .A2(n_9295),
    .B1(crac_out[17]),
    .B2(n_9347),
    .Y(n_5510));
 AOI22xp33_ASAP7_75t_R g152472__2346 (.A1(u0_slt1_r[11]),
    .A2(n_9630),
    .B1(crac_out[16]),
    .B2(n_9346),
    .Y(n_5509));
 NAND2xp33_ASAP7_75t_R g152474__1666 (.A(u0_slt1_r[10]),
    .B(n_9300),
    .Y(n_5508));
 NAND2xp33_ASAP7_75t_R g152476__7410 (.A(u0_slt1_r[9]),
    .B(n_9299),
    .Y(n_5507));
 NAND2xp33_ASAP7_75t_R g152478__6417 (.A(u0_slt1_r[8]),
    .B(n_9298),
    .Y(n_5506));
 NAND2xp33_ASAP7_75t_R g152480__5477 (.A(u0_slt1_r[7]),
    .B(n_9629),
    .Y(n_5505));
 NAND2xp33_ASAP7_75t_R g152482__2398 (.A(u0_slt1_r[6]),
    .B(n_9297),
    .Y(n_5504));
 NAND2xp33_ASAP7_75t_R g152484__5107 (.A(u0_slt1_r[5]),
    .B(n_9296),
    .Y(n_5503));
 NAND2xp33_ASAP7_75t_R g152486__6260 (.A(u0_slt1_r[4]),
    .B(n_9301),
    .Y(n_5502));
 NAND2xp33_ASAP7_75t_R g152488__4319 (.A(u0_slt1_r[3]),
    .B(n_9300),
    .Y(n_5501));
 NAND2xp33_ASAP7_75t_R g152490__8428 (.A(u0_slt1_r[2]),
    .B(n_5522),
    .Y(n_5500));
 NAND2xp33_ASAP7_75t_R g152492__5526 (.A(u0_slt1_r[1]),
    .B(n_9299),
    .Y(n_5499));
 NAND2xp33_ASAP7_75t_R g152494__6783 (.A(u0_slt1_r[0]),
    .B(n_9298),
    .Y(n_5498));
 NAND2xp33_ASAP7_75t_R g152496__3680 (.A(u0_slt2_r[19]),
    .B(n_9297),
    .Y(n_5497));
 AOI22xp33_ASAP7_75t_R g152498__1617 (.A1(u0_slt2_r[18]),
    .A2(n_9296),
    .B1(crac_out[15]),
    .B2(n_9396),
    .Y(n_5496));
 AOI22xp33_ASAP7_75t_R g152500__2802 (.A1(u0_slt2_r[17]),
    .A2(n_9299),
    .B1(crac_out[14]),
    .B2(n_9345),
    .Y(n_5495));
 AOI22xp33_ASAP7_75t_R g152502__1705 (.A1(u0_slt2_r[16]),
    .A2(n_9295),
    .B1(crac_out[13]),
    .B2(n_9344),
    .Y(n_5494));
 AOI22xp33_ASAP7_75t_R g152504__5122 (.A1(u0_slt2_r[15]),
    .A2(n_9294),
    .B1(crac_out[12]),
    .B2(n_9398),
    .Y(n_5493));
 AOI22xp33_ASAP7_75t_R g152506__8246 (.A1(u0_slt2_r[14]),
    .A2(n_9301),
    .B1(crac_out[11]),
    .B2(n_9351),
    .Y(n_5492));
 AOI22xp33_ASAP7_75t_R g152508__7098 (.A1(u0_slt2_r[13]),
    .A2(n_9300),
    .B1(crac_out[10]),
    .B2(n_9350),
    .Y(n_5491));
 AOI22xp33_ASAP7_75t_R g152510__6131 (.A1(u0_slt2_r[12]),
    .A2(n_9299),
    .B1(crac_out[9]),
    .B2(n_9398),
    .Y(n_5490));
 AOI22xp33_ASAP7_75t_R g152512__1881 (.A1(u0_slt2_r[11]),
    .A2(n_9298),
    .B1(crac_out[8]),
    .B2(n_9349),
    .Y(n_5489));
 AOI22xp33_ASAP7_75t_R g152514__5115 (.A1(u0_slt2_r[10]),
    .A2(n_9297),
    .B1(crac_out[7]),
    .B2(n_9348),
    .Y(n_5488));
 AOI22xp33_ASAP7_75t_R g152516__7482 (.A1(u0_slt2_r[9]),
    .A2(n_9296),
    .B1(crac_out[6]),
    .B2(n_9397),
    .Y(n_5487));
 AOI22xp33_ASAP7_75t_R g152518__4733 (.A1(u0_slt2_r[8]),
    .A2(n_9467),
    .B1(crac_out[5]),
    .B2(n_9347),
    .Y(n_5486));
 AOI22xp33_ASAP7_75t_R g152520__6161 (.A1(u0_slt2_r[7]),
    .A2(n_9295),
    .B1(crac_out[4]),
    .B2(n_9346),
    .Y(n_5485));
 AOI22xp33_ASAP7_75t_R g152522__9315 (.A1(u0_slt2_r[6]),
    .A2(n_9294),
    .B1(crac_out[3]),
    .B2(n_9345),
    .Y(n_5484));
 AOI22xp33_ASAP7_75t_R g152524__9945 (.A1(u0_slt2_r[5]),
    .A2(n_9629),
    .B1(crac_out[2]),
    .B2(n_9344),
    .Y(n_5483));
 AOI22xp33_ASAP7_75t_R g152526__2883 (.A1(u0_slt2_r[4]),
    .A2(n_9301),
    .B1(crac_out[1]),
    .B2(n_9351),
    .Y(n_5482));
 AOI22xp33_ASAP7_75t_R g152528__2346 (.A1(u0_slt2_r[3]),
    .A2(n_9300),
    .B1(crac_out[0]),
    .B2(n_9396),
    .Y(n_5481));
 NAND2xp33_ASAP7_75t_R g152530__1666 (.A(u0_slt2_r[2]),
    .B(n_9467),
    .Y(n_5480));
 NAND2xp33_ASAP7_75t_R g152532__7410 (.A(u0_slt2_r[1]),
    .B(n_9294),
    .Y(n_5479));
 NAND2xp33_ASAP7_75t_R g152534__6417 (.A(u0_slt2_r[0]),
    .B(n_9466),
    .Y(n_5478));
 NAND2xp33_ASAP7_75t_R g152536__5477 (.A(u0_slt3_r[19]),
    .B(n_9468),
    .Y(n_5477));
 AOI22xp33_ASAP7_75t_R g152538__2398 (.A1(u0_slt3_r[18]),
    .A2(n_9466),
    .B1(out_slt3[19]),
    .B2(n_9395),
    .Y(n_5476));
 AOI22xp33_ASAP7_75t_R g152540__5107 (.A1(u0_slt3_r[17]),
    .A2(n_9298),
    .B1(out_slt3[18]),
    .B2(n_9394),
    .Y(n_5475));
 AOI22xp33_ASAP7_75t_R g152542__6260 (.A1(u0_slt3_r[16]),
    .A2(n_9297),
    .B1(out_slt3[17]),
    .B2(n_9395),
    .Y(n_5474));
 AOI22xp33_ASAP7_75t_R g152544__4319 (.A1(u0_slt3_r[15]),
    .A2(n_9296),
    .B1(out_slt3[16]),
    .B2(n_9350),
    .Y(n_5473));
 AOI22xp33_ASAP7_75t_R g152546__8428 (.A1(u0_slt3_r[14]),
    .A2(n_9295),
    .B1(out_slt3[15]),
    .B2(n_9349),
    .Y(n_5472));
 AOI22xp33_ASAP7_75t_R g152548__5526 (.A1(u0_slt3_r[13]),
    .A2(n_9294),
    .B1(out_slt3[14]),
    .B2(n_9348),
    .Y(n_5471));
 AOI22xp33_ASAP7_75t_R g152550__6783 (.A1(u0_slt3_r[12]),
    .A2(n_5522),
    .B1(out_slt3[13]),
    .B2(n_9347),
    .Y(n_5470));
 AOI22xp33_ASAP7_75t_R g152552__3680 (.A1(u0_slt3_r[11]),
    .A2(n_9630),
    .B1(out_slt3[12]),
    .B2(n_9346),
    .Y(n_5469));
 AOI22xp33_ASAP7_75t_R g152554__1617 (.A1(u0_slt3_r[10]),
    .A2(n_9629),
    .B1(out_slt3[11]),
    .B2(n_9345),
    .Y(n_5468));
 AOI22xp33_ASAP7_75t_R g152556__2802 (.A1(u0_slt3_r[9]),
    .A2(n_9301),
    .B1(out_slt3[10]),
    .B2(n_9344),
    .Y(n_5467));
 AOI22xp33_ASAP7_75t_R g152558__1705 (.A1(u0_slt3_r[8]),
    .A2(n_9300),
    .B1(out_slt3[9]),
    .B2(n_9351),
    .Y(n_5466));
 AOI22xp33_ASAP7_75t_R g152560__5122 (.A1(u0_slt3_r[7]),
    .A2(n_9299),
    .B1(out_slt3[8]),
    .B2(n_9350),
    .Y(n_5465));
 AOI22xp33_ASAP7_75t_R g152562__8246 (.A1(u0_slt3_r[6]),
    .A2(n_9298),
    .B1(out_slt3[7]),
    .B2(n_9349),
    .Y(n_5464));
 AOI22xp33_ASAP7_75t_R g152564__7098 (.A1(u0_slt3_r[5]),
    .A2(n_9468),
    .B1(out_slt3[6]),
    .B2(n_9348),
    .Y(n_5463));
 AOI22xp33_ASAP7_75t_R g152566__6131 (.A1(u0_slt3_r[4]),
    .A2(n_9297),
    .B1(out_slt3[5]),
    .B2(n_9347),
    .Y(n_5462));
 AOI22xp33_ASAP7_75t_R g152568__1881 (.A1(u0_slt3_r[3]),
    .A2(n_9296),
    .B1(out_slt3[4]),
    .B2(n_9346),
    .Y(n_5461));
 AOI22xp33_ASAP7_75t_R g152570__5115 (.A1(u0_slt3_r[2]),
    .A2(n_9295),
    .B1(out_slt3[3]),
    .B2(n_9345),
    .Y(n_5460));
 AOI22xp33_ASAP7_75t_R g152572__7482 (.A1(u0_slt3_r[1]),
    .A2(n_9294),
    .B1(out_slt3[2]),
    .B2(n_9344),
    .Y(n_5459));
 AOI22xp33_ASAP7_75t_R g152574__4733 (.A1(u0_slt3_r[0]),
    .A2(n_9467),
    .B1(out_slt3[1]),
    .B2(n_9396),
    .Y(n_5458));
 AOI22xp33_ASAP7_75t_R g152576__6161 (.A1(u0_slt4_r[19]),
    .A2(n_9466),
    .B1(out_slt3[0]),
    .B2(n_9351),
    .Y(n_5457));
 AOI22xp33_ASAP7_75t_R g152578__9315 (.A1(u0_slt4_r[18]),
    .A2(n_9301),
    .B1(out_slt4[19]),
    .B2(n_9350),
    .Y(n_5456));
 AOI22xp33_ASAP7_75t_R g152580__9945 (.A1(u0_slt4_r[17]),
    .A2(n_9300),
    .B1(out_slt4[18]),
    .B2(n_9349),
    .Y(n_5455));
 AOI22xp33_ASAP7_75t_R g152582__2883 (.A1(u0_slt4_r[16]),
    .A2(n_9299),
    .B1(out_slt4[17]),
    .B2(n_9348),
    .Y(n_5454));
 AOI22xp33_ASAP7_75t_R g152584__2346 (.A1(u0_slt4_r[15]),
    .A2(n_9298),
    .B1(out_slt4[16]),
    .B2(n_9347),
    .Y(n_5453));
 AOI22xp33_ASAP7_75t_R g152586__1666 (.A1(u0_slt4_r[14]),
    .A2(n_9630),
    .B1(out_slt4[15]),
    .B2(n_9346),
    .Y(n_5452));
 AOI22xp33_ASAP7_75t_R g152588__7410 (.A1(u0_slt4_r[13]),
    .A2(n_9629),
    .B1(out_slt4[14]),
    .B2(n_9345),
    .Y(n_5451));
 AOI22xp33_ASAP7_75t_R g152590__6417 (.A1(u0_slt4_r[12]),
    .A2(n_9297),
    .B1(out_slt4[13]),
    .B2(n_9344),
    .Y(n_5450));
 AOI22xp33_ASAP7_75t_R g152592__5477 (.A1(u0_slt4_r[11]),
    .A2(n_9296),
    .B1(out_slt4[12]),
    .B2(n_9351),
    .Y(n_5449));
 AOI22xp33_ASAP7_75t_R g152594__2398 (.A1(u0_slt4_r[10]),
    .A2(n_9630),
    .B1(out_slt4[11]),
    .B2(n_9398),
    .Y(n_5448));
 AOI22xp33_ASAP7_75t_R g152596__5107 (.A1(u0_slt4_r[9]),
    .A2(n_9295),
    .B1(out_slt4[10]),
    .B2(n_9398),
    .Y(n_5447));
 AOI22xp33_ASAP7_75t_R g152598__6260 (.A1(u0_slt4_r[8]),
    .A2(n_9294),
    .B1(out_slt4[9]),
    .B2(n_9397),
    .Y(n_5446));
 AOI22xp33_ASAP7_75t_R g152600__4319 (.A1(u0_slt4_r[7]),
    .A2(n_9301),
    .B1(out_slt4[8]),
    .B2(n_9396),
    .Y(n_5445));
 AOI22xp33_ASAP7_75t_R g152602__8428 (.A1(u0_slt4_r[6]),
    .A2(n_5522),
    .B1(out_slt4[7]),
    .B2(n_9395),
    .Y(n_5444));
 AOI22xp33_ASAP7_75t_R g152604__5526 (.A1(u0_slt4_r[5]),
    .A2(n_9300),
    .B1(out_slt4[6]),
    .B2(n_9394),
    .Y(n_5443));
 AOI22xp33_ASAP7_75t_R g152606__6783 (.A1(u0_slt4_r[4]),
    .A2(n_9468),
    .B1(out_slt4[5]),
    .B2(n_9350),
    .Y(n_5442));
 AOI22xp33_ASAP7_75t_R g152608__3680 (.A1(u0_slt4_r[3]),
    .A2(n_9294),
    .B1(out_slt4[4]),
    .B2(n_9395),
    .Y(n_5441));
 AOI22xp33_ASAP7_75t_R g152610__1617 (.A1(u0_slt4_r[2]),
    .A2(n_9298),
    .B1(out_slt4[3]),
    .B2(n_9396),
    .Y(n_5440));
 AOI22xp33_ASAP7_75t_R g152612__2802 (.A1(u0_slt4_r[1]),
    .A2(n_9467),
    .B1(out_slt4[2]),
    .B2(n_9398),
    .Y(n_5439));
 AOI22xp33_ASAP7_75t_R g152614__1705 (.A1(u0_slt4_r[0]),
    .A2(n_9297),
    .B1(out_slt4[1]),
    .B2(n_9398),
    .Y(n_5438));
 AOI22xp33_ASAP7_75t_R g152616__5122 (.A1(u0_slt5_r[19]),
    .A2(n_9629),
    .B1(out_slt4[0]),
    .B2(n_9349),
    .Y(n_5437));
 NAND2xp33_ASAP7_75t_R g152618__8246 (.A(u0_slt5_r[18]),
    .B(n_9630),
    .Y(n_5436));
 NAND2xp33_ASAP7_75t_R g152620__7098 (.A(u0_slt5_r[17]),
    .B(n_9466),
    .Y(n_5435));
 NAND2xp33_ASAP7_75t_R g152622__6131 (.A(u0_slt5_r[16]),
    .B(n_9468),
    .Y(n_5434));
 NAND2xp33_ASAP7_75t_R g152624__1881 (.A(u0_slt5_r[15]),
    .B(n_9630),
    .Y(n_5433));
 NAND2xp33_ASAP7_75t_R g152626__5115 (.A(u0_slt5_r[14]),
    .B(n_9630),
    .Y(n_5432));
 NAND2xp33_ASAP7_75t_R g152628__7482 (.A(u0_slt5_r[13]),
    .B(n_9301),
    .Y(n_5431));
 NAND2xp33_ASAP7_75t_R g152630__4733 (.A(u0_slt5_r[12]),
    .B(n_9467),
    .Y(n_5430));
 NAND2xp33_ASAP7_75t_R g152632__6161 (.A(u0_slt5_r[11]),
    .B(n_9466),
    .Y(n_5429));
 NAND2xp33_ASAP7_75t_R g152634__9315 (.A(u0_slt5_r[10]),
    .B(n_9630),
    .Y(n_5428));
 NAND2xp33_ASAP7_75t_R g152636__9945 (.A(u0_slt5_r[9]),
    .B(n_9629),
    .Y(n_5427));
 NAND2xp33_ASAP7_75t_R g152638__2883 (.A(u0_slt5_r[8]),
    .B(n_9468),
    .Y(n_5426));
 NAND2xp33_ASAP7_75t_R g152640__2346 (.A(u0_slt5_r[7]),
    .B(n_9296),
    .Y(n_5425));
 NAND2xp33_ASAP7_75t_R g152642__1666 (.A(u0_slt5_r[6]),
    .B(n_9295),
    .Y(n_5424));
 NAND2xp33_ASAP7_75t_R g152644__7410 (.A(u0_slt5_r[5]),
    .B(n_9296),
    .Y(n_5423));
 NAND2xp33_ASAP7_75t_R g152646__6417 (.A(u0_slt5_r[4]),
    .B(n_9297),
    .Y(n_5422));
 NAND2xp33_ASAP7_75t_R g152648__5477 (.A(u0_slt5_r[3]),
    .B(n_9301),
    .Y(n_5421));
 NAND2xp33_ASAP7_75t_R g152650__2398 (.A(u0_slt5_r[2]),
    .B(n_9294),
    .Y(n_5420));
 NAND2xp33_ASAP7_75t_R g152652__5107 (.A(u0_slt5_r[1]),
    .B(n_9296),
    .Y(n_5419));
 NAND2xp33_ASAP7_75t_R g152654__6260 (.A(u0_slt5_r[0]),
    .B(n_9297),
    .Y(n_5418));
 NAND2xp33_ASAP7_75t_R g152656__4319 (.A(u0_slt6_r[19]),
    .B(n_9298),
    .Y(n_5417));
 AOI22xp33_ASAP7_75t_R g152658__8428 (.A1(u0_slt6_r[18]),
    .A2(n_9294),
    .B1(out_slt6[19]),
    .B2(n_9344),
    .Y(n_5416));
 AOI22xp33_ASAP7_75t_R g152660__5526 (.A1(u0_slt6_r[17]),
    .A2(n_9301),
    .B1(out_slt6[18]),
    .B2(n_9397),
    .Y(n_5415));
 AOI22xp33_ASAP7_75t_R g152662__6783 (.A1(u0_slt6_r[16]),
    .A2(n_9300),
    .B1(out_slt6[17]),
    .B2(n_9396),
    .Y(n_5414));
 AOI22xp33_ASAP7_75t_R g152664__3680 (.A1(u0_slt6_r[15]),
    .A2(n_5522),
    .B1(out_slt6[16]),
    .B2(n_9347),
    .Y(n_5413));
 AOI22xp33_ASAP7_75t_R g152666__1617 (.A1(u0_slt6_r[14]),
    .A2(n_9468),
    .B1(out_slt6[15]),
    .B2(n_9346),
    .Y(n_5412));
 AOI22xp33_ASAP7_75t_R g152668__2802 (.A1(u0_slt6_r[13]),
    .A2(n_9299),
    .B1(out_slt6[14]),
    .B2(n_9395),
    .Y(n_5411));
 AOI22xp33_ASAP7_75t_R g152670__1705 (.A1(u0_slt6_r[12]),
    .A2(n_9298),
    .B1(out_slt6[13]),
    .B2(n_9394),
    .Y(n_5410));
 AOI22xp33_ASAP7_75t_R g152672__5122 (.A1(u0_slt6_r[11]),
    .A2(n_9297),
    .B1(out_slt6[12]),
    .B2(n_9395),
    .Y(n_5409));
 AOI22xp33_ASAP7_75t_R g152674__8246 (.A1(u0_slt6_r[10]),
    .A2(n_9296),
    .B1(out_slt6[11]),
    .B2(n_9345),
    .Y(n_5408));
 AOI22xp33_ASAP7_75t_R g152676__7098 (.A1(u0_slt6_r[9]),
    .A2(n_9295),
    .B1(out_slt6[10]),
    .B2(n_9396),
    .Y(n_5407));
 AOI22xp33_ASAP7_75t_R g152678__6131 (.A1(u0_slt6_r[8]),
    .A2(n_9294),
    .B1(out_slt6[9]),
    .B2(n_9344),
    .Y(n_5406));
 AOI22xp33_ASAP7_75t_R g152680__1881 (.A1(u0_slt6_r[7]),
    .A2(n_9301),
    .B1(out_slt6[8]),
    .B2(n_9351),
    .Y(n_5405));
 AOI22xp33_ASAP7_75t_R g152682__5115 (.A1(u0_slt6_r[6]),
    .A2(n_5522),
    .B1(out_slt6[7]),
    .B2(n_9398),
    .Y(n_5404));
 AOI22xp33_ASAP7_75t_R g152684__7482 (.A1(u0_slt6_r[5]),
    .A2(n_9300),
    .B1(out_slt6[6]),
    .B2(n_9398),
    .Y(n_5403));
 AOI22xp33_ASAP7_75t_R g152686__4733 (.A1(u0_slt6_r[4]),
    .A2(n_9466),
    .B1(out_slt6[5]),
    .B2(n_9350),
    .Y(n_5402));
 AOI22xp33_ASAP7_75t_R g152688__6161 (.A1(u0_slt6_r[3]),
    .A2(n_5522),
    .B1(out_slt6[4]),
    .B2(n_9397),
    .Y(n_5401));
 AOI22xp33_ASAP7_75t_R g152690__9315 (.A1(u0_slt6_r[2]),
    .A2(n_9468),
    .B1(out_slt6[3]),
    .B2(n_9396),
    .Y(n_5400));
 AOI22xp33_ASAP7_75t_R g152692__9945 (.A1(u0_slt6_r[1]),
    .A2(n_9299),
    .B1(out_slt6[2]),
    .B2(n_9349),
    .Y(n_5399));
 AOI22xp33_ASAP7_75t_R g152694__2883 (.A1(u0_slt6_r[0]),
    .A2(n_9467),
    .B1(out_slt6[1]),
    .B2(n_9348),
    .Y(n_5398));
 AOI22xp33_ASAP7_75t_R g152696__2346 (.A1(u0_slt7_r[19]),
    .A2(n_9466),
    .B1(out_slt6[0]),
    .B2(n_9395),
    .Y(n_5397));
 AOI22xp33_ASAP7_75t_R g152698__1666 (.A1(u0_slt7_r[18]),
    .A2(n_5522),
    .B1(out_slt7[19]),
    .B2(n_9394),
    .Y(n_5396));
 AOI22xp33_ASAP7_75t_R g152700__7410 (.A1(u0_slt7_r[17]),
    .A2(n_9298),
    .B1(out_slt7[18]),
    .B2(n_9347),
    .Y(n_5395));
 AOI22xp33_ASAP7_75t_R g152702__6417 (.A1(u0_slt7_r[16]),
    .A2(n_9468),
    .B1(out_slt7[17]),
    .B2(n_9346),
    .Y(n_5394));
 AOI22xp33_ASAP7_75t_R g152704__5477 (.A1(u0_slt7_r[15]),
    .A2(n_9467),
    .B1(out_slt7[16]),
    .B2(n_9345),
    .Y(n_5393));
 AOI22xp33_ASAP7_75t_R g152706__2398 (.A1(u0_slt7_r[14]),
    .A2(n_9297),
    .B1(out_slt7[15]),
    .B2(n_9395),
    .Y(n_5392));
 AOI22xp33_ASAP7_75t_R g152708__5107 (.A1(u0_slt7_r[13]),
    .A2(n_9466),
    .B1(out_slt7[14]),
    .B2(n_9344),
    .Y(n_5391));
 AOI22xp33_ASAP7_75t_R g152710__6260 (.A1(u0_slt7_r[12]),
    .A2(n_9296),
    .B1(out_slt7[13]),
    .B2(n_9351),
    .Y(n_5390));
 AOI22xp33_ASAP7_75t_R g152712__4319 (.A1(u0_slt7_r[11]),
    .A2(n_9295),
    .B1(out_slt7[12]),
    .B2(n_9350),
    .Y(n_5389));
 AOI22xp33_ASAP7_75t_R g152714__8428 (.A1(u0_slt7_r[10]),
    .A2(n_9294),
    .B1(out_slt7[11]),
    .B2(n_9349),
    .Y(n_5388));
 AOI22xp33_ASAP7_75t_R g152716__5526 (.A1(u0_slt7_r[9]),
    .A2(n_9629),
    .B1(out_slt7[10]),
    .B2(n_9396),
    .Y(n_5387));
 AOI22xp33_ASAP7_75t_R g152718__6783 (.A1(u0_slt7_r[8]),
    .A2(n_9301),
    .B1(out_slt7[9]),
    .B2(n_9348),
    .Y(n_5386));
 AOI22xp33_ASAP7_75t_R g152720__3680 (.A1(u0_slt7_r[7]),
    .A2(n_9300),
    .B1(out_slt7[8]),
    .B2(n_9347),
    .Y(n_5385));
 AOI22xp33_ASAP7_75t_R g152722__1617 (.A1(u0_slt7_r[6]),
    .A2(n_9299),
    .B1(out_slt7[7]),
    .B2(n_9346),
    .Y(n_5384));
 AOI22xp33_ASAP7_75t_R g152724__2802 (.A1(u0_slt7_r[5]),
    .A2(n_9298),
    .B1(out_slt7[6]),
    .B2(n_9345),
    .Y(n_5383));
 AOI22xp33_ASAP7_75t_R g152726__1705 (.A1(u0_slt7_r[4]),
    .A2(n_9630),
    .B1(out_slt7[5]),
    .B2(n_9398),
    .Y(n_5382));
 AOI22xp33_ASAP7_75t_R g152728__5122 (.A1(u0_slt7_r[3]),
    .A2(n_9629),
    .B1(out_slt7[4]),
    .B2(n_9398),
    .Y(n_5381));
 AOI22xp33_ASAP7_75t_R g152730__8246 (.A1(u0_slt7_r[2]),
    .A2(n_9297),
    .B1(out_slt7[3]),
    .B2(n_9344),
    .Y(n_5380));
 AOI22xp33_ASAP7_75t_R g152732__7098 (.A1(u0_slt7_r[1]),
    .A2(n_9630),
    .B1(out_slt7[2]),
    .B2(n_9351),
    .Y(n_5379));
 AOI22xp33_ASAP7_75t_R g152734__6131 (.A1(u0_slt7_r[0]),
    .A2(n_9629),
    .B1(out_slt7[1]),
    .B2(n_9350),
    .Y(n_5378));
 AOI22xp33_ASAP7_75t_R g152736__1881 (.A1(u0_slt8_r[19]),
    .A2(n_9630),
    .B1(out_slt7[0]),
    .B2(n_9349),
    .Y(n_5377));
 AOI22xp33_ASAP7_75t_R g152738__5115 (.A1(u0_slt8_r[18]),
    .A2(n_9629),
    .B1(out_slt8[19]),
    .B2(n_9348),
    .Y(n_5376));
 AOI22xp33_ASAP7_75t_R g152740__7482 (.A1(u0_slt8_r[17]),
    .A2(n_9296),
    .B1(out_slt8[18]),
    .B2(n_9397),
    .Y(n_5375));
 AOI22xp33_ASAP7_75t_R g152742__4733 (.A1(u0_slt8_r[16]),
    .A2(n_9295),
    .B1(out_slt8[17]),
    .B2(n_9347),
    .Y(n_5374));
 AOI22xp33_ASAP7_75t_R g152744__6161 (.A1(u0_slt8_r[15]),
    .A2(n_9294),
    .B1(out_slt8[16]),
    .B2(n_9396),
    .Y(n_5373));
 AOI22xp33_ASAP7_75t_R g152746__9315 (.A1(u0_slt8_r[14]),
    .A2(n_9301),
    .B1(out_slt8[15]),
    .B2(n_9395),
    .Y(n_5372));
 AOI22xp33_ASAP7_75t_R g152748__9945 (.A1(u0_slt8_r[13]),
    .A2(n_5522),
    .B1(out_slt8[14]),
    .B2(n_9346),
    .Y(n_5371));
 AOI22xp33_ASAP7_75t_R g152750__2883 (.A1(u0_slt8_r[12]),
    .A2(n_9300),
    .B1(out_slt8[13]),
    .B2(n_9394),
    .Y(n_5370));
 AOI22xp33_ASAP7_75t_R g152752__2346 (.A1(u0_slt8_r[11]),
    .A2(n_9468),
    .B1(out_slt8[12]),
    .B2(n_9345),
    .Y(n_5369));
 AOI22xp33_ASAP7_75t_R g152754__1666 (.A1(u0_slt8_r[10]),
    .A2(n_9299),
    .B1(out_slt8[11]),
    .B2(n_9395),
    .Y(n_5368));
 AOI22xp33_ASAP7_75t_R g152756__7410 (.A1(u0_slt8_r[9]),
    .A2(n_9467),
    .B1(out_slt8[10]),
    .B2(n_9344),
    .Y(n_5367));
 AOI22xp33_ASAP7_75t_R g152758__6417 (.A1(u0_slt8_r[8]),
    .A2(n_9298),
    .B1(out_slt8[9]),
    .B2(n_9396),
    .Y(n_5366));
 AOI22xp33_ASAP7_75t_R g152760__5477 (.A1(u0_slt8_r[7]),
    .A2(n_9297),
    .B1(out_slt8[8]),
    .B2(n_9351),
    .Y(n_5365));
 AOI22xp33_ASAP7_75t_R g152762__2398 (.A1(u0_slt8_r[6]),
    .A2(n_9296),
    .B1(out_slt8[7]),
    .B2(n_9398),
    .Y(n_5364));
 AOI22xp33_ASAP7_75t_R g152764__5107 (.A1(u0_slt8_r[5]),
    .A2(n_9295),
    .B1(out_slt8[6]),
    .B2(n_9350),
    .Y(n_5363));
 AOI22xp33_ASAP7_75t_R g152766__6260 (.A1(u0_slt8_r[4]),
    .A2(n_9294),
    .B1(out_slt8[5]),
    .B2(n_9349),
    .Y(n_5362));
 AOI22xp33_ASAP7_75t_R g152768__4319 (.A1(u0_slt8_r[3]),
    .A2(n_9630),
    .B1(out_slt8[4]),
    .B2(n_9348),
    .Y(n_5361));
 AOI22xp33_ASAP7_75t_R g152770__8428 (.A1(u0_slt8_r[2]),
    .A2(n_9629),
    .B1(out_slt8[3]),
    .B2(n_9347),
    .Y(n_5360));
 AOI22xp33_ASAP7_75t_R g152772__5526 (.A1(u0_slt8_r[1]),
    .A2(n_9301),
    .B1(out_slt8[2]),
    .B2(n_9398),
    .Y(n_5359));
 AOI22xp33_ASAP7_75t_R g152774__6783 (.A1(u0_slt8_r[0]),
    .A2(n_9630),
    .B1(out_slt8[1]),
    .B2(n_9346),
    .Y(n_5358));
 AOI22xp33_ASAP7_75t_R g152776__3680 (.A1(u0_slt9_r[19]),
    .A2(n_9300),
    .B1(out_slt8[0]),
    .B2(n_9345),
    .Y(n_5357));
 AOI22xp33_ASAP7_75t_R g152778__1617 (.A1(u0_slt9_r[18]),
    .A2(n_9466),
    .B1(out_slt9[19]),
    .B2(n_9397),
    .Y(n_5356));
 AOI22xp33_ASAP7_75t_R g152780__2802 (.A1(u0_slt9_r[17]),
    .A2(n_9299),
    .B1(out_slt9[18]),
    .B2(n_9396),
    .Y(n_5355));
 AOI22xp33_ASAP7_75t_R g152782__1705 (.A1(u0_slt9_r[16]),
    .A2(n_9298),
    .B1(out_slt9[17]),
    .B2(n_9395),
    .Y(n_5354));
 AOI22xp33_ASAP7_75t_R g152784__5122 (.A1(u0_slt9_r[15]),
    .A2(n_9467),
    .B1(out_slt9[16]),
    .B2(n_9394),
    .Y(n_5353));
 AOI22xp33_ASAP7_75t_R g152786__8246 (.A1(u0_slt9_r[14]),
    .A2(n_9297),
    .B1(out_slt9[15]),
    .B2(n_9344),
    .Y(n_5352));
 AOI22xp33_ASAP7_75t_R g152788__7098 (.A1(u0_slt9_r[13]),
    .A2(n_9629),
    .B1(out_slt9[14]),
    .B2(n_9395),
    .Y(n_5351));
 AOI22xp33_ASAP7_75t_R g152790__6131 (.A1(u0_slt9_r[12]),
    .A2(n_9296),
    .B1(out_slt9[13]),
    .B2(n_9396),
    .Y(n_5350));
 AOI22xp33_ASAP7_75t_R g152792__1881 (.A1(u0_slt9_r[11]),
    .A2(n_9295),
    .B1(out_slt9[12]),
    .B2(n_9351),
    .Y(n_5349));
 AOI22xp33_ASAP7_75t_R g152794__5115 (.A1(u0_slt9_r[10]),
    .A2(n_9294),
    .B1(out_slt9[11]),
    .B2(n_9350),
    .Y(n_5348));
 AOI22xp33_ASAP7_75t_R g152796__7410 (.A1(u0_slt9_r[9]),
    .A2(n_9301),
    .B1(out_slt9[10]),
    .B2(n_9398),
    .Y(n_5332));
 AOI22xp33_ASAP7_75t_R g152798__6260 (.A1(u0_slt9_r[8]),
    .A2(n_9300),
    .B1(out_slt9[9]),
    .B2(n_9398),
    .Y(n_5325));
 AOI22xp33_ASAP7_75t_R g152800__8246 (.A1(u0_slt9_r[7]),
    .A2(n_9466),
    .B1(out_slt9[8]),
    .B2(n_9349),
    .Y(n_5314));
 AOI22xp33_ASAP7_75t_R g152802__9945 (.A1(u0_slt9_r[6]),
    .A2(n_9299),
    .B1(out_slt9[7]),
    .B2(n_9348),
    .Y(n_5303));
 AOI22xp33_ASAP7_75t_R g152804__2398 (.A1(u0_slt9_r[5]),
    .A2(n_9298),
    .B1(out_slt9[6]),
    .B2(n_9397),
    .Y(n_5293));
 AOI22xp33_ASAP7_75t_R g152814__7482 (.A1(u1_sr[19]),
    .A2(out_le[4]),
    .B1(in_slt4[19]),
    .B2(n_5341),
    .Y(n_5347));
 AOI22xp33_ASAP7_75t_R g152815__4733 (.A1(u1_sr[19]),
    .A2(out_le[3]),
    .B1(in_slt3[19]),
    .B2(n_5338),
    .Y(n_5346));
 AOI22xp33_ASAP7_75t_R g152816__6161 (.A1(u1_sr[19]),
    .A2(n_11046),
    .B1(in_slt2[19]),
    .B2(n_5336),
    .Y(n_5345));
 AOI22xp33_ASAP7_75t_R g152817__9315 (.A1(u1_sr[19]),
    .A2(out_le[5]),
    .B1(in_slt6[19]),
    .B2(n_5333),
    .Y(n_5344));
 AOI22xp33_ASAP7_75t_R g152818__5122 (.A1(u0_slt9_r[4]),
    .A2(n_9630),
    .B1(out_slt9[5]),
    .B2(n_9347),
    .Y(n_5279));
 AOI22xp33_ASAP7_75t_R g152823__9945 (.A1(u1_sr[18]),
    .A2(n_10709),
    .B1(in_slt4[18]),
    .B2(n_10787),
    .Y(n_5343));
 AOI22xp33_ASAP7_75t_R g152824__2883 (.A1(u1_sr[18]),
    .A2(n_10735),
    .B1(in_slt3[18]),
    .B2(n_10761),
    .Y(n_5340));
 AOI22xp33_ASAP7_75t_R g152825__2346 (.A1(u1_sr[18]),
    .A2(out_le[2]),
    .B1(in_slt2[18]),
    .B2(n_5336),
    .Y(n_5337));
 AOI22xp33_ASAP7_75t_R g152826__1666 (.A1(u1_sr[18]),
    .A2(n_10839),
    .B1(in_slt6[18]),
    .B2(n_10813),
    .Y(n_5335));
 AOI22xp33_ASAP7_75t_R g152832__6417 (.A1(u1_sr[17]),
    .A2(n_10735),
    .B1(in_slt3[17]),
    .B2(n_10761),
    .Y(n_5330));
 AOI22xp33_ASAP7_75t_R g152833__5477 (.A1(u1_sr[17]),
    .A2(out_le[2]),
    .B1(in_slt2[17]),
    .B2(n_5336),
    .Y(n_5329));
 AOI22xp33_ASAP7_75t_R g152835__2398 (.A1(u1_sr[17]),
    .A2(n_10709),
    .B1(in_slt4[17]),
    .B2(n_10787),
    .Y(n_5328));
 AOI22xp33_ASAP7_75t_R g152836__5107 (.A1(u1_sr[17]),
    .A2(n_10839),
    .B1(in_slt6[17]),
    .B2(n_10813),
    .Y(n_5327));
 INVxp33_ASAP7_75t_R g152837 (.A(u1_sr[18]),
    .Y(n_5331));
 AOI22xp33_ASAP7_75t_R g152843__4319 (.A1(u1_sr[16]),
    .A2(out_le[4]),
    .B1(in_slt4[16]),
    .B2(n_5341),
    .Y(n_5324));
 AOI22xp33_ASAP7_75t_R g152844__8428 (.A1(u1_sr[16]),
    .A2(out_le[3]),
    .B1(in_slt3[16]),
    .B2(n_5338),
    .Y(n_5323));
 AOI22xp33_ASAP7_75t_R g152845__5526 (.A1(u1_sr[16]),
    .A2(n_11046),
    .B1(in_slt2[16]),
    .B2(n_5336),
    .Y(n_5322));
 AOI22xp33_ASAP7_75t_R g152846__6783 (.A1(u1_sr[16]),
    .A2(out_le[5]),
    .B1(in_slt6[16]),
    .B2(n_5333),
    .Y(n_5321));
 AOI22xp33_ASAP7_75t_R g152847__2883 (.A1(u0_slt9_r[3]),
    .A2(n_9297),
    .B1(out_slt9[4]),
    .B2(n_9396),
    .Y(n_5266));
 INVxp33_ASAP7_75t_R g152849 (.A(u1_sr[17]),
    .Y(n_5326));
 AOI22xp33_ASAP7_75t_R g152855__3680 (.A1(u1_sr[15]),
    .A2(n_10709),
    .B1(in_slt4[15]),
    .B2(n_10787),
    .Y(n_5319));
 AOI22xp33_ASAP7_75t_R g152856__1617 (.A1(u1_sr[15]),
    .A2(n_10735),
    .B1(in_slt3[15]),
    .B2(n_10761),
    .Y(n_5318));
 AOI22xp33_ASAP7_75t_R g152857__5122 (.A1(u1_sr[15]),
    .A2(out_le[2]),
    .B1(in_slt2[15]),
    .B2(n_5336),
    .Y(n_5315));
 AOI22xp33_ASAP7_75t_R g152858__1705 (.A1(u1_sr[15]),
    .A2(n_10839),
    .B1(in_slt6[15]),
    .B2(n_10813),
    .Y(n_5316));
 AOI22xp33_ASAP7_75t_R g152859__2802 (.A1(out_le[0]),
    .A2(u1_sr[15]),
    .B1(in_slt0[15]),
    .B2(n_5296),
    .Y(n_5317));
 INVxp33_ASAP7_75t_R g152860 (.A(u1_sr[16]),
    .Y(n_5320));
 AOI22xp33_ASAP7_75t_R g152866__7098 (.A1(u1_sr[14]),
    .A2(out_le[3]),
    .B1(in_slt3[14]),
    .B2(n_5338),
    .Y(n_5312));
 AOI22xp33_ASAP7_75t_R g152867__6131 (.A1(u1_sr[14]),
    .A2(n_11046),
    .B1(in_slt2[14]),
    .B2(n_5336),
    .Y(n_5311));
 AOI22xp33_ASAP7_75t_R g152869__1881 (.A1(u1_sr[14]),
    .A2(out_le[4]),
    .B1(in_slt4[14]),
    .B2(n_5341),
    .Y(n_5310));
 AOI22xp33_ASAP7_75t_R g152870__5115 (.A1(u1_sr[14]),
    .A2(out_le[5]),
    .B1(in_slt6[14]),
    .B2(n_5333),
    .Y(n_5309));
 INVxp33_ASAP7_75t_R g152871 (.A(u1_sr[15]),
    .Y(n_5313));
 AOI22xp33_ASAP7_75t_R g152877__7482 (.A1(u1_sr[13]),
    .A2(n_10709),
    .B1(in_slt4[13]),
    .B2(n_10787),
    .Y(n_5307));
 AOI22xp33_ASAP7_75t_R g152878__4733 (.A1(u1_sr[13]),
    .A2(n_10735),
    .B1(in_slt3[13]),
    .B2(n_10761),
    .Y(n_5306));
 AOI22xp33_ASAP7_75t_R g152879__6161 (.A1(u1_sr[13]),
    .A2(out_le[2]),
    .B1(in_slt2[13]),
    .B2(n_5336),
    .Y(n_5305));
 AOI22xp33_ASAP7_75t_R g152880__9315 (.A1(u1_sr[13]),
    .A2(n_10839),
    .B1(in_slt6[13]),
    .B2(n_10813),
    .Y(n_5304));
 AOI22xp33_ASAP7_75t_R g152881__7410 (.A1(u0_slt9_r[2]),
    .A2(n_9296),
    .B1(out_slt9[3]),
    .B2(n_9346),
    .Y(n_4487));
 INVxp33_ASAP7_75t_R g152883 (.A(u1_sr[14]),
    .Y(n_5308));
 AOI22xp33_ASAP7_75t_R g152960__2883 (.A1(u1_sr[12]),
    .A2(out_le[5]),
    .B1(in_slt6[12]),
    .B2(n_5333),
    .Y(n_5301));
 AOI22xp33_ASAP7_75t_R g152961__2346 (.A1(u1_sr[12]),
    .A2(out_le[4]),
    .B1(in_slt4[12]),
    .B2(n_5341),
    .Y(n_5300));
 AOI22xp33_ASAP7_75t_R g152962__1666 (.A1(u1_sr[12]),
    .A2(out_le[3]),
    .B1(in_slt3[12]),
    .B2(n_5338),
    .Y(n_5299));
 AOI22xp33_ASAP7_75t_R g152963__7410 (.A1(u1_sr[12]),
    .A2(n_11046),
    .B1(in_slt2[12]),
    .B2(n_5336),
    .Y(n_5298));
 AOI22xp33_ASAP7_75t_R g152964__6417 (.A1(out_le[0]),
    .A2(u1_sr[12]),
    .B1(in_slt0[12]),
    .B2(n_5296),
    .Y(n_5297));
 NAND2x1_ASAP7_75t_SL g153 (.A(n_48972),
    .B(n_51500),
    .Y(n_48974));
 INVxp33_ASAP7_75t_R g153037 (.A(u1_sr[13]),
    .Y(n_5302));
 AOI22xp5_ASAP7_75t_SL g153290__5526 (.A1(n_30483),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [31]),
    .Y(n_4952));
 AOI22xp5_ASAP7_75t_SL g153291__3680 (.A1(n_4919),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [30]),
    .Y(n_4950));
 AOI22xp5_ASAP7_75t_SL g153292__1705 (.A1(n_4917),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [29]),
    .Y(n_4945));
 AOI22xp5_ASAP7_75t_SL g153293__7098 (.A1(n_4915),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [28]),
    .Y(n_4942));
 AOI22xp5_ASAP7_75t_SL g153294__1881 (.A1(n_4913),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [27]),
    .Y(n_4940));
 AOI22xp5_ASAP7_75t_SL g153295__5115 (.A1(n_4911),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [26]),
    .Y(n_4939));
 AOI22xp5_ASAP7_75t_SL g153296__7482 (.A1(n_4909),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [25]),
    .Y(n_4938));
 AOI22xp5_ASAP7_75t_SL g153297__4733 (.A1(n_4907),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [24]),
    .Y(n_4937));
 AOI22xp33_ASAP7_75t_SL g153298__6161 (.A1(n_4905),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [23]),
    .Y(n_4936));
 AOI22xp5_ASAP7_75t_SL g153299__2883 (.A1(n_4903),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [22]),
    .Y(n_4932));
 AOI22xp33_ASAP7_75t_SL g153300__7410 (.A1(n_4901),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [21]),
    .Y(n_4929));
 AOI22xp5_ASAP7_75t_SL g153301__6417 (.A1(n_4899),
    .A2(n_28953),
    .B1(n_21553),
    .B2(\u11_mem[1] [20]),
    .Y(n_4928));
 AOI22xp5_ASAP7_75t_SL g153302__5122 (.A1(n_24734),
    .A2(n_25681),
    .B1(\u9_mem[1] [31]),
    .B2(n_60873),
    .Y(n_5208));
 AOI22xp5_ASAP7_75t_SL g153303__8246 (.A1(n_24734),
    .A2(n_25680),
    .B1(\u9_mem[1] [30]),
    .B2(n_60873),
    .Y(n_5207));
 AOI22xp5_ASAP7_75t_SL g153304__7098 (.A1(n_25679),
    .A2(n_24734),
    .B1(\u9_mem[1] [29]),
    .B2(n_60873),
    .Y(n_5204));
 AOI22xp5_ASAP7_75t_SL g153305__6131 (.A1(n_25682),
    .A2(n_24734),
    .B1(\u9_mem[1] [28]),
    .B2(n_60873),
    .Y(n_5203));
 AOI22xp5_ASAP7_75t_SL g153306__1881 (.A1(n_5177),
    .A2(n_24734),
    .B1(\u9_mem[1] [27]),
    .B2(n_60873),
    .Y(n_5202));
 AOI22xp5_ASAP7_75t_SL g153307__5115 (.A1(n_5171),
    .A2(n_24734),
    .B1(\u9_mem[1] [26]),
    .B2(n_60873),
    .Y(n_5201));
 AOI22xp5_ASAP7_75t_SL g153308__7482 (.A1(n_24734),
    .A2(n_5173),
    .B1(\u9_mem[1] [25]),
    .B2(n_60873),
    .Y(n_5200));
 AOI22xp5_ASAP7_75t_SL g153309__4733 (.A1(n_25674),
    .A2(n_24734),
    .B1(\u9_mem[1] [24]),
    .B2(n_60873),
    .Y(n_5199));
 AOI22xp5_ASAP7_75t_SL g153310__6161 (.A1(n_25673),
    .A2(n_24734),
    .B1(\u9_mem[1] [23]),
    .B2(n_60873),
    .Y(n_5198));
 AOI22xp5_ASAP7_75t_SL g153311__9315 (.A1(n_5181),
    .A2(n_24734),
    .B1(\u9_mem[1] [22]),
    .B2(n_60873),
    .Y(n_5197));
 AOI22xp5_ASAP7_75t_SL g153312__9945 (.A1(n_5185),
    .A2(n_24734),
    .B1(\u9_mem[1] [21]),
    .B2(n_60873),
    .Y(n_5196));
 AOI22xp5_ASAP7_75t_SL g153313__2883 (.A1(n_25675),
    .A2(n_24734),
    .B1(\u9_mem[1] [20]),
    .B2(n_60873),
    .Y(n_5195));
 AOI22xp5_ASAP7_75t_SL g153314__8428 (.A1(n_29006),
    .A2(n_30483),
    .B1(n_20595),
    .B2(\u11_mem[3] [31]),
    .Y(n_4922));
 AOI22xp5_ASAP7_75t_SL g153315__5526 (.A1(n_4919),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [30]),
    .Y(n_4920));
 AOI22xp5_ASAP7_75t_SL g153316__6783 (.A1(n_4917),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [29]),
    .Y(n_4918));
 AOI22xp5_ASAP7_75t_SL g153317__3680 (.A1(n_4915),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [28]),
    .Y(n_4916));
 AOI22xp5_ASAP7_75t_SL g153318__1617 (.A1(n_4913),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [27]),
    .Y(n_4914));
 AOI22xp33_ASAP7_75t_SL g153319__2802 (.A1(n_4911),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [26]),
    .Y(n_4912));
 AOI22xp5_ASAP7_75t_SL g153320__1705 (.A1(n_4909),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [25]),
    .Y(n_4910));
 AOI22xp5_ASAP7_75t_SL g153321__5122 (.A1(n_4907),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [24]),
    .Y(n_4908));
 AOI22xp33_ASAP7_75t_SL g153322__8246 (.A1(n_4905),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [23]),
    .Y(n_4906));
 AOI22xp33_ASAP7_75t_SL g153323__7098 (.A1(n_4903),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [22]),
    .Y(n_4904));
 AOI22xp5_ASAP7_75t_SL g153324__6131 (.A1(n_4901),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [21]),
    .Y(n_4902));
 AOI22xp33_ASAP7_75t_SL g153325__1881 (.A1(n_29006),
    .A2(n_4899),
    .B1(n_20595),
    .B2(\u11_mem[3] [20]),
    .Y(n_4900));
 AOI22xp5_ASAP7_75t_SL g153330__4319 (.A1(n_24735),
    .A2(n_5177),
    .B1(\u9_mem[3] [27]),
    .B2(n_45330),
    .Y(n_5178));
 AOI22xp5_ASAP7_75t_SL g153331__6783 (.A1(n_5171),
    .A2(n_24735),
    .B1(\u9_mem[3] [26]),
    .B2(n_45330),
    .Y(n_5172));
 AOI22xp5_ASAP7_75t_SL g153335__5115 (.A1(n_24735),
    .A2(n_5181),
    .B1(\u9_mem[3] [22]),
    .B2(n_45330),
    .Y(n_5161));
 AOI22xp5_ASAP7_75t_SL g153336__7482 (.A1(n_24735),
    .A2(n_5185),
    .B1(\u9_mem[3] [21]),
    .B2(n_45330),
    .Y(n_5160));
 AOI22xp5_ASAP7_75t_SL g153337__4733 (.A1(n_24735),
    .A2(n_25675),
    .B1(\u9_mem[3] [20]),
    .B2(n_45330),
    .Y(n_5159));
 O2A1O1Ixp33_ASAP7_75t_SL g153338__5122 (.A1(n_4078),
    .A2(n_24763),
    .B(u26_cnt[2]),
    .C(n_21778),
    .Y(n_4505));
 AOI22xp33_ASAP7_75t_R g153339__5477 (.A1(u1_sr[11]),
    .A2(n_10839),
    .B1(in_slt6[11]),
    .B2(n_10813),
    .Y(n_5294));
 AOI22xp33_ASAP7_75t_R g153340__5107 (.A1(u1_sr[11]),
    .A2(n_10709),
    .B1(in_slt4[11]),
    .B2(n_10787),
    .Y(n_5292));
 AOI22xp33_ASAP7_75t_R g153341__8428 (.A1(u1_sr[11]),
    .A2(n_10735),
    .B1(in_slt3[11]),
    .B2(n_10761),
    .Y(n_5289));
 AOI22xp5_ASAP7_75t_SL g153342__2398 (.A1(n_28953),
    .A2(n_45624),
    .B1(n_21553),
    .B2(\u11_mem[1] [19]),
    .Y(n_4886));
 AOI22xp5_ASAP7_75t_SL g153343__5107 (.A1(n_28953),
    .A2(n_4883),
    .B1(n_21553),
    .B2(\u11_mem[1] [18]),
    .Y(n_4884));
 AOI22xp5_ASAP7_75t_SL g153344__6260 (.A1(n_28953),
    .A2(n_4881),
    .B1(n_21553),
    .B2(\u11_mem[1] [17]),
    .Y(n_4882));
 AOI22xp5_ASAP7_75t_SL g153345__175619 (.A1(n_28953),
    .A2(n_21552),
    .B1(n_21553),
    .B2(\u11_mem[1] [16]),
    .Y(n_21554));
 AOI22xp33_ASAP7_75t_SL g153346__8428 (.A1(n_4877),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [15]),
    .Y(n_4878));
 AOI22xp5_ASAP7_75t_SL g153347__6783 (.A1(n_28953),
    .A2(n_31779),
    .B1(n_20593),
    .B2(\u11_mem[1] [14]),
    .Y(n_4875));
 AOI22xp33_ASAP7_75t_SL g153348__1705 (.A1(n_4869),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [13]),
    .Y(n_4870));
 AOI22xp33_ASAP7_75t_SL g153350__5115 (.A1(n_4956),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [11]),
    .Y(n_4863));
 AOI22xp33_ASAP7_75t_SL g153351__6161 (.A1(n_21317),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [10]),
    .Y(n_4860));
 AOI22xp33_ASAP7_75t_SL g153353__2346 (.A1(n_21321),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [8]),
    .Y(n_4856));
 AOI22xp33_ASAP7_75t_SL g153355__7410 (.A1(n_4851),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [6]),
    .Y(n_4852));
 AOI22xp33_ASAP7_75t_SL g153356__6417 (.A1(n_4849),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [5]),
    .Y(n_4850));
 AOI22xp33_ASAP7_75t_SL g153357__5477 (.A1(n_28953),
    .A2(n_21325),
    .B1(n_20593),
    .B2(\u11_mem[1] [4]),
    .Y(n_4848));
 AOI22xp5_ASAP7_75t_SL g153358__2398 (.A1(n_28953),
    .A2(n_27878),
    .B1(n_20593),
    .B2(\u11_mem[1] [3]),
    .Y(n_4846));
 AOI22xp5_ASAP7_75t_SL g153359__5107 (.A1(n_28953),
    .A2(n_15136),
    .B1(n_20593),
    .B2(\u11_mem[1] [2]),
    .Y(n_4844));
 AOI22xp33_ASAP7_75t_SL g153360__6260 (.A1(n_28953),
    .A2(n_25530),
    .B1(n_20593),
    .B2(\u11_mem[1] [1]),
    .Y(n_4842));
 AOI22xp33_ASAP7_75t_SL g153361__4319 (.A1(n_28953),
    .A2(n_66076),
    .B1(n_20593),
    .B2(\u11_mem[1] [0]),
    .Y(n_4840));
 AOI22xp5_ASAP7_75t_SL g153362__6161 (.A1(n_5211),
    .A2(n_24734),
    .B1(\u9_mem[1] [19]),
    .B2(n_60873),
    .Y(n_5158));
 AOI22xp5_ASAP7_75t_SL g153363__9315 (.A1(n_24734),
    .A2(n_49625),
    .B1(\u9_mem[1] [18]),
    .B2(n_60873),
    .Y(n_5157));
 AOI22xp5_ASAP7_75t_SL g153364__9945 (.A1(n_24734),
    .A2(n_25678),
    .B1(\u9_mem[1] [17]),
    .B2(n_60873),
    .Y(n_5156));
 AOI22xp5_ASAP7_75t_SL g153365__2883 (.A1(n_24734),
    .A2(n_25677),
    .B1(\u9_mem[1] [16]),
    .B2(n_60873),
    .Y(n_5154));
 AOI22xp5_ASAP7_75t_SL g153366__2346 (.A1(n_17599),
    .A2(n_24734),
    .B1(\u9_mem[1] [15]),
    .B2(n_60873),
    .Y(n_5153));
 AOI22xp33_ASAP7_75t_SL g153367__1666 (.A1(n_24734),
    .A2(n_17595),
    .B1(n_60873),
    .B2(\u9_mem[1] [14]),
    .Y(n_5152));
 AOI22xp33_ASAP7_75t_SL g153368__6417 (.A1(n_24734),
    .A2(n_17596),
    .B1(n_60873),
    .B2(\u9_mem[1] [13]),
    .Y(n_5149));
 AOI22xp33_ASAP7_75t_SL g153369__176525 (.A1(n_24734),
    .A2(n_48055),
    .B1(n_60873),
    .B2(\u9_mem[1] [12]),
    .Y(n_22629));
 AOI22xp5_ASAP7_75t_SL g153371__5107 (.A1(n_21534),
    .A2(n_24734),
    .B1(\u9_mem[1] [10]),
    .B2(n_60873),
    .Y(n_5143));
 AOI22xp33_ASAP7_75t_SL g153372__4319 (.A1(n_24734),
    .A2(n_21530),
    .B1(n_60873),
    .B2(\u9_mem[1] [9]),
    .Y(n_5139));
 AOI22xp33_ASAP7_75t_SL g153373__178344 (.A1(n_24734),
    .A2(n_24888),
    .B1(n_60873),
    .B2(\u9_mem[1] [8]),
    .Y(n_24892));
 AOI22xp33_ASAP7_75t_SL g153374__5526 (.A1(n_17591),
    .A2(n_24734),
    .B1(\u9_mem[1] [7]),
    .B2(n_60873),
    .Y(n_5135));
 AOI22xp33_ASAP7_75t_SL g153375__6783 (.A1(n_24734),
    .A2(n_17597),
    .B1(n_60873),
    .B2(\u9_mem[1] [6]),
    .Y(n_5133));
 AOI22xp33_ASAP7_75t_SL g153376__176531 (.A1(n_22632),
    .A2(n_24734),
    .B1(n_60873),
    .B2(\u9_mem[1] [5]),
    .Y(n_22635));
 AOI22xp33_ASAP7_75t_SL g153377__1617 (.A1(n_48642),
    .A2(n_24734),
    .B1(\u9_mem[1] [4]),
    .B2(n_60873),
    .Y(n_5129));
 AOI22xp5_ASAP7_75t_SL g153378__2802 (.A1(n_46562),
    .A2(n_24734),
    .B1(\u9_mem[1] [3]),
    .B2(n_60873),
    .Y(n_5127));
 AOI22xp5_ASAP7_75t_SL g153379__1705 (.A1(n_46558),
    .A2(n_24734),
    .B1(\u9_mem[1] [2]),
    .B2(n_60873),
    .Y(n_5125));
 AOI22xp5_ASAP7_75t_SL g153381__8246 (.A1(n_40712),
    .A2(n_24734),
    .B1(\u9_mem[1] [0]),
    .B2(n_60873),
    .Y(n_5121));
 AOI21xp5_ASAP7_75t_SL g153382__176747 (.A1(n_22922),
    .A2(u16_u5_dma_req_r1),
    .B(n_22923),
    .Y(n_22924));
 AOI21xp5_ASAP7_75t_SL g153386__176754 (.A1(n_30062),
    .A2(u16_u1_dma_req_r1),
    .B(n_22932),
    .Y(n_22933));
 AOI21xp5_ASAP7_75t_SL g153387__176895 (.A1(n_23099),
    .A2(u16_u0_dma_req_r1),
    .B(n_23100),
    .Y(n_23101));
 AOI22xp33_ASAP7_75t_SL g153388__3680 (.A1(n_45624),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [19]),
    .Y(n_4835));
 AOI22xp33_ASAP7_75t_SL g153389__1617 (.A1(n_4883),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [18]),
    .Y(n_4834));
 AOI22xp33_ASAP7_75t_SL g153390__2802 (.A1(n_29006),
    .A2(n_4881),
    .B1(n_20594),
    .B2(\u11_mem[3] [17]),
    .Y(n_4833));
 AOI22xp33_ASAP7_75t_SL g153391__1705 (.A1(n_29006),
    .A2(n_21552),
    .B1(n_20594),
    .B2(\u11_mem[3] [16]),
    .Y(n_4832));
 AOI22xp33_ASAP7_75t_SL g153392__5122 (.A1(n_4877),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [15]),
    .Y(n_4831));
 AOI22xp33_ASAP7_75t_SL g153394__7098 (.A1(n_4869),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [13]),
    .Y(n_4829));
 A2O1A1Ixp33_ASAP7_75t_SL g153395__175376 (.A1(n_340),
    .A2(n_21263),
    .B(n_24734),
    .C(n_521),
    .Y(n_21264));
 A2O1A1Ixp33_ASAP7_75t_SL g153396__174767 (.A1(u11_wp[2]),
    .A2(n_41248),
    .B(n_28953),
    .C(n_659),
    .Y(n_20597));
 OAI21xp5_ASAP7_75t_SL g153397__1881 (.A1(n_24735),
    .A2(n_786),
    .B(n_4544),
    .Y(n_4827));
 OAI21xp5_ASAP7_75t_SL g153398__1617 (.A1(n_29006),
    .A2(n_660),
    .B(n_4392),
    .Y(n_4641));
 NAND2xp5_ASAP7_75t_SL g153399__5115 (.A(n_47616),
    .B(n_521),
    .Y(n_4826));
 AOI22xp33_ASAP7_75t_R g153401__4319 (.A1(out_le[0]),
    .A2(u1_sr[11]),
    .B1(in_slt0[11]),
    .B2(n_5296),
    .Y(n_5290));
 AOI22xp33_ASAP7_75t_R g153402__6260 (.A1(out_le[1]),
    .A2(u1_sr[11]),
    .B1(in_slt1[11]),
    .B2(n_5284),
    .Y(n_5291));
 AOI22xp33_ASAP7_75t_R g153403__5526 (.A1(u1_sr[11]),
    .A2(out_le[2]),
    .B1(in_slt2[11]),
    .B2(n_5336),
    .Y(n_5288));
 AOI22xp5_ASAP7_75t_SL g153404__6131 (.A1(n_24735),
    .A2(n_40712),
    .B1(\u9_mem[3] [0]),
    .B2(n_45330),
    .Y(n_5118));
 AOI22xp33_ASAP7_75t_SL g153408__4733 (.A1(n_24735),
    .A2(n_48642),
    .B1(\u9_mem[3] [4]),
    .B2(n_45330),
    .Y(n_5114));
 AOI22xp33_ASAP7_75t_SL g153409__6161 (.A1(n_24735),
    .A2(n_22632),
    .B1(\u9_mem[3] [5]),
    .B2(n_45330),
    .Y(n_5113));
 AOI22xp33_ASAP7_75t_SL g153410__9315 (.A1(n_24735),
    .A2(n_17597),
    .B1(\u9_mem[3] [6]),
    .B2(n_45330),
    .Y(n_5112));
 AOI22xp33_ASAP7_75t_SL g153411__9945 (.A1(n_24735),
    .A2(n_17591),
    .B1(\u9_mem[3] [7]),
    .B2(n_45330),
    .Y(n_5111));
 AOI22xp33_ASAP7_75t_SL g153412__178339 (.A1(n_24735),
    .A2(n_24888),
    .B1(\u9_mem[3] [8]),
    .B2(n_45330),
    .Y(n_24889));
 AOI22xp33_ASAP7_75t_SL g153413__175598 (.A1(n_24735),
    .A2(n_21530),
    .B1(\u9_mem[3] [9]),
    .B2(n_45330),
    .Y(n_21532));
 AOI22xp33_ASAP7_75t_SL g153414__175602 (.A1(n_24735),
    .A2(n_21534),
    .B1(\u9_mem[3] [10]),
    .B2(n_45330),
    .Y(n_21536));
 AOI22xp33_ASAP7_75t_SL g153416__6417 (.A1(n_24735),
    .A2(n_48055),
    .B1(\u9_mem[3] [12]),
    .B2(n_45330),
    .Y(n_5106));
 AOI22xp5_ASAP7_75t_SL g153417__5477 (.A1(n_24735),
    .A2(n_17596),
    .B1(\u9_mem[3] [13]),
    .B2(n_45330),
    .Y(n_5105));
 AOI22xp33_ASAP7_75t_SL g153418__2398 (.A1(n_24735),
    .A2(n_17595),
    .B1(\u9_mem[3] [14]),
    .B2(n_45330),
    .Y(n_5104));
 AOI22xp33_ASAP7_75t_SL g153419__5107 (.A1(n_24735),
    .A2(n_17599),
    .B1(n_45330),
    .B2(\u9_mem[3] [15]),
    .Y(n_5103));
 AOI22xp5_ASAP7_75t_SL g153420__6260 (.A1(n_24735),
    .A2(n_25677),
    .B1(\u9_mem[3] [16]),
    .B2(n_45330),
    .Y(n_5101));
 AOI22xp5_ASAP7_75t_SL g153421__4319 (.A1(n_24735),
    .A2(n_25678),
    .B1(\u9_mem[3] [17]),
    .B2(n_45330),
    .Y(n_5100));
 AOI22xp5_ASAP7_75t_SL g153423__1705 (.A1(n_5211),
    .A2(n_24735),
    .B1(\u9_mem[3] [19]),
    .B2(n_45330),
    .Y(n_5212));
 AOI22xp5_ASAP7_75t_SL g153424__4733 (.A1(n_29006),
    .A2(n_66076),
    .B1(n_20594),
    .B2(\u11_mem[3] [0]),
    .Y(n_4824));
 AOI22xp33_ASAP7_75t_SL g153425__6161 (.A1(n_29006),
    .A2(n_25530),
    .B1(n_20594),
    .B2(\u11_mem[3] [1]),
    .Y(n_4823));
 AOI22xp33_ASAP7_75t_SL g153428__2346 (.A1(n_21325),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [4]),
    .Y(n_4819));
 AOI22xp33_ASAP7_75t_SL g153429__7410 (.A1(n_4849),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [5]),
    .Y(n_4817));
 AOI22xp33_ASAP7_75t_SL g153430__1666 (.A1(n_4851),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [6]),
    .Y(n_4818));
 AOI22xp33_ASAP7_75t_SL g153432__7482 (.A1(n_21321),
    .A2(n_29006),
    .B1(n_20594),
    .B2(\u11_mem[3] [8]),
    .Y(n_4825));
 AOI22xp33_ASAP7_75t_SL g153433__8428 (.A1(n_31777),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [9]),
    .Y(n_4992));
 AOI22xp33_ASAP7_75t_SL g153434__5526 (.A1(n_21317),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [10]),
    .Y(n_5098));
 AOI22xp33_ASAP7_75t_SL g153435__6783 (.A1(n_4956),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [11]),
    .Y(n_5097));
 AOI22xp33_ASAP7_75t_SL g153436__3680 (.A1(n_31781),
    .A2(n_29006),
    .B1(n_20595),
    .B2(\u11_mem[3] [12]),
    .Y(n_5094));
 INVxp33_ASAP7_75t_R g153542 (.A(u1_sr[12]),
    .Y(n_5295));
 AOI22xp33_ASAP7_75t_SL g153543__168321 (.A1(n_12871),
    .A2(n_17599),
    .B1(\u9_mem[2] [15]),
    .B2(n_5258),
    .Y(n_12895));
 AOI22xp33_ASAP7_75t_SL g153544__168301 (.A1(n_12869),
    .A2(n_17595),
    .B1(\u9_mem[2] [14]),
    .B2(n_5258),
    .Y(n_12875));
 AOI22xp33_ASAP7_75t_SL g153545__168318 (.A1(n_12871),
    .A2(n_17596),
    .B1(n_5258),
    .B2(\u9_mem[2] [13]),
    .Y(n_12892));
 AOI22xp33_ASAP7_75t_SL g153546__168328 (.A1(n_12871),
    .A2(n_48055),
    .B1(\u9_mem[2] [12]),
    .B2(n_5258),
    .Y(n_12902));
 AOI22xp33_ASAP7_75t_SL g153547__168319 (.A1(n_12871),
    .A2(n_15693),
    .B1(\u9_mem[2] [11]),
    .B2(n_5258),
    .Y(n_12893));
 AOI22xp33_ASAP7_75t_SL g153548__168315 (.A1(n_12871),
    .A2(n_21534),
    .B1(\u9_mem[2] [10]),
    .B2(n_5258),
    .Y(n_12889));
 AOI22xp33_ASAP7_75t_SL g153549__168316 (.A1(n_12871),
    .A2(n_21530),
    .B1(\u9_mem[2] [9]),
    .B2(n_5258),
    .Y(n_12890));
 AOI22xp33_ASAP7_75t_SL g153550__178342 (.A1(n_12871),
    .A2(n_24888),
    .B1(\u9_mem[2] [8]),
    .B2(n_5258),
    .Y(n_24890));
 AOI22xp33_ASAP7_75t_SL g153551__168327 (.A1(n_12871),
    .A2(n_17591),
    .B1(n_5258),
    .B2(\u9_mem[2] [7]),
    .Y(n_12901));
 AOI22xp33_ASAP7_75t_SL g153552__168299 (.A1(n_12869),
    .A2(n_17597),
    .B1(n_5258),
    .B2(\u9_mem[2] [6]),
    .Y(n_12873));
 AOI22xp33_ASAP7_75t_SL g153553__168326 (.A1(n_12871),
    .A2(n_22632),
    .B1(\u9_mem[2] [5]),
    .B2(n_5258),
    .Y(n_12900));
 AOI22xp5_ASAP7_75t_SL g153555__168325 (.A1(n_46562),
    .A2(n_12871),
    .B1(\u9_mem[2] [3]),
    .B2(n_5258),
    .Y(n_12899));
 AOI22xp5_ASAP7_75t_SL g153556__168324 (.A1(n_46558),
    .A2(n_12871),
    .B1(\u9_mem[2] [2]),
    .B2(n_5258),
    .Y(n_12898));
 AOI22xp5_ASAP7_75t_SL g153557__168323 (.A1(n_12482),
    .A2(n_12871),
    .B1(\u9_mem[2] [1]),
    .B2(n_5258),
    .Y(n_12897));
 AOI22xp5_ASAP7_75t_SL g153558__168322 (.A1(n_40712),
    .A2(n_12871),
    .B1(\u9_mem[2] [0]),
    .B2(n_5258),
    .Y(n_12896));
 AOI22xp5_ASAP7_75t_SL g153559__3680 (.A1(n_5211),
    .A2(n_31720),
    .B1(\u9_mem[0] [19]),
    .B2(n_46587),
    .Y(n_5020));
 AOI22xp5_ASAP7_75t_SL g153561__2802 (.A1(n_31720),
    .A2(n_25678),
    .B1(\u9_mem[0] [17]),
    .B2(n_46587),
    .Y(n_5016));
 AOI22xp5_ASAP7_75t_SL g153562__1705 (.A1(n_31720),
    .A2(n_25677),
    .B1(\u9_mem[0] [16]),
    .B2(n_46587),
    .Y(n_5015));
 AOI22xp33_ASAP7_75t_SL g153563__5122 (.A1(n_17599),
    .A2(n_31720),
    .B1(\u9_mem[0] [15]),
    .B2(n_46587),
    .Y(n_5014));
 AOI22xp33_ASAP7_75t_SL g153564__8246 (.A1(n_17595),
    .A2(n_31720),
    .B1(\u9_mem[0] [14]),
    .B2(n_46587),
    .Y(n_5012));
 AOI22xp33_ASAP7_75t_SL g153565__7098 (.A1(n_17596),
    .A2(n_31720),
    .B1(\u9_mem[0] [13]),
    .B2(n_46587),
    .Y(n_5011));
 AOI22xp5_ASAP7_75t_SL g153566__6131 (.A1(n_48055),
    .A2(n_31720),
    .B1(\u9_mem[0] [12]),
    .B2(n_46587),
    .Y(n_5010));
 AOI22xp5_ASAP7_75t_SL g153567__1881 (.A1(n_15693),
    .A2(n_31720),
    .B1(\u9_mem[0] [11]),
    .B2(n_46587),
    .Y(n_5009));
 AOI22xp33_ASAP7_75t_SL g153568__5115 (.A1(n_21534),
    .A2(n_31720),
    .B1(\u9_mem[0] [10]),
    .B2(n_46587),
    .Y(n_5008));
 AOI22xp33_ASAP7_75t_SL g153569__7482 (.A1(n_21530),
    .A2(n_31720),
    .B1(\u9_mem[0] [9]),
    .B2(n_46587),
    .Y(n_5007));
 AOI22xp5_ASAP7_75t_SL g153570__178343 (.A1(n_24888),
    .A2(n_31720),
    .B1(\u9_mem[0] [8]),
    .B2(n_46587),
    .Y(n_24891));
 AOI22xp5_ASAP7_75t_SL g153571__6161 (.A1(n_17591),
    .A2(n_31720),
    .B1(\u9_mem[0] [7]),
    .B2(n_46587),
    .Y(n_5005));
 AOI22xp33_ASAP7_75t_SL g153572__9315 (.A1(n_17597),
    .A2(n_31720),
    .B1(\u9_mem[0] [6]),
    .B2(n_46587),
    .Y(n_5004));
 AOI22xp33_ASAP7_75t_SL g153573__9945 (.A1(n_22632),
    .A2(n_31720),
    .B1(\u9_mem[0] [5]),
    .B2(n_46587),
    .Y(n_5003));
 AOI22xp33_ASAP7_75t_SL g153574__2883 (.A1(n_48642),
    .A2(n_31720),
    .B1(\u9_mem[0] [4]),
    .B2(n_46587),
    .Y(n_5002));
 AOI22xp5_ASAP7_75t_SL g153575__1666 (.A1(n_31720),
    .A2(n_46562),
    .B1(\u9_mem[0] [3]),
    .B2(n_46587),
    .Y(n_5000));
 AOI22xp5_ASAP7_75t_SL g153576__7410 (.A1(n_31720),
    .A2(n_46558),
    .B1(\u9_mem[0] [2]),
    .B2(n_46587),
    .Y(n_4999));
 AOI22xp5_ASAP7_75t_SL g153577__6417 (.A1(n_12482),
    .A2(n_31720),
    .B1(\u9_mem[0] [1]),
    .B2(n_46587),
    .Y(n_4998));
 AOI221xp5_ASAP7_75t_SL g153579__213705 (.A1(n_15094),
    .A2(n_79104),
    .B1(out_slt6[19]),
    .B2(n_66659),
    .C(n_38375),
    .Y(n_66663));
 AOI221xp5_ASAP7_75t_SL g153584__6783 (.A1(n_31863),
    .A2(out_slt3[18]),
    .B1(n_25405),
    .B2(n_2539),
    .C(n_4408),
    .Y(n_5021));
 AOI221xp5_ASAP7_75t_SL g153585__5526 (.A1(n_31863),
    .A2(out_slt3[17]),
    .B1(n_25405),
    .B2(n_14864),
    .C(n_4407),
    .Y(n_5022));
 AOI21xp5_ASAP7_75t_SL g153586__8428 (.A1(n_25405),
    .A2(n_2686),
    .B(n_4495),
    .Y(n_5023));
 AOI22xp33_ASAP7_75t_R g153589__6783 (.A1(u1_sr[10]),
    .A2(n_11046),
    .B1(in_slt2[10]),
    .B2(n_5336),
    .Y(n_5286));
 AOI22xp33_ASAP7_75t_R g153590__3680 (.A1(u1_sr[10]),
    .A2(out_le[1]),
    .B1(in_slt1[10]),
    .B2(n_5284),
    .Y(n_5285));
 NAND2xp5_ASAP7_75t_SL g153591__6783 (.A(n_4232),
    .B(n_557),
    .Y(n_4578));
 AOI221xp5_ASAP7_75t_SL g153592__219228 (.A1(n_5028),
    .A2(n_79208),
    .B1(out_slt9[7]),
    .B2(n_73301),
    .C(n_4369),
    .Y(n_73310));
 AOI221xp5_ASAP7_75t_SL g153593__219227 (.A1(n_5028),
    .A2(n_23661),
    .B1(out_slt9[6]),
    .B2(n_73301),
    .C(n_4371),
    .Y(n_73309));
 AOI221xp5_ASAP7_75t_SL g153594__219232 (.A1(n_73301),
    .A2(out_slt9[5]),
    .B1(n_5028),
    .B2(n_2435),
    .C(n_4372),
    .Y(n_73314));
 AOI221xp5_ASAP7_75t_SL g153595__219229 (.A1(n_73301),
    .A2(out_slt9[4]),
    .B1(n_5028),
    .B2(n_2433),
    .C(n_4374),
    .Y(n_73311));
 AOI221x1_ASAP7_75t_SL g153599__2346 (.A1(n_31863),
    .A2(out_slt3[4]),
    .B1(n_25405),
    .B2(n_7572),
    .C(n_4451),
    .Y(n_5036));
 AOI221xp5_ASAP7_75t_SL g153600__193163 (.A1(n_42253),
    .A2(out_slt8[7]),
    .B1(n_50295),
    .B2(n_5077),
    .C(n_4450),
    .Y(n_42264));
 AOI221xp5_ASAP7_75t_SL g153601__193160 (.A1(n_42253),
    .A2(out_slt8[6]),
    .B1(n_5077),
    .B2(n_36843),
    .C(n_4445),
    .Y(n_42261));
 AOI221xp5_ASAP7_75t_SL g153602__193161 (.A1(n_42253),
    .A2(out_slt8[5]),
    .B1(n_5077),
    .B2(n_2385),
    .C(n_4441),
    .Y(n_42262));
 AOI221xp5_ASAP7_75t_SL g153603__6161 (.A1(n_4225),
    .A2(out_slt8[4]),
    .B1(n_5077),
    .B2(n_2429),
    .C(n_4438),
    .Y(n_5041));
 AOI221xp5_ASAP7_75t_SL g153607__179418 (.A1(n_36361),
    .A2(out_slt7[4]),
    .B1(n_25954),
    .B2(n_49182),
    .C(n_4410),
    .Y(n_26103));
 AOI221xp5_ASAP7_75t_SL g153611__185128 (.A1(n_43087),
    .A2(out_slt4[4]),
    .B1(n_32582),
    .B2(n_36013),
    .C(n_4541),
    .Y(n_32600));
 OAI21xp5_ASAP7_75t_SL g153616__5526 (.A1(n_61242),
    .A2(n_1029),
    .B(n_4224),
    .Y(n_4579));
 AOI221xp5_ASAP7_75t_SL g153618__185117 (.A1(n_2337),
    .A2(n_32582),
    .B1(n_43087),
    .B2(out_slt4[17]),
    .C(n_4572),
    .Y(n_32589));
 AOI21xp5_ASAP7_75t_SL g153619__185121 (.A1(n_32582),
    .A2(n_2579),
    .B(n_4614),
    .Y(n_32593));
 AOI21xp5_ASAP7_75t_SL g153624__185113 (.A1(n_32582),
    .A2(n_49320),
    .B(n_46701),
    .Y(n_32584));
 A2O1A1Ixp33_ASAP7_75t_SL g153625__179916 (.A1(u10_wp[2]),
    .A2(n_26645),
    .B(n_24803),
    .C(n_557),
    .Y(n_26646));
 O2A1O1Ixp5_ASAP7_75t_SL g153627__169861 (.A1(n_36082),
    .A2(n_4146),
    .B(u15_crac_rd),
    .C(n_2947),
    .Y(n_14816));
 O2A1O1Ixp33_ASAP7_75t_SL g153628__178191 (.A1(n_24730),
    .A2(n_13420),
    .B(n_24732),
    .C(n_4542),
    .Y(n_24733));
 O2A1O1Ixp33_ASAP7_75t_SL g153629__182014 (.A1(n_28948),
    .A2(n_23286),
    .B(n_28950),
    .C(n_4390),
    .Y(n_28951));
 AOI221xp5_ASAP7_75t_SL g153631__1617 (.A1(n_5024),
    .A2(out_slt3[19]),
    .B1(n_25405),
    .B2(n_2594),
    .C(n_4409),
    .Y(n_5054));
 AOI21xp5_ASAP7_75t_SL g153632__179287 (.A1(n_2363),
    .A2(n_25954),
    .B(n_28412),
    .Y(n_25955));
 AOI21xp5_ASAP7_75t_SL g153633__188954 (.A1(n_37140),
    .A2(n_25956),
    .B(n_34841),
    .Y(n_37141));
 AOI221xp5_ASAP7_75t_SL g153634__188333 (.A1(n_22060),
    .A2(n_25954),
    .B1(out_slt7[10]),
    .B2(n_36361),
    .C(n_4418),
    .Y(n_36366));
 AOI221xp5_ASAP7_75t_SL g153635__188335 (.A1(n_25956),
    .A2(n_78813),
    .B1(out_slt7[11]),
    .B2(n_36361),
    .C(n_22842),
    .Y(n_36367));
 AOI221xp5_ASAP7_75t_SL g153639__182909 (.A1(n_36361),
    .A2(out_slt7[15]),
    .B1(n_25956),
    .B2(n_17706),
    .C(n_4430),
    .Y(n_29948));
 AOI21xp5_ASAP7_75t_SL g153643__1666 (.A1(n_2509),
    .A2(n_5077),
    .B(n_4464),
    .Y(n_5071));
 AOI21xp5_ASAP7_75t_SL g153644__2346 (.A1(n_2513),
    .A2(n_5077),
    .B(n_4462),
    .Y(n_5072));
 AOI21xp5_ASAP7_75t_SL g153645__2883 (.A1(n_2541),
    .A2(n_5077),
    .B(n_4461),
    .Y(n_5073));
 AOI21xp5_ASAP7_75t_SL g153646__9945 (.A1(n_43721),
    .A2(n_5077),
    .B(n_4460),
    .Y(n_5074));
 AOI21xp5_ASAP7_75t_SL g153648__196988 (.A1(n_5077),
    .A2(n_46566),
    .B(n_51160),
    .Y(n_46567));
 AOI21xp5_ASAP7_75t_SL g153651__5115 (.A1(n_25405),
    .A2(n_49500),
    .B(n_4484),
    .Y(n_5081));
 AOI21xp5_ASAP7_75t_SL g153652__1881 (.A1(n_25405),
    .A2(n_46231),
    .B(n_4486),
    .Y(n_5082));
 AOI21xp5_ASAP7_75t_SL g153655__8246 (.A1(n_36531),
    .A2(n_5091),
    .B(n_4525),
    .Y(n_5087));
 AOI21xp5_ASAP7_75t_SL g153656__5122 (.A1(n_2447),
    .A2(n_5091),
    .B(n_17184),
    .Y(n_5088));
 AOI221xp5_ASAP7_75t_SL g153659__1617 (.A1(n_4988),
    .A2(out_slt9[12]),
    .B1(n_5091),
    .B2(n_2348),
    .C(n_4361),
    .Y(n_5093));
 AOI221xp5_ASAP7_75t_SL g153662__6783 (.A1(n_4988),
    .A2(out_slt9[18]),
    .B1(n_5028),
    .B2(n_27136),
    .C(n_4342),
    .Y(n_4990));
 OAI21xp33_ASAP7_75t_SL g153664__176232 (.A1(oc0_int_set[0]),
    .A2(n_2079),
    .B(n_22268),
    .Y(n_22271));
 OAI21xp33_ASAP7_75t_SL g153665__176236 (.A1(oc1_int_set[0]),
    .A2(n_2106),
    .B(n_22268),
    .Y(n_22275));
 OAI21xp33_ASAP7_75t_SL g153666__176235 (.A1(oc2_int_set[0]),
    .A2(n_2095),
    .B(n_22268),
    .Y(n_22274));
 OAI21xp33_ASAP7_75t_SL g153667__176231 (.A1(oc3_int_set[0]),
    .A2(n_2065),
    .B(n_22268),
    .Y(n_22270));
 OAI21xp33_ASAP7_75t_SL g153668__176233 (.A1(oc4_int_set[0]),
    .A2(n_2130),
    .B(n_22268),
    .Y(n_22272));
 OAI21xp33_ASAP7_75t_SL g153669__176234 (.A1(oc5_int_set[0]),
    .A2(u13_ints_r[17]),
    .B(n_22268),
    .Y(n_22273));
 AOI21xp5_ASAP7_75t_SL g153675__171918 (.A1(n_7511),
    .A2(n_4976),
    .B(n_38370),
    .Y(n_17304));
 AOI21xp5_ASAP7_75t_SL g153677__185118 (.A1(n_2584),
    .A2(n_32585),
    .B(n_4617),
    .Y(n_32590));
 AOI322xp5_ASAP7_75t_SL g153760__193866 (.A1(n_32582),
    .A2(n_1892),
    .A3(n_4548),
    .B1(n_31748),
    .B2(n_7803),
    .C1(n_43088),
    .C2(n_42779),
    .Y(n_43091));
 AOI22xp5_ASAP7_75t_SL g153761__168317 (.A1(n_12871),
    .A2(n_25678),
    .B1(\u9_mem[2] [17]),
    .B2(n_5258),
    .Y(n_12891));
 AOI22xp5_ASAP7_75t_SL g153762__168314 (.A1(n_12871),
    .A2(n_49625),
    .B1(\u9_mem[2] [18]),
    .B2(n_5258),
    .Y(n_12888));
 AOI22xp33_ASAP7_75t_SL g153763__168294 (.A1(n_12869),
    .A2(n_5211),
    .B1(n_5258),
    .B2(\u9_mem[2] [19]),
    .Y(n_12870));
 AOI221xp5_ASAP7_75t_SL g153764__169153 (.A1(n_27128),
    .A2(n_36383),
    .B1(n_34235),
    .B2(n_36628),
    .C(n_4092),
    .Y(n_13976));
 AOI22xp5_ASAP7_75t_SL g153766__178451 (.A1(n_61242),
    .A2(n_40956),
    .B1(\u10_mem[3] [0]),
    .B2(n_61244),
    .Y(n_25004));
 AOI22xp5_ASAP7_75t_SL g153767__178449 (.A1(n_61242),
    .A2(n_48456),
    .B1(n_61244),
    .B2(\u10_mem[3] [1]),
    .Y(n_25002));
 AOI22xp5_ASAP7_75t_SL g153768__178448 (.A1(n_61242),
    .A2(n_62614),
    .B1(\u10_mem[3] [2]),
    .B2(n_61244),
    .Y(n_25001));
 AOI22xp5_ASAP7_75t_SL g153770__178446 (.A1(n_50555),
    .A2(n_61242),
    .B1(\u10_mem[3] [4]),
    .B2(n_61244),
    .Y(n_24999));
 AOI22xp5_ASAP7_75t_SL g153771__178445 (.A1(n_61242),
    .A2(n_50553),
    .B1(n_61244),
    .B2(\u10_mem[3] [5]),
    .Y(n_24998));
 AOI22xp5_ASAP7_75t_SL g153772__178444 (.A1(n_61242),
    .A2(n_65879),
    .B1(\u10_mem[3] [6]),
    .B2(n_61244),
    .Y(n_24997));
 AOI22xp33_ASAP7_75t_SL g153773__188371 (.A1(n_61242),
    .A2(n_50552),
    .B1(n_61244),
    .B2(\u10_mem[3] [7]),
    .Y(n_36405));
 AOI22xp5_ASAP7_75t_SL g153774__178442 (.A1(n_61242),
    .A2(n_31786),
    .B1(\u10_mem[3] [8]),
    .B2(n_61244),
    .Y(n_24995));
 AOI22xp5_ASAP7_75t_SL g153775__178441 (.A1(n_61242),
    .A2(n_18707),
    .B1(\u10_mem[3] [9]),
    .B2(n_35121),
    .Y(n_24993));
 AOI22xp5_ASAP7_75t_SL g153776__178440 (.A1(n_61242),
    .A2(n_46479),
    .B1(\u10_mem[3] [10]),
    .B2(n_35121),
    .Y(n_24992));
 AOI22xp5_ASAP7_75t_SL g153778__178439 (.A1(n_61242),
    .A2(n_28747),
    .B1(n_35121),
    .B2(\u10_mem[3] [12]),
    .Y(n_24991));
 AOI22xp33_ASAP7_75t_SL g153779__178438 (.A1(n_61242),
    .A2(n_17613),
    .B1(n_35121),
    .B2(\u10_mem[3] [13]),
    .Y(n_24990));
 AOI22xp33_ASAP7_75t_SL g153780__178437 (.A1(n_61242),
    .A2(n_17614),
    .B1(n_35121),
    .B2(\u10_mem[3] [14]),
    .Y(n_24989));
 AOI22xp33_ASAP7_75t_SL g153781__178436 (.A1(n_61242),
    .A2(n_17615),
    .B1(n_35121),
    .B2(\u10_mem[3] [15]),
    .Y(n_24988));
 AOI22xp5_ASAP7_75t_SL g153782__178435 (.A1(n_61242),
    .A2(n_4712),
    .B1(n_35121),
    .B2(\u10_mem[3] [16]),
    .Y(n_24987));
 AOI22xp5_ASAP7_75t_SL g153783__178434 (.A1(n_61242),
    .A2(n_4710),
    .B1(n_35121),
    .B2(\u10_mem[3] [17]),
    .Y(n_24986));
 AOI22xp5_ASAP7_75t_SL g153784__178433 (.A1(n_61242),
    .A2(n_50549),
    .B1(n_35121),
    .B2(\u10_mem[3] [18]),
    .Y(n_24985));
 AOI22xp33_ASAP7_75t_SL g153788__182080 (.A1(n_66076),
    .A2(n_29008),
    .B1(\u11_mem[0] [0]),
    .B2(n_4784),
    .Y(n_29019));
 AOI22xp5_ASAP7_75t_SL g153790__182072 (.A1(n_25530),
    .A2(n_29011),
    .B1(\u11_mem[0] [1]),
    .B2(n_4784),
    .Y(n_29012));
 AOI22xp5_ASAP7_75t_SL g153791__182078 (.A1(n_15136),
    .A2(n_29008),
    .B1(\u11_mem[0] [2]),
    .B2(n_4784),
    .Y(n_29017));
 AOI22xp5_ASAP7_75t_SL g153792__182075 (.A1(n_27878),
    .A2(n_29008),
    .B1(\u11_mem[0] [3]),
    .B2(n_4784),
    .Y(n_29014));
 AOI22xp33_ASAP7_75t_SL g153793__182084 (.A1(n_21325),
    .A2(n_29008),
    .B1(\u11_mem[0] [4]),
    .B2(n_4784),
    .Y(n_29023));
 AOI22xp33_ASAP7_75t_SL g153794__182094 (.A1(n_29011),
    .A2(n_4849),
    .B1(n_4784),
    .B2(\u11_mem[0] [5]),
    .Y(n_29033));
 AOI22xp5_ASAP7_75t_SL g153795__182086 (.A1(n_4851),
    .A2(n_29008),
    .B1(\u11_mem[0] [6]),
    .B2(n_4784),
    .Y(n_29025));
 AOI22xp33_ASAP7_75t_SL g153797__182082 (.A1(n_21321),
    .A2(n_29008),
    .B1(n_4784),
    .B2(\u11_mem[0] [8]),
    .Y(n_29021));
 AOI22xp33_ASAP7_75t_SL g153798__182071 (.A1(n_31777),
    .A2(n_29008),
    .B1(n_4784),
    .B2(\u11_mem[0] [9]),
    .Y(n_29010));
 AOI22xp33_ASAP7_75t_SL g153799__182068 (.A1(n_29008),
    .A2(n_21317),
    .B1(n_4784),
    .B2(\u11_mem[0] [10]),
    .Y(n_29009));
 AOI22xp5_ASAP7_75t_SL g153801__182083 (.A1(n_31781),
    .A2(n_29008),
    .B1(\u11_mem[0] [12]),
    .B2(n_4784),
    .Y(n_29022));
 AOI22xp33_ASAP7_75t_SL g153802__182074 (.A1(n_4869),
    .A2(n_29008),
    .B1(\u11_mem[0] [13]),
    .B2(n_4784),
    .Y(n_29013));
 AOI22xp33_ASAP7_75t_SL g153803__182081 (.A1(n_31779),
    .A2(n_29008),
    .B1(\u11_mem[0] [14]),
    .B2(n_4784),
    .Y(n_29020));
 AOI22xp33_ASAP7_75t_SL g153804__182077 (.A1(n_4877),
    .A2(n_29008),
    .B1(\u11_mem[0] [15]),
    .B2(n_4784),
    .Y(n_29016));
 AOI22xp5_ASAP7_75t_SL g153805__182079 (.A1(n_21552),
    .A2(n_29008),
    .B1(\u11_mem[0] [16]),
    .B2(n_4784),
    .Y(n_29018));
 AOI22xp5_ASAP7_75t_SL g153806__182097 (.A1(n_29011),
    .A2(n_4881),
    .B1(\u11_mem[0] [17]),
    .B2(n_4784),
    .Y(n_29036));
 AOI22xp33_ASAP7_75t_SL g153807__182076 (.A1(n_4883),
    .A2(n_29008),
    .B1(\u11_mem[0] [18]),
    .B2(n_4784),
    .Y(n_29015));
 AOI22xp5_ASAP7_75t_SL g153808__182089 (.A1(n_29011),
    .A2(n_45624),
    .B1(\u11_mem[0] [19]),
    .B2(n_4784),
    .Y(n_29028));
 AOI22xp5_ASAP7_75t_SL g153810__168293 (.A1(n_25530),
    .A2(n_28520),
    .B1(\u11_mem[2] [1]),
    .B2(n_61785),
    .Y(n_12867));
 AOI22xp5_ASAP7_75t_SL g153811__168291 (.A1(n_15136),
    .A2(n_28520),
    .B1(\u11_mem[2] [2]),
    .B2(n_61785),
    .Y(n_12865));
 AOI22xp33_ASAP7_75t_SL g153813__175430 (.A1(n_45625),
    .A2(n_21325),
    .B1(n_61785),
    .B2(\u11_mem[2] [4]),
    .Y(n_21328));
 AOI22xp33_ASAP7_75t_SL g153814__168277 (.A1(n_45625),
    .A2(n_4849),
    .B1(\u11_mem[2] [5]),
    .B2(n_61785),
    .Y(n_12851));
 AOI22xp5_ASAP7_75t_SL g153815__168289 (.A1(n_28520),
    .A2(n_4851),
    .B1(\u11_mem[2] [6]),
    .B2(n_61785),
    .Y(n_12863));
 AOI22xp33_ASAP7_75t_SL g153817__175426 (.A1(n_28520),
    .A2(n_21321),
    .B1(\u11_mem[2] [8]),
    .B2(n_61785),
    .Y(n_21324));
 AOI22xp5_ASAP7_75t_SL g153818__168287 (.A1(n_31777),
    .A2(n_28520),
    .B1(\u11_mem[2] [9]),
    .B2(n_61785),
    .Y(n_12861));
 AOI22xp33_ASAP7_75t_SL g153819__175422 (.A1(n_28520),
    .A2(n_21317),
    .B1(\u11_mem[2] [10]),
    .B2(n_61785),
    .Y(n_21320));
 AOI22xp33_ASAP7_75t_SL g153820__168262 (.A1(n_28520),
    .A2(n_4956),
    .B1(\u11_mem[2] [11]),
    .B2(n_61785),
    .Y(n_12837));
 AOI22xp33_ASAP7_75t_SL g153821__168285 (.A1(n_31781),
    .A2(n_28520),
    .B1(n_61785),
    .B2(\u11_mem[2] [12]),
    .Y(n_12859));
 AOI22xp33_ASAP7_75t_SL g153822__168284 (.A1(n_28520),
    .A2(n_4869),
    .B1(n_61785),
    .B2(\u11_mem[2] [13]),
    .Y(n_12858));
 AOI22xp33_ASAP7_75t_SL g153824__168280 (.A1(n_28520),
    .A2(n_4877),
    .B1(\u11_mem[2] [15]),
    .B2(n_61785),
    .Y(n_12854));
 AOI22xp5_ASAP7_75t_SL g153825__168282 (.A1(n_28520),
    .A2(n_21552),
    .B1(\u11_mem[2] [16]),
    .B2(n_61785),
    .Y(n_12856));
 AOI22xp5_ASAP7_75t_SL g153826__168281 (.A1(n_28520),
    .A2(n_4881),
    .B1(\u11_mem[2] [17]),
    .B2(n_61785),
    .Y(n_12855));
 AOI22xp5_ASAP7_75t_SL g153827__168283 (.A1(n_28520),
    .A2(n_4883),
    .B1(\u11_mem[2] [18]),
    .B2(n_61785),
    .Y(n_12857));
 AOI221xp5_ASAP7_75t_SL g153829__173944 (.A1(n_4788),
    .A2(n_28239),
    .B1(n_49131),
    .B2(n_4787),
    .C(n_4087),
    .Y(n_19688));
 AOI221xp5_ASAP7_75t_SL g153830__205422 (.A1(n_4788),
    .A2(n_56868),
    .B1(n_36107),
    .B2(n_4787),
    .C(n_4086),
    .Y(n_56870));
 AOI221xp5_ASAP7_75t_SL g153833__178097 (.A1(n_4792),
    .A2(n_43320),
    .B1(n_70649),
    .B2(n_14006),
    .C(n_24595),
    .Y(n_24596));
 AOI221xp5_ASAP7_75t_SL g153835__6131 (.A1(n_4792),
    .A2(n_31058),
    .B1(n_70649),
    .B2(n_4515),
    .C(n_4084),
    .Y(n_4794));
 AOI21xp5_ASAP7_75t_SL g153837__9945 (.A1(n_64813),
    .A2(n_5077),
    .B(n_4456),
    .Y(n_4933));
 AOI221xp5_ASAP7_75t_SL g153839__180563 (.A1(n_27372),
    .A2(n_5077),
    .B1(n_4225),
    .B2(out_slt8[19]),
    .C(n_4375),
    .Y(n_27373));
 AOI22xp33_ASAP7_75t_R g153840 (.A1(u0_slt9_r[1]),
    .A2(n_9295),
    .B1(out_slt9[2]),
    .B2(n_9345),
    .Y(n_3985));
 AOI221xp5_ASAP7_75t_SL g153841__191897 (.A1(n_1723),
    .A2(n_79196),
    .B1(n_4795),
    .B2(n_40902),
    .C(n_4083),
    .Y(n_40905));
 AOI221xp5_ASAP7_75t_SL g153842__8246 (.A1(n_1838),
    .A2(n_79196),
    .B1(n_4795),
    .B2(n_59477),
    .C(n_4082),
    .Y(n_4798));
 AOI221xp5_ASAP7_75t_SL g153843__5477 (.A1(n_31863),
    .A2(out_slt3[12]),
    .B1(n_25405),
    .B2(n_22064),
    .C(n_4359),
    .Y(n_4927));
 AOI221x1_ASAP7_75t_SL g153844__219225 (.A1(out_slt9[14]),
    .A2(n_73307),
    .B1(n_5028),
    .B2(n_13738),
    .C(n_79200),
    .Y(n_73308));
 AOI221x1_ASAP7_75t_SL g153845__200405 (.A1(n_73313),
    .A2(out_slt9[15]),
    .B1(n_5091),
    .B2(n_2603),
    .C(n_79201),
    .Y(n_50541));
 AOI22xp5_ASAP7_75t_SL g153859__4319 (.A1(n_24803),
    .A2(n_31786),
    .B1(\u10_mem[1] [8]),
    .B2(n_78621),
    .Y(n_4807));
 AOI22xp5_ASAP7_75t_SL g153862__6417 (.A1(n_24803),
    .A2(n_61243),
    .B1(\u10_mem[1] [11]),
    .B2(n_32302),
    .Y(n_4656));
 AOI22xp5_ASAP7_75t_SL g153863__2802 (.A1(n_28747),
    .A2(n_24803),
    .B1(\u10_mem[1] [12]),
    .B2(n_32302),
    .Y(n_4721));
 AOI22xp33_ASAP7_75t_SL g153864__1705 (.A1(n_17613),
    .A2(n_24803),
    .B1(\u10_mem[1] [13]),
    .B2(n_32302),
    .Y(n_4719));
 AOI22xp33_ASAP7_75t_SL g153865__5122 (.A1(n_17614),
    .A2(n_24803),
    .B1(\u10_mem[1] [14]),
    .B2(n_32302),
    .Y(n_4717));
 AOI22xp5_ASAP7_75t_SL g153866__8246 (.A1(n_24803),
    .A2(n_17615),
    .B1(n_32302),
    .B2(\u10_mem[1] [15]),
    .Y(n_4715));
 AOI22xp5_ASAP7_75t_SL g153867__7098 (.A1(n_24803),
    .A2(n_4712),
    .B1(\u10_mem[1] [16]),
    .B2(n_32302),
    .Y(n_4713));
 AOI22xp5_ASAP7_75t_SL g153868__6131 (.A1(n_24803),
    .A2(n_4710),
    .B1(\u10_mem[1] [17]),
    .B2(n_32302),
    .Y(n_4711));
 AOI22xp5_ASAP7_75t_SL g153869__167224 (.A1(n_50549),
    .A2(n_24803),
    .B1(\u10_mem[1] [18]),
    .B2(n_32302),
    .Y(n_11699));
 AOI22xp5_ASAP7_75t_SL g153870__5115 (.A1(n_24803),
    .A2(n_50551),
    .B1(\u10_mem[1] [19]),
    .B2(n_32302),
    .Y(n_4707));
 OAI211xp5_ASAP7_75t_SL g153871__223685 (.A1(n_13266),
    .A2(n_78137),
    .B(n_78139),
    .C(n_78140),
    .Y(n_78141));
 OAI211xp5_ASAP7_75t_SL g153873__167561 (.A1(n_12098),
    .A2(n_18743),
    .B(n_4048),
    .C(n_4081),
    .Y(n_12099));
 AOI22xp33_ASAP7_75t_R g153875__1705 (.A1(u1_sr[10]),
    .A2(out_le[3]),
    .B1(in_slt3[10]),
    .B2(n_5338),
    .Y(n_5281));
 AOI22xp33_ASAP7_75t_R g153876__2802 (.A1(u1_sr[10]),
    .A2(out_le[4]),
    .B1(in_slt4[10]),
    .B2(n_5341),
    .Y(n_5282));
 AOI22xp33_ASAP7_75t_R g153877__1617 (.A1(u1_sr[10]),
    .A2(out_le[5]),
    .B1(in_slt6[10]),
    .B2(n_5333),
    .Y(n_5283));
 AOI22xp33_ASAP7_75t_SL g153879__193871 (.A1(n_8112),
    .A2(n_26806),
    .B1(n_43088),
    .B2(out_slt4[0]),
    .Y(n_43096));
 AOI22xp33_ASAP7_75t_SL g153880__193867 (.A1(n_18684),
    .A2(n_26806),
    .B1(n_43088),
    .B2(out_slt4[1]),
    .Y(n_43092));
 AOI22xp33_ASAP7_75t_SL g153882__213722 (.A1(n_26098),
    .A2(n_28690),
    .B1(n_66672),
    .B2(out_slt6[1]),
    .Y(n_66681));
 AOI22xp5_ASAP7_75t_SL g153883__196657 (.A1(n_36628),
    .A2(n_4527),
    .B1(out_slt7[0]),
    .B2(n_46184),
    .Y(n_46188));
 AOI22xp33_ASAP7_75t_SL g153886__205418 (.A1(n_56868),
    .A2(n_49719),
    .B1(n_51158),
    .B2(out_slt8[1]),
    .Y(n_56869));
 AOI22xp5_ASAP7_75t_SL g153887__169189 (.A1(n_14006),
    .A2(n_4514),
    .B1(out_slt3[0]),
    .B2(n_4513),
    .Y(n_14008));
 AOI22xp33_ASAP7_75t_SL g153888__3680 (.A1(n_4515),
    .A2(n_4514),
    .B1(n_4513),
    .B2(out_slt3[1]),
    .Y(n_4516));
 AOI22xp33_ASAP7_75t_SL g153889__219219 (.A1(n_79195),
    .A2(n_40902),
    .B1(n_73301),
    .B2(out_slt9[0]),
    .Y(n_73302));
 AOI22xp33_ASAP7_75t_SL g153890__219221 (.A1(n_59477),
    .A2(n_79195),
    .B1(n_73301),
    .B2(out_slt9[1]),
    .Y(n_73303));
 OAI222xp33_ASAP7_75t_SL g153891__176455 (.A1(n_7863),
    .A2(n_66670),
    .B1(n_34479),
    .B2(n_22530),
    .C1(n_50463),
    .C2(n_19593),
    .Y(n_22532));
 AOI22xp5_ASAP7_75t_SL g153893__168312 (.A1(n_25675),
    .A2(n_12869),
    .B1(\u9_mem[2] [20]),
    .B2(n_5258),
    .Y(n_12886));
 AOI22xp5_ASAP7_75t_SL g153894__168311 (.A1(n_5185),
    .A2(n_12869),
    .B1(\u9_mem[2] [21]),
    .B2(n_5258),
    .Y(n_12885));
 AOI22xp5_ASAP7_75t_SL g153895__168310 (.A1(n_5181),
    .A2(n_12869),
    .B1(\u9_mem[2] [22]),
    .B2(n_5258),
    .Y(n_12884));
 AOI22xp5_ASAP7_75t_SL g153896__168309 (.A1(n_25673),
    .A2(n_12869),
    .B1(\u9_mem[2] [23]),
    .B2(n_5258),
    .Y(n_12883));
 AOI22xp5_ASAP7_75t_SL g153897__168308 (.A1(n_25674),
    .A2(n_12869),
    .B1(\u9_mem[2] [24]),
    .B2(n_5258),
    .Y(n_12882));
 AOI22xp5_ASAP7_75t_SL g153898__168307 (.A1(n_12869),
    .A2(n_5173),
    .B1(\u9_mem[2] [25]),
    .B2(n_5258),
    .Y(n_12881));
 AOI22xp5_ASAP7_75t_SL g153899__168306 (.A1(n_5171),
    .A2(n_12869),
    .B1(\u9_mem[2] [26]),
    .B2(n_5258),
    .Y(n_12880));
 AOI22xp5_ASAP7_75t_SL g153900__168305 (.A1(n_5177),
    .A2(n_12869),
    .B1(\u9_mem[2] [27]),
    .B2(n_5258),
    .Y(n_12879));
 AOI22xp5_ASAP7_75t_SL g153901__168297 (.A1(n_12871),
    .A2(n_25682),
    .B1(\u9_mem[2] [28]),
    .B2(n_5258),
    .Y(n_12872));
 AOI22xp5_ASAP7_75t_SL g153902__168304 (.A1(n_25679),
    .A2(n_12869),
    .B1(\u9_mem[2] [29]),
    .B2(n_5258),
    .Y(n_12878));
 AOI22xp5_ASAP7_75t_SL g153903__168303 (.A1(n_25680),
    .A2(n_12869),
    .B1(\u9_mem[2] [30]),
    .B2(n_5258),
    .Y(n_12877));
 AOI22xp5_ASAP7_75t_SL g153904__168302 (.A1(n_12869),
    .A2(n_25681),
    .B1(\u9_mem[2] [31]),
    .B2(n_5258),
    .Y(n_12876));
 AOI22xp5_ASAP7_75t_SL g153906__168272 (.A1(n_45625),
    .A2(n_4901),
    .B1(\u11_mem[2] [21]),
    .B2(n_61785),
    .Y(n_12846));
 AOI22xp5_ASAP7_75t_SL g153907__168268 (.A1(n_45625),
    .A2(n_4903),
    .B1(\u11_mem[2] [22]),
    .B2(n_61785),
    .Y(n_12842));
 AOI22xp5_ASAP7_75t_SL g153908__168265 (.A1(n_45625),
    .A2(n_4905),
    .B1(\u11_mem[2] [23]),
    .B2(n_61785),
    .Y(n_12839));
 AOI22xp5_ASAP7_75t_SL g153909__168264 (.A1(n_45625),
    .A2(n_4907),
    .B1(\u11_mem[2] [24]),
    .B2(n_61785),
    .Y(n_12838));
 AOI22xp5_ASAP7_75t_SL g153911__168274 (.A1(n_45625),
    .A2(n_4911),
    .B1(\u11_mem[2] [26]),
    .B2(n_61785),
    .Y(n_12848));
 AOI22xp5_ASAP7_75t_SL g153912__168269 (.A1(n_45625),
    .A2(n_4913),
    .B1(\u11_mem[2] [27]),
    .B2(n_61785),
    .Y(n_12843));
 AOI22xp5_ASAP7_75t_SL g153913__168273 (.A1(n_45625),
    .A2(n_4915),
    .B1(\u11_mem[2] [28]),
    .B2(n_61785),
    .Y(n_12847));
 AOI22xp5_ASAP7_75t_SL g153914__168271 (.A1(n_45625),
    .A2(n_4917),
    .B1(\u11_mem[2] [29]),
    .B2(n_61785),
    .Y(n_12845));
 AOI22xp5_ASAP7_75t_SL g153915__168275 (.A1(n_45625),
    .A2(n_4919),
    .B1(\u11_mem[2] [30]),
    .B2(n_61785),
    .Y(n_12849));
 AOI22xp5_ASAP7_75t_SL g153917__178432 (.A1(n_61242),
    .A2(n_4675),
    .B1(\u10_mem[3] [20]),
    .B2(n_35121),
    .Y(n_24984));
 AOI22xp5_ASAP7_75t_SL g153918__178455 (.A1(n_61242),
    .A2(n_4673),
    .B1(\u10_mem[3] [21]),
    .B2(n_61244),
    .Y(n_25008));
 AOI22xp5_ASAP7_75t_SL g153919__178452 (.A1(n_61242),
    .A2(n_4671),
    .B1(\u10_mem[3] [22]),
    .B2(n_61244),
    .Y(n_25005));
 AOI22xp5_ASAP7_75t_SL g153920__187221 (.A1(n_61242),
    .A2(n_35120),
    .B1(n_35121),
    .B2(\u10_mem[3] [23]),
    .Y(n_35122));
 AOI22xp5_ASAP7_75t_SL g153921__178429 (.A1(n_61242),
    .A2(n_4667),
    .B1(\u10_mem[3] [24]),
    .B2(n_35121),
    .Y(n_24981));
 AOI22xp5_ASAP7_75t_SL g153922__178454 (.A1(n_61242),
    .A2(n_4665),
    .B1(\u10_mem[3] [25]),
    .B2(n_61244),
    .Y(n_25007));
 AOI22xp5_ASAP7_75t_SL g153923__178453 (.A1(n_61242),
    .A2(n_4663),
    .B1(\u10_mem[3] [26]),
    .B2(n_61244),
    .Y(n_25006));
 AOI22xp5_ASAP7_75t_SL g153924__178430 (.A1(n_61242),
    .A2(n_4661),
    .B1(\u10_mem[3] [27]),
    .B2(n_35121),
    .Y(n_24982));
 AOI22xp5_ASAP7_75t_SL g153925__178457 (.A1(n_61242),
    .A2(n_4695),
    .B1(\u10_mem[3] [28]),
    .B2(n_61244),
    .Y(n_25010));
 AOI22xp5_ASAP7_75t_SL g153926__178427 (.A1(n_61242),
    .A2(n_4693),
    .B1(\u10_mem[3] [29]),
    .B2(n_35121),
    .Y(n_24979));
 AOI22xp5_ASAP7_75t_SL g153927__178456 (.A1(n_61242),
    .A2(n_4691),
    .B1(\u10_mem[3] [30]),
    .B2(n_61244),
    .Y(n_25009));
 AOI22xp5_ASAP7_75t_SL g153928__178428 (.A1(n_61242),
    .A2(n_4689),
    .B1(\u10_mem[3] [31]),
    .B2(n_35121),
    .Y(n_24980));
 AOI22xp5_ASAP7_75t_SL g153929__5526 (.A1(n_25675),
    .A2(n_31720),
    .B1(\u9_mem[0] [20]),
    .B2(n_46587),
    .Y(n_4876));
 AOI22xp5_ASAP7_75t_SL g153930__3680 (.A1(n_5185),
    .A2(n_31720),
    .B1(\u9_mem[0] [21]),
    .B2(n_46587),
    .Y(n_4873));
 AOI22xp5_ASAP7_75t_SL g153931__1617 (.A1(n_5181),
    .A2(n_31720),
    .B1(\u9_mem[0] [22]),
    .B2(n_46587),
    .Y(n_4872));
 AOI22xp5_ASAP7_75t_SL g153932__2802 (.A1(n_25673),
    .A2(n_31720),
    .B1(\u9_mem[0] [23]),
    .B2(n_46587),
    .Y(n_4871));
 AOI22xp5_ASAP7_75t_SL g153933__5122 (.A1(n_25674),
    .A2(n_31720),
    .B1(\u9_mem[0] [24]),
    .B2(n_46587),
    .Y(n_4868));
 AOI22xp5_ASAP7_75t_SL g153934__8246 (.A1(n_31720),
    .A2(n_5173),
    .B1(\u9_mem[0] [25]),
    .B2(n_46587),
    .Y(n_4867));
 AOI22xp5_ASAP7_75t_SL g153935__6131 (.A1(n_5171),
    .A2(n_31720),
    .B1(\u9_mem[0] [26]),
    .B2(n_46587),
    .Y(n_4865));
 AOI22xp5_ASAP7_75t_SL g153936__1881 (.A1(n_5177),
    .A2(n_31720),
    .B1(\u9_mem[0] [27]),
    .B2(n_46587),
    .Y(n_4864));
 AOI22xp5_ASAP7_75t_SL g153937__7482 (.A1(n_25682),
    .A2(n_31720),
    .B1(\u9_mem[0] [28]),
    .B2(n_46587),
    .Y(n_4862));
 AOI22xp5_ASAP7_75t_SL g153938__4733 (.A1(n_25679),
    .A2(n_31720),
    .B1(\u9_mem[0] [29]),
    .B2(n_46587),
    .Y(n_4861));
 AOI22xp5_ASAP7_75t_SL g153939__9315 (.A1(n_25680),
    .A2(n_31720),
    .B1(\u9_mem[0] [30]),
    .B2(n_46587),
    .Y(n_4859));
 AOI22xp5_ASAP7_75t_SL g153940__9945 (.A1(n_25681),
    .A2(n_31720),
    .B1(\u9_mem[0] [31]),
    .B2(n_46587),
    .Y(n_4858));
 AOI22xp5_ASAP7_75t_SL g153941__182091 (.A1(n_4899),
    .A2(n_29011),
    .B1(\u11_mem[0] [20]),
    .B2(n_4784),
    .Y(n_29030));
 AOI22xp5_ASAP7_75t_SL g153942__182098 (.A1(n_4901),
    .A2(n_29011),
    .B1(\u11_mem[0] [21]),
    .B2(n_4784),
    .Y(n_29037));
 AOI22xp5_ASAP7_75t_SL g153943__182099 (.A1(n_4903),
    .A2(n_29011),
    .B1(\u11_mem[0] [22]),
    .B2(n_4784),
    .Y(n_29038));
 AOI22xp5_ASAP7_75t_SL g153944__182088 (.A1(n_29011),
    .A2(n_4905),
    .B1(\u11_mem[0] [23]),
    .B2(n_4784),
    .Y(n_29027));
 AOI22xp5_ASAP7_75t_SL g153945__182096 (.A1(n_4907),
    .A2(n_29011),
    .B1(\u11_mem[0] [24]),
    .B2(n_4784),
    .Y(n_29035));
 AOI22xp5_ASAP7_75t_SL g153946__182093 (.A1(n_4909),
    .A2(n_29011),
    .B1(\u11_mem[0] [25]),
    .B2(n_4784),
    .Y(n_29032));
 AOI22xp5_ASAP7_75t_SL g153947__182090 (.A1(n_4911),
    .A2(n_29011),
    .B1(\u11_mem[0] [26]),
    .B2(n_4784),
    .Y(n_29029));
 AOI22xp5_ASAP7_75t_SL g153948__182101 (.A1(n_4913),
    .A2(n_29011),
    .B1(\u11_mem[0] [27]),
    .B2(n_4784),
    .Y(n_29040));
 AOI22xp5_ASAP7_75t_SL g153949__182092 (.A1(n_4915),
    .A2(n_29011),
    .B1(\u11_mem[0] [28]),
    .B2(n_4784),
    .Y(n_29031));
 AOI22xp5_ASAP7_75t_SL g153950__182087 (.A1(n_4917),
    .A2(n_29011),
    .B1(\u11_mem[0] [29]),
    .B2(n_4784),
    .Y(n_29026));
 AOI22xp5_ASAP7_75t_SL g153951__182100 (.A1(n_4919),
    .A2(n_29011),
    .B1(\u11_mem[0] [30]),
    .B2(n_4784),
    .Y(n_29039));
 AOI22xp5_ASAP7_75t_SL g153952__182095 (.A1(n_30483),
    .A2(n_29011),
    .B1(\u11_mem[0] [31]),
    .B2(n_4784),
    .Y(n_29034));
 AOI22xp5_ASAP7_75t_SL g153954__1881 (.A1(n_4673),
    .A2(n_24803),
    .B1(\u10_mem[1] [21]),
    .B2(n_32302),
    .Y(n_4674));
 AOI22xp5_ASAP7_75t_SL g153956__7482 (.A1(n_35120),
    .A2(n_24803),
    .B1(\u10_mem[1] [23]),
    .B2(n_32302),
    .Y(n_4670));
 AOI22xp5_ASAP7_75t_SL g153959__9315 (.A1(n_24803),
    .A2(n_4663),
    .B1(\u10_mem[1] [26]),
    .B2(n_32302),
    .Y(n_4664));
 AOI22xp5_ASAP7_75t_SL g153960__9945 (.A1(n_24803),
    .A2(n_4661),
    .B1(\u10_mem[1] [27]),
    .B2(n_32302),
    .Y(n_4662));
 AOI22xp5_ASAP7_75t_SL g153963__1666 (.A1(n_24803),
    .A2(n_4691),
    .B1(\u10_mem[1] [30]),
    .B2(n_32302),
    .Y(n_4658));
 AOI22xp5_ASAP7_75t_SL g153964__7410 (.A1(n_24803),
    .A2(n_4689),
    .B1(\u10_mem[1] [31]),
    .B2(n_32302),
    .Y(n_4657));
 OAI221xp5_ASAP7_75t_SL g153971__218177 (.A1(n_3996),
    .A2(n_72059),
    .B1(n_72060),
    .B2(n_79204),
    .C(n_51479),
    .Y(n_72061));
 OAI221xp5_ASAP7_75t_SL g153972__182369 (.A1(n_17616),
    .A2(n_6242),
    .B1(n_20317),
    .B2(n_29312),
    .C(n_33796),
    .Y(n_29313));
 OAI221xp5_ASAP7_75t_SL g153973__5526 (.A1(n_6115),
    .A2(n_3999),
    .B1(n_4645),
    .B2(n_2458),
    .C(n_48426),
    .Y(n_4646));
 OAI221xp5_ASAP7_75t_SL g153974__6783 (.A1(n_42249),
    .A2(n_7656),
    .B1(n_52770),
    .B2(n_2462),
    .C(n_51036),
    .Y(n_4644));
 AOI322xp5_ASAP7_75t_SL g153975__213703 (.A1(n_34475),
    .A2(n_725),
    .A3(n_37311),
    .B1(n_56850),
    .B2(n_64847),
    .C1(u5_rp[3]),
    .C2(n_66659),
    .Y(n_66661));
 AOI22xp5_ASAP7_75t_SL g153976__168300 (.A1(n_12869),
    .A2(n_25677),
    .B1(\u9_mem[2] [16]),
    .B2(n_5258),
    .Y(n_12874));
 INVxp33_ASAP7_75t_R g153977 (.A(u1_sr[11]),
    .Y(n_5287));
 AOI22xp5_ASAP7_75t_SL g153978__7098 (.A1(n_46478),
    .A2(n_48456),
    .B1(\u10_mem[0] [1]),
    .B2(n_46477),
    .Y(n_4502));
 O2A1O1Ixp33_ASAP7_75t_SL g153979__173338 (.A1(n_19045),
    .A2(n_47768),
    .B(n_19046),
    .C(n_17686),
    .Y(n_19047));
 AOI22xp5_ASAP7_75t_SL g153985__1881 (.A1(n_50555),
    .A2(n_46478),
    .B1(\u10_mem[0] [4]),
    .B2(n_46477),
    .Y(n_4500));
 AOI22xp5_ASAP7_75t_SL g153986__5115 (.A1(n_35392),
    .A2(n_46478),
    .B1(\u10_mem[0] [3]),
    .B2(n_46477),
    .Y(n_4498));
 AOI22xp33_ASAP7_75t_R g153994__8246 (.A1(out_le[0]),
    .A2(u1_sr[9]),
    .B1(in_slt0[9]),
    .B2(n_5296),
    .Y(n_5278));
 AOI22xp33_ASAP7_75t_R g153995__7098 (.A1(u1_sr[9]),
    .A2(out_le[2]),
    .B1(in_slt2[9]),
    .B2(n_5336),
    .Y(n_5277));
 A2O1A1Ixp33_ASAP7_75t_SL g153996__4733 (.A1(n_31872),
    .A2(n_2685),
    .B(n_4485),
    .C(n_4258),
    .Y(n_4495));
 A2O1A1Ixp33_ASAP7_75t_SL g153997__189853 (.A1(n_43205),
    .A2(n_64713),
    .B(n_38374),
    .C(n_66674),
    .Y(n_38380));
 A2O1A1Ixp33_ASAP7_75t_SL g153998__189854 (.A1(n_4332),
    .A2(n_2486),
    .B(n_38374),
    .C(n_66673),
    .Y(n_38381));
 AOI22xp5_ASAP7_75t_SL g154 (.A1(\u8_mem[3] [4]),
    .A2(n_78273),
    .B1(\u8_mem[1] [4]),
    .B2(n_78274),
    .Y(n_48972));
 A2O1A1Ixp33_ASAP7_75t_SL g154000__189844 (.A1(n_21027),
    .A2(n_31869),
    .B(n_38364),
    .C(n_66664),
    .Y(n_38370));
 AOI22xp5_ASAP7_75t_SL g154002__2346 (.A1(n_46478),
    .A2(n_40956),
    .B1(\u10_mem[0] [0]),
    .B2(n_46477),
    .Y(n_4489));
 AOI22xp5_ASAP7_75t_SL g154003__1666 (.A1(n_46478),
    .A2(n_62614),
    .B1(\u10_mem[0] [2]),
    .B2(n_46477),
    .Y(n_4488));
 AND3x4_ASAP7_75t_SL g154062__178195 (.A(n_21261),
    .B(n_203),
    .C(u9_wp[1]),
    .Y(n_24735));
 OR2x6_ASAP7_75t_SL g154063__174765 (.A(n_28952),
    .B(n_225),
    .Y(n_20594));
 OR2x6_ASAP7_75t_SL g154063__9945_dup174766 (.A(n_28952),
    .B(n_225),
    .Y(n_20595));
 OR2x6_ASAP7_75t_SL g154065__175620 (.A(n_28952),
    .B(n_29003),
    .Y(n_21553));
 OR2x6_ASAP7_75t_SL g154065__9315_dup174764 (.A(n_28952),
    .B(n_29003),
    .Y(n_20593));
 AND3x4_ASAP7_75t_SL g154068__178190 (.A(n_259),
    .B(n_21261),
    .C(u9_wp[1]),
    .Y(n_24734));
 AOI22xp5_ASAP7_75t_SL g154069__2398 (.A1(n_46478),
    .A2(n_50553),
    .B1(\u10_mem[0] [5]),
    .B2(n_46477),
    .Y(n_4483));
 AOI22xp33_ASAP7_75t_SL g154071__6260 (.A1(n_46478),
    .A2(n_50552),
    .B1(\u10_mem[0] [7]),
    .B2(n_46477),
    .Y(n_4481));
 AOI22xp33_ASAP7_75t_SL g154077__1617 (.A1(n_46478),
    .A2(n_17613),
    .B1(n_46477),
    .B2(\u10_mem[0] [13]),
    .Y(n_4475));
 AOI22xp33_ASAP7_75t_SL g154078__2802 (.A1(n_17614),
    .A2(n_46478),
    .B1(\u10_mem[0] [14]),
    .B2(n_46477),
    .Y(n_4474));
 AOI22xp33_ASAP7_75t_SL g154079__1705 (.A1(n_17615),
    .A2(n_46478),
    .B1(\u10_mem[0] [15]),
    .B2(n_46477),
    .Y(n_4473));
 AOI22xp5_ASAP7_75t_SL g154080__5122 (.A1(n_46478),
    .A2(n_4712),
    .B1(\u10_mem[0] [16]),
    .B2(n_46477),
    .Y(n_4472));
 AOI22xp5_ASAP7_75t_SL g154081__7098 (.A1(n_46478),
    .A2(n_4710),
    .B1(\u10_mem[0] [17]),
    .B2(n_46477),
    .Y(n_4470));
 AOI22xp5_ASAP7_75t_SL g154082__167222 (.A1(n_50549),
    .A2(n_46478),
    .B1(\u10_mem[0] [18]),
    .B2(n_46477),
    .Y(n_11697));
 AOI22xp5_ASAP7_75t_SL g154085__198354 (.A1(n_48456),
    .A2(n_36975),
    .B1(\u10_mem[2] [1]),
    .B2(n_48146),
    .Y(n_48159));
 AOI22xp5_ASAP7_75t_SL g154087__198359 (.A1(n_35392),
    .A2(n_36971),
    .B1(\u10_mem[2] [3]),
    .B2(n_48146),
    .Y(n_48164));
 AOI22xp33_ASAP7_75t_SL g154088__198370 (.A1(n_50555),
    .A2(n_36975),
    .B1(\u10_mem[2] [4]),
    .B2(n_48153),
    .Y(n_48175));
 AOI22xp33_ASAP7_75t_SL g154089__198371 (.A1(n_50553),
    .A2(n_36971),
    .B1(\u10_mem[2] [5]),
    .B2(n_48153),
    .Y(n_48176));
 AOI22xp33_ASAP7_75t_SL g154091__198355 (.A1(n_36971),
    .A2(n_50552),
    .B1(n_48146),
    .B2(\u10_mem[2] [7]),
    .Y(n_48160));
 AOI22xp5_ASAP7_75t_SL g154092__198348 (.A1(n_31786),
    .A2(n_36975),
    .B1(\u10_mem[2] [8]),
    .B2(n_48153),
    .Y(n_48154));
 AOI22xp5_ASAP7_75t_SL g154093__198350 (.A1(n_18707),
    .A2(n_36975),
    .B1(\u10_mem[2] [9]),
    .B2(n_48146),
    .Y(n_48155));
 AOI22xp33_ASAP7_75t_SL g154094__198366 (.A1(n_36971),
    .A2(n_46479),
    .B1(\u10_mem[2] [10]),
    .B2(n_48153),
    .Y(n_48171));
 AOI22xp5_ASAP7_75t_SL g154095__198358 (.A1(n_36971),
    .A2(n_61243),
    .B1(\u10_mem[2] [11]),
    .B2(n_48146),
    .Y(n_48163));
 AOI22xp5_ASAP7_75t_SL g154096__198353 (.A1(n_28747),
    .A2(n_36975),
    .B1(\u10_mem[2] [12]),
    .B2(n_48146),
    .Y(n_48158));
 AOI22xp33_ASAP7_75t_SL g154097__198367 (.A1(n_36971),
    .A2(n_17613),
    .B1(n_48153),
    .B2(\u10_mem[2] [13]),
    .Y(n_48172));
 A2O1A1Ixp33_ASAP7_75t_SL g154098__181547 (.A1(n_37367),
    .A2(n_2362),
    .B(n_48223),
    .C(n_46189),
    .Y(n_28412));
 AOI22xp33_ASAP7_75t_SL g154099__198356 (.A1(n_36971),
    .A2(n_17614),
    .B1(n_48146),
    .B2(\u10_mem[2] [14]),
    .Y(n_48161));
 AOI22xp33_ASAP7_75t_SL g154100__198368 (.A1(n_36971),
    .A2(n_17615),
    .B1(n_48153),
    .B2(\u10_mem[2] [15]),
    .Y(n_48173));
 AOI22xp5_ASAP7_75t_SL g154101__198351 (.A1(n_4712),
    .A2(n_36975),
    .B1(\u10_mem[2] [16]),
    .B2(n_48146),
    .Y(n_48156));
 AOI22xp5_ASAP7_75t_SL g154102__198352 (.A1(n_4710),
    .A2(n_36975),
    .B1(\u10_mem[2] [17]),
    .B2(n_48146),
    .Y(n_48157));
 AOI22xp33_ASAP7_75t_SL g154103__198365 (.A1(n_50549),
    .A2(n_36971),
    .B1(\u10_mem[2] [18]),
    .B2(n_48153),
    .Y(n_48170));
 AOI22xp33_ASAP7_75t_SL g154104__198357 (.A1(n_36971),
    .A2(n_50551),
    .B1(n_48146),
    .B2(\u10_mem[2] [19]),
    .Y(n_48162));
 A2O1A1Ixp33_ASAP7_75t_SL g154106__6260 (.A1(n_7754),
    .A2(n_7806),
    .B(n_64852),
    .C(n_43086),
    .Y(n_4617));
 A2O1A1Ixp33_ASAP7_75t_L g154108__4733 (.A1(n_34434),
    .A2(n_2508),
    .B(n_27225),
    .C(n_42252),
    .Y(n_4464));
 A2O1A1Ixp33_ASAP7_75t_L g154109__6161 (.A1(n_4448),
    .A2(n_2511),
    .B(n_27225),
    .C(n_42254),
    .Y(n_4462));
 A2O1A1Ixp33_ASAP7_75t_SL g154110__8428 (.A1(n_1850),
    .A2(n_2578),
    .B(n_64852),
    .C(n_4254),
    .Y(n_4614));
 A2O1A1Ixp33_ASAP7_75t_L g154111__9315 (.A1(n_2498),
    .A2(n_2540),
    .B(n_27225),
    .C(n_42251),
    .Y(n_4461));
 A2O1A1Ixp33_ASAP7_75t_L g154112__9945 (.A1(n_15101),
    .A2(n_2503),
    .B(n_27225),
    .C(n_4186),
    .Y(n_4460));
 A2O1A1Ixp33_ASAP7_75t_SL g154114__200937 (.A1(n_56060),
    .A2(n_1872),
    .B(n_27225),
    .C(n_51159),
    .Y(n_51160));
 A2O1A1Ixp33_ASAP7_75t_SL g154115__1666 (.A1(n_1845),
    .A2(n_2500),
    .B(n_27225),
    .C(n_42255),
    .Y(n_4457));
 A2O1A1Ixp33_ASAP7_75t_SL g154116__7410 (.A1(n_1736),
    .A2(n_2403),
    .B(n_27225),
    .C(n_42256),
    .Y(n_4456));
 A2O1A1Ixp33_ASAP7_75t_SL g154117__8246 (.A1(n_41492),
    .A2(n_2401),
    .B(n_27225),
    .C(n_42257),
    .Y(n_4471));
 A2O1A1Ixp33_ASAP7_75t_SL g154118__5477 (.A1(n_4381),
    .A2(n_49499),
    .B(n_4485),
    .C(n_4180),
    .Y(n_4484));
 A2O1A1Ixp33_ASAP7_75t_SL g154119__6417 (.A1(n_4377),
    .A2(n_46230),
    .B(n_4485),
    .C(n_4179),
    .Y(n_4486));
 A2O1A1Ixp33_ASAP7_75t_SL g154120__4319 (.A1(n_57041),
    .A2(n_2444),
    .B(n_4524),
    .C(n_73304),
    .Y(n_4525));
 A2O1A1Ixp33_ASAP7_75t_SL g154121__171814 (.A1(n_17617),
    .A2(n_2446),
    .B(n_4524),
    .C(n_73305),
    .Y(n_17184));
 XNOR2xp5_ASAP7_75t_SL g154122__6417 (.A(n_402),
    .B(n_3991),
    .Y(n_4232));
 AOI22xp33_ASAP7_75t_SL g154123__175580 (.A1(n_21513),
    .A2(crac_wr),
    .B1(u15_crac_we_r),
    .B2(n_21514),
    .Y(n_21515));
 AOI21xp5_ASAP7_75t_SL g154125 (.A1(n_28880),
    .A2(u16_u7_dma_req_r1),
    .B(n_487),
    .Y(n_4161));
 AOI21xp5_ASAP7_75t_SL g154126 (.A1(n_18873),
    .A2(u16_u8_dma_req_r1),
    .B(n_391),
    .Y(n_4162));
 AOI22xp33_ASAP7_75t_R g154127__6131 (.A1(u1_sr[9]),
    .A2(n_10735),
    .B1(in_slt3[9]),
    .B2(n_10761),
    .Y(n_5276));
 AOI22xp33_ASAP7_75t_R g154128__1881 (.A1(u1_sr[9]),
    .A2(n_10709),
    .B1(in_slt4[9]),
    .B2(n_10787),
    .Y(n_5275));
 AOI22xp33_ASAP7_75t_R g154129__5115 (.A1(u1_sr[9]),
    .A2(n_10839),
    .B1(in_slt6[9]),
    .B2(n_10813),
    .Y(n_5274));
 AOI22xp5_ASAP7_75t_SL g154130__198343 (.A1(n_4675),
    .A2(n_36975),
    .B1(\u10_mem[2] [20]),
    .B2(n_48146),
    .Y(n_48148));
 AOI22xp5_ASAP7_75t_SL g154131__198347 (.A1(n_4673),
    .A2(n_36971),
    .B1(\u10_mem[2] [21]),
    .B2(n_48146),
    .Y(n_48152));
 AOI22xp5_ASAP7_75t_SL g154132__198345 (.A1(n_4671),
    .A2(n_36971),
    .B1(\u10_mem[2] [22]),
    .B2(n_48146),
    .Y(n_48150));
 AOI22xp5_ASAP7_75t_SL g154133__198344 (.A1(n_35120),
    .A2(n_36971),
    .B1(\u10_mem[2] [23]),
    .B2(n_48146),
    .Y(n_48149));
 AOI22xp5_ASAP7_75t_SL g154135__198360 (.A1(n_4665),
    .A2(n_36975),
    .B1(\u10_mem[2] [25]),
    .B2(n_48146),
    .Y(n_48165));
 AOI22xp5_ASAP7_75t_SL g154136__198361 (.A1(n_4663),
    .A2(n_36971),
    .B1(\u10_mem[2] [26]),
    .B2(n_48146),
    .Y(n_48166));
 AOI22xp5_ASAP7_75t_SL g154137__198363 (.A1(n_4661),
    .A2(n_36975),
    .B1(\u10_mem[2] [27]),
    .B2(n_48146),
    .Y(n_48168));
 AOI22xp5_ASAP7_75t_SL g154138__198364 (.A1(n_36975),
    .A2(n_4695),
    .B1(\u10_mem[2] [28]),
    .B2(n_48146),
    .Y(n_48169));
 AOI22xp5_ASAP7_75t_SL g154139__198340 (.A1(n_36975),
    .A2(n_4693),
    .B1(\u10_mem[2] [29]),
    .B2(n_48146),
    .Y(n_48147));
 AOI22xp5_ASAP7_75t_SL g154140__198346 (.A1(n_4691),
    .A2(n_36971),
    .B1(\u10_mem[2] [30]),
    .B2(n_48146),
    .Y(n_48151));
 AOI22xp5_ASAP7_75t_SL g154141__198362 (.A1(n_4689),
    .A2(n_36971),
    .B1(\u10_mem[2] [31]),
    .B2(n_48146),
    .Y(n_48167));
 AOI22xp5_ASAP7_75t_SL g154142__6417 (.A1(n_4675),
    .A2(n_46478),
    .B1(\u10_mem[0] [20]),
    .B2(n_46477),
    .Y(n_4588));
 AOI22xp5_ASAP7_75t_SL g154143__6131 (.A1(n_4673),
    .A2(n_46478),
    .B1(\u10_mem[0] [21]),
    .B2(n_46477),
    .Y(n_4604));
 AOI22xp5_ASAP7_75t_SL g154144__1881 (.A1(n_4671),
    .A2(n_46478),
    .B1(\u10_mem[0] [22]),
    .B2(n_46477),
    .Y(n_4603));
 AOI22xp5_ASAP7_75t_SL g154145__5115 (.A1(n_35120),
    .A2(n_46478),
    .B1(\u10_mem[0] [23]),
    .B2(n_46477),
    .Y(n_4600));
 AOI22xp5_ASAP7_75t_SL g154146__7482 (.A1(n_4667),
    .A2(n_46478),
    .B1(\u10_mem[0] [24]),
    .B2(n_46477),
    .Y(n_4599));
 AOI22xp5_ASAP7_75t_SL g154147__4733 (.A1(n_4665),
    .A2(n_46478),
    .B1(\u10_mem[0] [25]),
    .B2(n_46477),
    .Y(n_4598));
 AOI22xp5_ASAP7_75t_SL g154148__6161 (.A1(n_4663),
    .A2(n_46478),
    .B1(\u10_mem[0] [26]),
    .B2(n_46477),
    .Y(n_4597));
 AOI22xp5_ASAP7_75t_SL g154149__9315 (.A1(n_4661),
    .A2(n_46478),
    .B1(\u10_mem[0] [27]),
    .B2(n_46477),
    .Y(n_4596));
 AOI22xp5_ASAP7_75t_SL g154150__9945 (.A1(n_4695),
    .A2(n_46478),
    .B1(\u10_mem[0] [28]),
    .B2(n_46477),
    .Y(n_4595));
 AOI22xp5_ASAP7_75t_SL g154151__2883 (.A1(n_46478),
    .A2(n_4693),
    .B1(\u10_mem[0] [29]),
    .B2(n_46477),
    .Y(n_4594));
 AOI22xp5_ASAP7_75t_SL g154152__2346 (.A1(n_4691),
    .A2(n_46478),
    .B1(\u10_mem[0] [30]),
    .B2(n_46477),
    .Y(n_4593));
 AOI22xp5_ASAP7_75t_SL g154153__1666 (.A1(n_4689),
    .A2(n_46478),
    .B1(\u10_mem[0] [31]),
    .B2(n_46477),
    .Y(n_4592));
 AOI21xp5_ASAP7_75t_SL g154154__7410 (.A1(n_4202),
    .A2(u15_crac_rd),
    .B(n_460),
    .Y(n_4591));
 INVxp33_ASAP7_75t_R g154157 (.A(u1_sr[10]),
    .Y(n_5280));
 NAND2xp33_ASAP7_75t_SL g154171__185111 (.A(n_32582),
    .B(n_36012),
    .Y(n_32583));
 NOR2xp33_ASAP7_75t_SL g154184__193872 (.A(n_43088),
    .B(n_7803),
    .Y(n_43097));
 NOR2xp33_ASAP7_75t_SL g154186__6783 (.A(n_64102),
    .B(n_42248),
    .Y(n_4443));
 NOR2xp33_ASAP7_75t_SL g154187__4733 (.A(n_46182),
    .B(n_12100),
    .Y(n_4312));
 NOR2xp33_ASAP7_75t_SL g154189__2802 (.A(n_73300),
    .B(n_13269),
    .Y(n_4439));
 NAND2xp33_ASAP7_75t_R g154190 (.A(n_6144),
    .B(n_42248),
    .Y(n_4098));
 NAND2xp33_ASAP7_75t_L g154191 (.A(n_18743),
    .B(n_46182),
    .Y(n_4081));
 NAND2xp5_ASAP7_75t_L g154200__6783 (.A(out_slt3[16]),
    .B(n_4513),
    .Y(n_4258));
 AND2x2_ASAP7_75t_SL g154206 (.A(out_slt7[2]),
    .B(n_46182),
    .Y(n_4092));
 AND2x2_ASAP7_75t_L g154215 (.A(out_slt8[2]),
    .B(n_42248),
    .Y(n_4087));
 AND2x2_ASAP7_75t_L g154216 (.A(out_slt8[3]),
    .B(n_42248),
    .Y(n_4086));
 NAND2xp5_ASAP7_75t_L g154219__2802 (.A(out_slt4[16]),
    .B(n_4253),
    .Y(n_4254));
 NAND2xp5_ASAP7_75t_L g154221 (.A(out_slt8[11]),
    .B(n_51158),
    .Y(n_4186));
 AND2x2_ASAP7_75t_SL g154223 (.A(out_slt3[3]),
    .B(n_24594),
    .Y(n_4084));
 NAND2xp5_ASAP7_75t_R g154228 (.A(out_slt3[8]),
    .B(n_5024),
    .Y(n_4180));
 NAND2xp5_ASAP7_75t_R g154229 (.A(out_slt3[9]),
    .B(n_5024),
    .Y(n_4179));
 AND2x2_ASAP7_75t_L g154230 (.A(out_slt9[2]),
    .B(n_73300),
    .Y(n_4083));
 AND2x2_ASAP7_75t_L g154231 (.A(out_slt9[3]),
    .B(n_73300),
    .Y(n_4082));
 NAND2xp5_ASAP7_75t_R g154233__219223 (.A(n_73301),
    .B(out_slt9[9]),
    .Y(n_73305));
 NOR3xp33_ASAP7_75t_SL g154241 (.A(n_4117),
    .B(n_6138),
    .C(n_4027),
    .Y(n_4527));
 NOR3xp33_ASAP7_75t_SL g154244 (.A(n_4028),
    .B(n_29310),
    .C(n_4114),
    .Y(n_4514));
 NAND2xp5_ASAP7_75t_SL g154249 (.A(n_21784),
    .B(n_21874),
    .Y(n_4078));
 OR2x6_ASAP7_75t_SL g154290__179919_dup (.A(n_32299),
    .B(n_32300),
    .Y(n_32302));
 AOI21xp33_ASAP7_75t_SL g154305__182132 (.A1(n_29074),
    .A2(u11_din_tmp1[15]),
    .B(n_29076),
    .Y(n_29077));
 AOI21xp33_ASAP7_75t_SL g154306__182151 (.A1(n_29074),
    .A2(u11_din_tmp1[14]),
    .B(n_29092),
    .Y(n_29093));
 AOI21xp33_ASAP7_75t_SL g154307__182161 (.A1(n_29074),
    .A2(u11_din_tmp1[13]),
    .B(n_29102),
    .Y(n_29103));
 AOI21xp33_ASAP7_75t_SL g154308__182153 (.A1(n_29074),
    .A2(u11_din_tmp1[12]),
    .B(n_29094),
    .Y(n_29095));
 AOI21xp33_ASAP7_75t_SL g154309__182163 (.A1(n_29074),
    .A2(u11_din_tmp1[11]),
    .B(n_29104),
    .Y(n_29105));
 AOI21xp33_ASAP7_75t_SL g154310__182141 (.A1(n_29074),
    .A2(u11_din_tmp1[10]),
    .B(n_29082),
    .Y(n_29083));
 AOI21xp33_ASAP7_75t_SL g154311 (.A1(n_12119),
    .A2(n_3908),
    .B(ic1_int_set[2]),
    .Y(n_4077));
 AOI21xp33_ASAP7_75t_SL g154313__182139 (.A1(n_36289),
    .A2(u11_din_tmp1[9]),
    .B(n_29080),
    .Y(n_29081));
 OR5x1_ASAP7_75t_SL g154314__9315 (.A(n_13420),
    .B(n_4542),
    .C(n_532),
    .D(n_24737),
    .E(u9_wp[3]),
    .Y(n_4544));
 AOI21xp33_ASAP7_75t_SL g154315__182159 (.A1(n_29074),
    .A2(u11_din_tmp1[8]),
    .B(n_29100),
    .Y(n_29101));
 OR5x1_ASAP7_75t_SL g154316__3680 (.A(n_23286),
    .B(n_4390),
    .C(n_543),
    .D(n_28954),
    .E(u11_wp[3]),
    .Y(n_4392));
 OAI21xp5_ASAP7_75t_SL g154317__201203 (.A1(n_51478),
    .A2(n_7335),
    .B(n_13269),
    .Y(n_51479));
 OAI21xp33_ASAP7_75t_SL g154318__186128 (.A1(n_7408),
    .A2(n_33795),
    .B(n_21507),
    .Y(n_33796));
 OAI21xp33_ASAP7_75t_SL g154319__198592 (.A1(n_48425),
    .A2(n_11874),
    .B(n_12100),
    .Y(n_48426));
 OAI21xp33_ASAP7_75t_SL g154320__200834 (.A1(n_51035),
    .A2(n_6299),
    .B(n_64102),
    .Y(n_51036));
 O2A1O1Ixp33_ASAP7_75t_SL g154321__6260 (.A1(n_31872),
    .A2(n_2524),
    .B(n_66198),
    .C(n_4485),
    .Y(n_4401));
 O2A1O1Ixp33_ASAP7_75t_L g154322__2398 (.A1(n_5674),
    .A2(n_2524),
    .B(n_4346),
    .C(n_4485),
    .Y(n_4404));
 O2A1O1Ixp33_ASAP7_75t_SL g154323__5477 (.A1(n_2524),
    .A2(n_4405),
    .B(n_5674),
    .C(n_4485),
    .Y(n_4407));
 AOI21xp33_ASAP7_75t_L g154324__6417 (.A1(n_7571),
    .A2(n_28893),
    .B(n_4485),
    .Y(n_4408));
 AOI21xp33_ASAP7_75t_L g154325__7410 (.A1(n_4405),
    .A2(n_20760),
    .B(n_4485),
    .Y(n_4409));
 AOI21xp33_ASAP7_75t_L g154326__1666 (.A1(n_2375),
    .A2(n_36771),
    .B(n_48223),
    .Y(n_4410));
 O2A1O1Ixp33_ASAP7_75t_L g154328__2883 (.A1(n_6122),
    .A2(n_37367),
    .B(n_36770),
    .C(n_48223),
    .Y(n_4413));
 O2A1O1Ixp33_ASAP7_75t_L g154329__9945 (.A1(n_6122),
    .A2(n_34837),
    .B(n_1742),
    .C(n_48223),
    .Y(n_4415));
 O2A1O1Ixp33_ASAP7_75t_SL g154330__9315 (.A1(n_6122),
    .A2(n_4416),
    .B(n_1853),
    .C(n_48223),
    .Y(n_4418));
 O2A1O1Ixp33_ASAP7_75t_SL g154331__176675 (.A1(n_22839),
    .A2(n_6122),
    .B(n_22841),
    .C(n_48223),
    .Y(n_22842));
 O2A1O1Ixp33_ASAP7_75t_SL g154332__4733 (.A1(n_4422),
    .A2(n_6122),
    .B(n_4416),
    .C(n_48223),
    .Y(n_4423));
 O2A1O1Ixp33_ASAP7_75t_SL g154333__7482 (.A1(n_6122),
    .A2(n_4424),
    .B(n_22839),
    .C(n_48223),
    .Y(n_4425));
 O2A1O1Ixp33_ASAP7_75t_SL g154334__5115 (.A1(n_6122),
    .A2(n_4426),
    .B(n_4422),
    .C(n_48223),
    .Y(n_4427));
 O2A1O1Ixp33_ASAP7_75t_SL g154335__1881 (.A1(n_6122),
    .A2(n_4428),
    .B(n_4424),
    .C(n_48223),
    .Y(n_4430));
 O2A1O1Ixp33_ASAP7_75t_L g154336__199215 (.A1(n_6122),
    .A2(n_49178),
    .B(n_4426),
    .C(n_48223),
    .Y(n_49179));
 O2A1O1Ixp33_ASAP7_75t_SL g154337__7098 (.A1(n_6122),
    .A2(n_70415),
    .B(n_4428),
    .C(n_48223),
    .Y(n_4434));
 AOI21xp33_ASAP7_75t_SL g154339__198418 (.A1(n_78040),
    .A2(n_70415),
    .B(n_48223),
    .Y(n_48224));
 O2A1O1Ixp33_ASAP7_75t_SL g154340__1705 (.A1(n_2428),
    .A2(n_65298),
    .B(n_14963),
    .C(n_27225),
    .Y(n_4438));
 O2A1O1Ixp33_ASAP7_75t_L g154341__1617 (.A1(n_50292),
    .A2(n_34649),
    .B(n_2424),
    .C(n_27225),
    .Y(n_4441));
 O2A1O1Ixp33_ASAP7_75t_SL g154342__5526 (.A1(n_50292),
    .A2(n_34434),
    .B(n_65298),
    .C(n_27225),
    .Y(n_4445));
 O2A1O1Ixp33_ASAP7_75t_R g154343__4319 (.A1(n_50292),
    .A2(n_4448),
    .B(n_34649),
    .C(n_27225),
    .Y(n_4450));
 O2A1O1Ixp33_ASAP7_75t_SL g154344__6260 (.A1(n_16672),
    .A2(n_2524),
    .B(n_14794),
    .C(n_4485),
    .Y(n_4451));
 O2A1O1Ixp33_ASAP7_75t_SL g154345__5107 (.A1(n_50292),
    .A2(n_41492),
    .B(n_56062),
    .C(n_27225),
    .Y(n_4453));
 AOI21xp33_ASAP7_75t_SL g154346__5122 (.A1(n_2427),
    .A2(n_50291),
    .B(n_27225),
    .Y(n_4384));
 O2A1O1Ixp33_ASAP7_75t_L g154347__8246 (.A1(n_2524),
    .A2(n_46228),
    .B(n_17489),
    .C(n_4485),
    .Y(n_4383));
 O2A1O1Ixp33_ASAP7_75t_SL g154349__6131 (.A1(n_4377),
    .A2(n_2524),
    .B(n_46228),
    .C(n_4485),
    .Y(n_4379));
 AOI21xp33_ASAP7_75t_SL g154350__1881 (.A1(n_2384),
    .A2(n_27368),
    .B(n_27225),
    .Y(n_4375));
 AOI21xp33_ASAP7_75t_SL g154351__5115 (.A1(n_23656),
    .A2(n_2432),
    .B(n_4524),
    .Y(n_4374));
 O2A1O1Ixp33_ASAP7_75t_SL g154352__7482 (.A1(n_176),
    .A2(n_4357),
    .B(n_1957),
    .C(n_4485),
    .Y(n_4373));
 AOI21xp33_ASAP7_75t_SL g154353__4733 (.A1(n_2440),
    .A2(n_2434),
    .B(n_4524),
    .Y(n_4372));
 O2A1O1Ixp33_ASAP7_75t_SL g154354__6161 (.A1(n_13734),
    .A2(n_57041),
    .B(n_1849),
    .C(n_4524),
    .Y(n_4371));
 O2A1O1Ixp33_ASAP7_75t_SL g154355__9315 (.A1(n_13734),
    .A2(n_17617),
    .B(n_1734),
    .C(n_4524),
    .Y(n_4369));
 O2A1O1Ixp33_ASAP7_75t_SL g154356__9945 (.A1(n_176),
    .A2(n_4345),
    .B(n_1959),
    .C(n_4485),
    .Y(n_4366));
 O2A1O1Ixp33_ASAP7_75t_SL g154357__2883 (.A1(n_4362),
    .A2(n_50319),
    .B(n_1846),
    .C(n_4524),
    .Y(n_4364));
 O2A1O1Ixp33_ASAP7_75t_SL g154358__2346 (.A1(n_4362),
    .A2(n_4355),
    .B(n_1852),
    .C(n_4524),
    .Y(n_4363));
 O2A1O1Ixp33_ASAP7_75t_SL g154359__1666 (.A1(n_4353),
    .A2(n_4362),
    .B(n_50319),
    .C(n_4524),
    .Y(n_4361));
 O2A1O1Ixp33_ASAP7_75t_SL g154360__7410 (.A1(n_176),
    .A2(n_66198),
    .B(n_4357),
    .C(n_4485),
    .Y(n_4359));
 O2A1O1Ixp33_ASAP7_75t_SL g154361__6417 (.A1(n_4362),
    .A2(n_4350),
    .B(n_4355),
    .C(n_4524),
    .Y(n_4356));
 O2A1O1Ixp33_ASAP7_75t_SL g154362__224659 (.A1(n_79194),
    .A2(n_41434),
    .B(n_4353),
    .C(n_4524),
    .Y(n_79200));
 O2A1O1Ixp33_ASAP7_75t_SL g154363__224660 (.A1(n_79194),
    .A2(n_4343),
    .B(n_4350),
    .C(n_4524),
    .Y(n_79201));
 O2A1O1Ixp33_ASAP7_75t_L g154364__224657 (.A1(n_79198),
    .A2(n_4341),
    .B(n_41434),
    .C(n_4524),
    .Y(n_79199));
 O2A1O1Ixp33_ASAP7_75t_SL g154365__6260 (.A1(n_4346),
    .A2(n_2524),
    .B(n_4345),
    .C(n_4485),
    .Y(n_4347));
 O2A1O1Ixp33_ASAP7_75t_L g154366__224661 (.A1(n_79194),
    .A2(n_4339),
    .B(n_4343),
    .C(n_4524),
    .Y(n_79202));
 AOI21xp33_ASAP7_75t_L g154367__8428 (.A1(n_4341),
    .A2(n_2345),
    .B(n_4524),
    .Y(n_4342));
 AOI21xp33_ASAP7_75t_SL g154368__5526 (.A1(n_79197),
    .A2(n_4339),
    .B(n_4524),
    .Y(n_4340));
 AOI21xp33_ASAP7_75t_SL g154369__188260 (.A1(n_29074),
    .A2(u11_din_tmp1[7]),
    .B(n_36290),
    .Y(n_36291));
 O2A1O1Ixp33_ASAP7_75t_SL g154370__189852 (.A1(n_725),
    .A2(n_27013),
    .B(n_59640),
    .C(n_38374),
    .Y(n_38379));
 O2A1O1Ixp33_ASAP7_75t_SL g154372__189851 (.A1(n_4332),
    .A2(n_842),
    .B(n_27013),
    .C(n_38374),
    .Y(n_38378));
 O2A1O1Ixp33_ASAP7_75t_SL g154375__189850 (.A1(n_4318),
    .A2(n_4320),
    .B(n_5706),
    .C(n_38374),
    .Y(n_38377));
 O2A1O1Ixp33_ASAP7_75t_SL g154376__189849 (.A1(n_725),
    .A2(n_4316),
    .B(n_4324),
    .C(n_38374),
    .Y(n_38376));
 AOI21xp33_ASAP7_75t_L g154380__189848 (.A1(n_16781),
    .A2(n_15090),
    .B(n_38374),
    .Y(n_38375));
 O2A1O1Ixp33_ASAP7_75t_L g154381__9945 (.A1(n_4548),
    .A2(n_4540),
    .B(n_43305),
    .C(n_64852),
    .Y(n_4541));
 O2A1O1Ixp33_ASAP7_75t_L g154382__6161 (.A1(n_4548),
    .A2(n_23671),
    .B(n_18679),
    .C(n_64852),
    .Y(n_4546));
 O2A1O1Ixp33_ASAP7_75t_SL g154383__4733 (.A1(n_7754),
    .A2(n_4548),
    .B(n_4540),
    .C(n_64852),
    .Y(n_4549));
 O2A1O1Ixp33_ASAP7_75t_L g154384__7482 (.A1(n_46697),
    .A2(n_4548),
    .B(n_23671),
    .C(n_64852),
    .Y(n_4557));
 O2A1O1Ixp33_ASAP7_75t_SL g154386__1881 (.A1(n_14918),
    .A2(n_13825),
    .B(n_1847),
    .C(n_64852),
    .Y(n_4562));
 AOI21xp33_ASAP7_75t_SL g154389__170080 (.A1(n_15080),
    .A2(n_15079),
    .B(n_64852),
    .Y(n_15082));
 O2A1O1Ixp5_ASAP7_75t_SL g154391__1705 (.A1(n_7319),
    .A2(n_14918),
    .B(n_4568),
    .C(n_64852),
    .Y(n_4572));
 AOI21xp33_ASAP7_75t_L g154392__2802 (.A1(n_2393),
    .A2(n_50712),
    .B(n_64852),
    .Y(n_4573));
 AOI21xp33_ASAP7_75t_SL g154393__1617 (.A1(n_2332),
    .A2(n_7319),
    .B(n_64852),
    .Y(n_4574));
 AOI22xp33_ASAP7_75t_R g154395__7482 (.A1(u1_sr[8]),
    .A2(out_le[1]),
    .B1(in_slt1[8]),
    .B2(n_5284),
    .Y(n_5272));
 AOI22xp33_ASAP7_75t_R g154396__4733 (.A1(u1_sr[8]),
    .A2(n_11046),
    .B1(in_slt2[8]),
    .B2(n_5336),
    .Y(n_5271));
 AOI22xp33_ASAP7_75t_R g154399__9945 (.A1(u1_sr[8]),
    .A2(out_le[3]),
    .B1(in_slt3[8]),
    .B2(n_5338),
    .Y(n_5267));
 AOI22xp33_ASAP7_75t_R g154400__9315 (.A1(u1_sr[8]),
    .A2(out_le[4]),
    .B1(in_slt4[8]),
    .B2(n_5341),
    .Y(n_5268));
 AOI22xp33_ASAP7_75t_R g154401__6161 (.A1(u1_sr[8]),
    .A2(out_le[5]),
    .B1(in_slt6[8]),
    .B2(n_5333),
    .Y(n_5269));
 AOI21xp33_ASAP7_75t_SL g154402__182543 (.A1(n_34505),
    .A2(u9_din_tmp1[0]),
    .B(n_29553),
    .Y(n_29554));
 AOI21xp33_ASAP7_75t_SL g154403__182545 (.A1(n_34505),
    .A2(u9_din_tmp1[1]),
    .B(n_29555),
    .Y(n_29556));
 AOI21xp33_ASAP7_75t_SL g154404__182514 (.A1(n_34505),
    .A2(u9_din_tmp1[2]),
    .B(n_29527),
    .Y(n_29528));
 AOI21xp33_ASAP7_75t_SL g154405__182519 (.A1(n_34505),
    .A2(u9_din_tmp1[3]),
    .B(n_29529),
    .Y(n_29530));
 AOI21xp33_ASAP7_75t_SL g154406__186720 (.A1(n_34505),
    .A2(u9_din_tmp1[4]),
    .B(n_34490),
    .Y(n_34491));
 AOI21xp33_ASAP7_75t_SL g154407__182539 (.A1(n_34505),
    .A2(u9_din_tmp1[5]),
    .B(n_29549),
    .Y(n_29550));
 AOI21xp33_ASAP7_75t_SL g154408__182537 (.A1(n_34505),
    .A2(u9_din_tmp1[6]),
    .B(n_29547),
    .Y(n_29548));
 AOI21xp33_ASAP7_75t_SL g154409__182535 (.A1(n_34505),
    .A2(u9_din_tmp1[7]),
    .B(n_29545),
    .Y(n_29546));
 AOI21xp33_ASAP7_75t_SL g154410__182533 (.A1(n_34505),
    .A2(u9_din_tmp1[8]),
    .B(n_29543),
    .Y(n_29544));
 AOI21xp33_ASAP7_75t_SL g154411__186724 (.A1(n_34505),
    .A2(u9_din_tmp1[9]),
    .B(n_34494),
    .Y(n_34495));
 AOI21xp33_ASAP7_75t_SL g154412__186728 (.A1(n_34505),
    .A2(u9_din_tmp1[10]),
    .B(n_34498),
    .Y(n_34499));
 AOI21xp33_ASAP7_75t_SL g154413__186732 (.A1(n_34505),
    .A2(u9_din_tmp1[11]),
    .B(n_34502),
    .Y(n_34503));
 AOI21xp33_ASAP7_75t_SL g154414__182547 (.A1(n_34505),
    .A2(u9_din_tmp1[12]),
    .B(n_29557),
    .Y(n_29558));
 AOI21xp33_ASAP7_75t_SL g154415__186736 (.A1(n_34505),
    .A2(u9_din_tmp1[13]),
    .B(n_34506),
    .Y(n_34507));
 AOI21xp33_ASAP7_75t_SL g154416__182523 (.A1(n_34505),
    .A2(u9_din_tmp1[14]),
    .B(n_29533),
    .Y(n_29534));
 AOI21xp33_ASAP7_75t_SL g154417__182521 (.A1(n_34505),
    .A2(u9_din_tmp1[15]),
    .B(n_29531),
    .Y(n_29532));
 AOI21xp33_ASAP7_75t_SL g154418__182147 (.A1(n_29074),
    .A2(u11_din_tmp1[0]),
    .B(n_29088),
    .Y(n_29089));
 AOI21xp33_ASAP7_75t_SL g154419__186712 (.A1(n_29074),
    .A2(u11_din_tmp1[1]),
    .B(n_34482),
    .Y(n_34483));
 AOI21xp33_ASAP7_75t_SL g154420__182137 (.A1(n_29074),
    .A2(u11_din_tmp1[2]),
    .B(n_29078),
    .Y(n_29079));
 AOI21xp33_ASAP7_75t_SL g154421__186716 (.A1(n_29074),
    .A2(u11_din_tmp1[3]),
    .B(n_34486),
    .Y(n_34487));
 AOI21xp33_ASAP7_75t_SL g154422__182165 (.A1(n_29074),
    .A2(u11_din_tmp1[4]),
    .B(n_29106),
    .Y(n_29107));
 AOI21xp33_ASAP7_75t_SL g154423__182155 (.A1(n_29074),
    .A2(u11_din_tmp1[5]),
    .B(n_29096),
    .Y(n_29097));
 AOI21xp33_ASAP7_75t_SL g154424__182157 (.A1(n_29074),
    .A2(u11_din_tmp1[6]),
    .B(n_29098),
    .Y(n_29099));
 OR2x6_ASAP7_75t_SL g154431__2883 (.A(n_13420),
    .B(n_4276),
    .Y(n_5258));
 OR2x6_ASAP7_75t_SL g154432__168296 (.A(n_4276),
    .B(n_13420),
    .Y(n_12868));
 OR2x6_ASAP7_75t_SL g154433__5122 (.A(n_625),
    .B(n_23286),
    .Y(n_4784));
 OR2x2_ASAP7_75t_SL g154436__168261_dup (.A(n_23285),
    .B(n_23286),
    .Y(n_23289));
 OR2x2_ASAP7_75t_SL g154436__177060 (.A(n_23285),
    .B(n_23286),
    .Y(n_23287));
 INVxp33_ASAP7_75t_R g154437 (.A(u1_sr[9]),
    .Y(n_5273));
 INVx1_ASAP7_75t_SL g154724 (.A(n_7803),
    .Y(n_4496));
 INVxp67_ASAP7_75t_SL g154725 (.A(n_21513),
    .Y(n_4202));
 INVx3_ASAP7_75t_SL g154729 (.A(n_4795),
    .Y(n_4524));
 INVx4_ASAP7_75t_SL g154731 (.A(n_70649),
    .Y(n_4485));
 HB1xp67_ASAP7_75t_R g154739 (.A(n_28696),
    .Y(n_4976));
 INVxp67_ASAP7_75t_R g154745 (.A(n_42249),
    .Y(n_4225));
 INVx1_ASAP7_75t_SL g154757 (.A(n_43090),
    .Y(n_4253));
 INVx1_ASAP7_75t_SL g154759 (.A(n_46183),
    .Y(n_5062));
 INVx1_ASAP7_75t_SL g154762 (.A(n_46182),
    .Y(n_3999));
 INVx1_ASAP7_75t_SL g154770 (.A(n_34541),
    .Y(n_4513));
 INVx1_ASAP7_75t_L g154774 (.A(n_3996),
    .Y(n_4988));
 INVx1_ASAP7_75t_SL g154776 (.A(n_73300),
    .Y(n_3996));
 AOI22xp5_ASAP7_75t_L g154785 (.A1(n_17403),
    .A2(n_3063),
    .B1(u14_u6_full_empty_r),
    .B2(n_20824),
    .Y(n_4070));
 NAND2xp33_ASAP7_75t_R g154792 (.A(n_28884),
    .B(u15_rdd1),
    .Y(n_4146));
 AOI22xp33_ASAP7_75t_R g154838__6417 (.A1(u1_sr[7]),
    .A2(n_10839),
    .B1(in_slt6[7]),
    .B2(n_10813),
    .Y(n_5225));
 AOI22xp33_ASAP7_75t_R g154839__5477 (.A1(u1_sr[7]),
    .A2(n_10709),
    .B1(in_slt4[7]),
    .B2(n_10787),
    .Y(n_5224));
 AOI22xp33_ASAP7_75t_R g154840__2398 (.A1(u1_sr[7]),
    .A2(n_10735),
    .B1(in_slt3[7]),
    .B2(n_10761),
    .Y(n_5223));
 AOI22xp33_ASAP7_75t_R g154841 (.A1(u0_slt9_r[0]),
    .A2(n_9299),
    .B1(out_slt9[1]),
    .B2(n_9348),
    .Y(n_2741));
 A2O1A1Ixp33_ASAP7_75t_SL g154846 (.A1(resume_req),
    .A2(n_2467),
    .B(u2_sync_resume),
    .C(n_607),
    .Y(n_2976));
 A2O1A1Ixp33_ASAP7_75t_SL g154849 (.A1(n_78810),
    .A2(n_18743),
    .B(n_37338),
    .C(n_13968),
    .Y(n_4048));
 AOI22xp33_ASAP7_75t_R g154857__5107 (.A1(u1_sr[7]),
    .A2(out_le[2]),
    .B1(in_slt2[7]),
    .B2(n_5336),
    .Y(n_5222));
 AOI22xp33_ASAP7_75t_R g154858__6260 (.A1(u1_sr[7]),
    .A2(out_le[1]),
    .B1(in_slt1[7]),
    .B2(n_5284),
    .Y(n_5221));
 OR5x1_ASAP7_75t_SL g154859__4319 (.A(n_47768),
    .B(n_17686),
    .C(n_534),
    .D(n_25438),
    .E(u10_wp[3]),
    .Y(n_4224));
 AOI22xp5_ASAP7_75t_SL g154862 (.A1(n_22938),
    .A2(n_2967),
    .B1(u14_u8_full_empty_r),
    .B2(n_18933),
    .Y(n_3993));
 NAND2xp33_ASAP7_75t_SL g154983 (.A(n_684),
    .B(n_12119),
    .Y(n_3991));
 OAI21xp5_ASAP7_75t_SL g154994 (.A1(n_24624),
    .A2(n_24625),
    .B(oc3_cfg[0]),
    .Y(n_4280));
 INVxp67_ASAP7_75t_R g155 (.A(i6_dout[30]),
    .Y(n_65895));
 NOR2xp33_ASAP7_75t_SL g155024 (.A(n_52768),
    .B(n_4116),
    .Y(n_4787));
 NOR2xp33_ASAP7_75t_SL g155025 (.A(n_29310),
    .B(n_4114),
    .Y(n_4792));
 NAND2xp5_ASAP7_75t_SL g155029 (.A(n_13968),
    .B(n_6136),
    .Y(n_4645));
 OAI21xp5_ASAP7_75t_SL g155037 (.A1(n_332),
    .A2(n_425),
    .B(n_70648),
    .Y(n_4261));
 AND2x2_ASAP7_75t_SL g155046 (.A(n_21343),
    .B(n_477),
    .Y(n_4795));
 AND2x2_ASAP7_75t_SL g155050 (.A(n_247),
    .B(n_70324),
    .Y(n_4788));
 INVxp33_ASAP7_75t_R g155073 (.A(u1_sr[8]),
    .Y(n_5263));
 INVxp67_ASAP7_75t_SL g155528 (.A(n_70648),
    .Y(n_4114));
 INVxp67_ASAP7_75t_SL g155529 (.A(n_34234),
    .Y(n_4117));
 INVxp67_ASAP7_75t_SL g155530 (.A(n_70324),
    .Y(n_4116));
 INVxp67_ASAP7_75t_SL g155531 (.A(n_21343),
    .Y(n_4119));
 BUFx3_ASAP7_75t_L g155541 (.A(n_52769),
    .Y(n_5077));
 BUFx2_ASAP7_75t_L g155542 (.A(n_15007),
    .Y(n_5091));
 BUFx2_ASAP7_75t_L g155543 (.A(n_15007),
    .Y(n_5028));
 INVx3_ASAP7_75t_SL g155546_dup188259 (.A(n_29073),
    .Y(n_36289));
 A2O1A1Ixp33_ASAP7_75t_SL g155567 (.A1(n_2454),
    .A2(n_2767),
    .B(n_16009),
    .C(n_552),
    .Y(n_3913));
 AOI31xp33_ASAP7_75t_SL g155573 (.A1(n_21550),
    .A2(n_552),
    .A3(u3_wp[2]),
    .B(n_24374),
    .Y(n_3081));
 AOI31xp33_ASAP7_75t_SL g155575 (.A1(n_33772),
    .A2(n_549),
    .A3(u7_wp[2]),
    .B(n_29365),
    .Y(n_3077));
 NAND4xp25_ASAP7_75t_SL g155577 (.A(n_10622),
    .B(n_7225),
    .C(n_8242),
    .D(n_2281),
    .Y(n_2683));
 AOI22xp33_ASAP7_75t_R g155578__2346 (.A1(u1_sr[6]),
    .A2(out_le[5]),
    .B1(in_slt6[6]),
    .B2(n_5333),
    .Y(n_4537));
 AOI22xp33_ASAP7_75t_R g155579 (.A1(u1_sr[5]),
    .A2(n_10839),
    .B1(in_slt6[5]),
    .B2(n_10813),
    .Y(n_4155));
 AOI22xp5_ASAP7_75t_L g155580 (.A1(n_3908),
    .A2(n_2953),
    .B1(u14_u7_full_empty_r),
    .B2(n_2952),
    .Y(n_3909));
 AOI22xp33_ASAP7_75t_R g155581__1666 (.A1(u1_sr[6]),
    .A2(out_le[4]),
    .B1(in_slt4[6]),
    .B2(n_5341),
    .Y(n_4536));
 AOI22xp33_ASAP7_75t_R g155582__7410 (.A1(u1_sr[6]),
    .A2(out_le[3]),
    .B1(in_slt3[6]),
    .B2(n_5338),
    .Y(n_4535));
 OAI22xp5_ASAP7_75t_SL g155583 (.A1(u14_u7_en_out_l_44),
    .A2(in_valid_s[1]),
    .B1(in_slt0[11]),
    .B2(n_2645),
    .Y(n_2965));
 AOI22xp33_ASAP7_75t_R g155584 (.A1(u1_sr[4]),
    .A2(out_le[5]),
    .B1(in_slt6[4]),
    .B2(n_5333),
    .Y(n_3907));
 AOI22xp33_ASAP7_75t_R g155585 (.A1(u1_sr[3]),
    .A2(n_10839),
    .B1(in_slt6[3]),
    .B2(n_10813),
    .Y(n_2940));
 AOI22xp33_ASAP7_75t_R g155586 (.A1(u1_sr[2]),
    .A2(out_le[5]),
    .B1(in_slt6[2]),
    .B2(n_5333),
    .Y(n_2612));
 AOI22xp33_ASAP7_75t_R g155587 (.A1(u1_sr[1]),
    .A2(out_le[5]),
    .B1(in_slt6[1]),
    .B2(n_5333),
    .Y(n_2574));
 AOI22xp33_ASAP7_75t_R g155588 (.A1(u1_sr[0]),
    .A2(n_10839),
    .B1(in_slt6[0]),
    .B2(n_10813),
    .Y(n_2575));
 AOI22xp33_ASAP7_75t_R g155589__6417 (.A1(u1_sr[6]),
    .A2(n_11046),
    .B1(in_slt2[6]),
    .B2(n_5336),
    .Y(n_4534));
 AOI22xp33_ASAP7_75t_R g155590 (.A1(u1_sr[5]),
    .A2(out_le[2]),
    .B1(in_slt2[5]),
    .B2(n_5336),
    .Y(n_4156));
 AOI22xp33_ASAP7_75t_R g155591 (.A1(u1_sr[4]),
    .A2(n_11046),
    .B1(in_slt2[4]),
    .B2(n_5336),
    .Y(n_3906));
 AOI22xp33_ASAP7_75t_R g155592__5477 (.A1(u1_sr[6]),
    .A2(out_le[1]),
    .B1(in_slt1[6]),
    .B2(n_5284),
    .Y(n_4533));
 AOI22xp33_ASAP7_75t_SL g155600 (.A1(n_64819),
    .A2(n_3815),
    .B1(\u8_mem[3] [1]),
    .B2(n_70622),
    .Y(n_3900));
 AOI22xp5_ASAP7_75t_SL g155631 (.A1(n_11128),
    .A2(n_33203),
    .B1(\u5_mem[3] [0]),
    .B2(n_9476),
    .Y(n_3862));
 AOI22xp5_ASAP7_75t_SL g155632 (.A1(n_11126),
    .A2(n_3815),
    .B1(\u5_mem[3] [1]),
    .B2(n_9476),
    .Y(n_3858));
 AOI22xp5_ASAP7_75t_SL g155658 (.A1(n_11126),
    .A2(n_65910),
    .B1(\u5_mem[3] [27]),
    .B2(n_9476),
    .Y(n_3959));
 AOI22xp33_ASAP7_75t_SL g155732 (.A1(n_66869),
    .A2(n_14570),
    .B1(\u7_mem[3] [5]),
    .B2(n_33772),
    .Y(n_3722));
 AOI22xp33_ASAP7_75t_SL g155733 (.A1(n_32650),
    .A2(n_14570),
    .B1(\u7_mem[3] [6]),
    .B2(n_33772),
    .Y(n_3721));
 AOI22xp33_ASAP7_75t_SL g155734 (.A1(n_65969),
    .A2(n_14570),
    .B1(\u7_mem[3] [7]),
    .B2(n_33772),
    .Y(n_3720));
 AOI22xp33_ASAP7_75t_SL g155735 (.A1(n_65980),
    .A2(n_14570),
    .B1(\u7_mem[3] [8]),
    .B2(n_33772),
    .Y(n_3719));
 AOI22xp33_ASAP7_75t_SL g155736 (.A1(n_79971),
    .A2(n_14570),
    .B1(\u7_mem[3] [9]),
    .B2(n_33772),
    .Y(n_3718));
 AOI22xp33_ASAP7_75t_SL g155737 (.A1(n_65975),
    .A2(n_14570),
    .B1(\u7_mem[3] [10]),
    .B2(n_33772),
    .Y(n_3717));
 AOI22xp33_ASAP7_75t_SL g155738 (.A1(n_66843),
    .A2(n_14570),
    .B1(\u7_mem[3] [11]),
    .B2(n_33772),
    .Y(n_3716));
 AOI22xp33_ASAP7_75t_SL g155740 (.A1(n_35041),
    .A2(n_14570),
    .B1(\u7_mem[3] [13]),
    .B2(n_33772),
    .Y(n_3714));
 AOI22xp33_ASAP7_75t_SL g155741 (.A1(n_66032),
    .A2(n_14570),
    .B1(\u7_mem[3] [14]),
    .B2(n_33772),
    .Y(n_3713));
 AOI22xp33_ASAP7_75t_SL g155742 (.A1(n_28913),
    .A2(n_14570),
    .B1(\u7_mem[3] [15]),
    .B2(n_33772),
    .Y(n_3712));
 AOI22xp33_ASAP7_75t_SL g155744 (.A1(n_65952),
    .A2(n_14570),
    .B1(\u7_mem[3] [17]),
    .B2(n_33772),
    .Y(n_3710));
 AOI22xp33_ASAP7_75t_SL g155745 (.A1(n_14570),
    .A2(n_10194),
    .B1(\u7_mem[3] [18]),
    .B2(n_33772),
    .Y(n_3709));
 AOI22xp33_ASAP7_75t_SL g155759 (.A1(n_47390),
    .A2(n_75733),
    .B1(\u4_mem[3] [0]),
    .B2(n_35908),
    .Y(n_3933));
 AOI22xp5_ASAP7_75t_SL g155760 (.A1(n_30253),
    .A2(n_3815),
    .B1(\u4_mem[3] [1]),
    .B2(n_35908),
    .Y(n_3934));
 AOI22xp5_ASAP7_75t_SL g155761 (.A1(n_66000),
    .A2(n_47390),
    .B1(\u4_mem[3] [2]),
    .B2(n_35908),
    .Y(n_3935));
 AOI22xp5_ASAP7_75t_SL g155762 (.A1(n_66855),
    .A2(n_30253),
    .B1(\u4_mem[3] [3]),
    .B2(n_35908),
    .Y(n_3941));
 AOI22xp33_ASAP7_75t_SL g155767 (.A1(n_65980),
    .A2(n_47390),
    .B1(\u4_mem[3] [8]),
    .B2(n_35908),
    .Y(n_3955));
 AOI22xp5_ASAP7_75t_SL g155768 (.A1(n_30253),
    .A2(n_79972),
    .B1(n_35908),
    .B2(\u4_mem[3] [9]),
    .Y(n_3956));
 AOI22xp33_ASAP7_75t_SL g155770 (.A1(n_66843),
    .A2(n_47390),
    .B1(\u4_mem[3] [11]),
    .B2(n_35908),
    .Y(n_3703));
 AOI22xp5_ASAP7_75t_SL g155771 (.A1(n_65997),
    .A2(n_30253),
    .B1(\u4_mem[3] [12]),
    .B2(n_35908),
    .Y(n_3702));
 AOI22xp5_ASAP7_75t_SL g155772 (.A1(n_47390),
    .A2(n_35041),
    .B1(n_35908),
    .B2(\u4_mem[3] [13]),
    .Y(n_3701));
 AOI22xp33_ASAP7_75t_SL g155773 (.A1(n_66032),
    .A2(n_30253),
    .B1(\u4_mem[3] [14]),
    .B2(n_35908),
    .Y(n_3700));
 AOI22xp33_ASAP7_75t_SL g155774 (.A1(n_28913),
    .A2(n_47390),
    .B1(\u4_mem[3] [15]),
    .B2(n_35908),
    .Y(n_3699));
 AOI22xp33_ASAP7_75t_SL g155775 (.A1(n_47390),
    .A2(n_65949),
    .B1(\u4_mem[3] [16]),
    .B2(n_35908),
    .Y(n_3698));
 AOI22xp33_ASAP7_75t_SL g155776 (.A1(n_65952),
    .A2(n_30253),
    .B1(\u4_mem[3] [17]),
    .B2(n_35908),
    .Y(n_3697));
 AOI22xp5_ASAP7_75t_SL g155827 (.A1(n_33203),
    .A2(n_32163),
    .B1(\u5_mem[1] [0]),
    .B2(n_13500),
    .Y(n_3638));
 AOI22xp33_ASAP7_75t_SL g155828 (.A1(n_3815),
    .A2(n_32164),
    .B1(\u5_mem[1] [1]),
    .B2(n_13508),
    .Y(n_3635));
 AOI22xp5_ASAP7_75t_SL g155838 (.A1(n_16009),
    .A2(n_3815),
    .B1(n_22505),
    .B2(\u3_mem[1] [1]),
    .Y(n_3621));
 INVx1_ASAP7_75t_L g155999 (.A(n_18933),
    .Y(n_2967));
 AOI22xp5_ASAP7_75t_SL g156 (.A1(n_24803),
    .A2(n_50554),
    .B1(\u10_mem[1] [7]),
    .B2(n_32302),
    .Y(n_42801));
 INVx1_ASAP7_75t_SL g156001 (.A(n_20824),
    .Y(n_3063));
 INVxp33_ASAP7_75t_R g156003 (.A(u1_sr[7]),
    .Y(n_4624));
 AOI22xp33_ASAP7_75t_R g156114 (.A1(u1_sr[5]),
    .A2(n_10709),
    .B1(in_slt4[5]),
    .B2(n_10787),
    .Y(n_4177));
 AOI22xp33_ASAP7_75t_R g156115__1881 (.A1(u1_sr[5]),
    .A2(n_10735),
    .B1(in_slt3[5]),
    .B2(n_10761),
    .Y(n_4208));
 AOI22xp33_ASAP7_75t_R g156116__5115 (.A1(u1_sr[5]),
    .A2(out_le[1]),
    .B1(in_slt1[5]),
    .B2(n_5284),
    .Y(n_4207));
 NAND2xp5_ASAP7_75t_SL g156117 (.A(n_13749),
    .B(n_281),
    .Y(n_2957));
 NAND2xp5_ASAP7_75t_SL g156119 (.A(n_64133),
    .B(n_375),
    .Y(n_2956));
 NOR2xp33_ASAP7_75t_SL g156124 (.A(n_2475),
    .B(n_2655),
    .Y(n_2935));
 NOR2xp33_ASAP7_75t_SL g156125 (.A(n_2477),
    .B(n_2657),
    .Y(n_2934));
 NAND3xp33_ASAP7_75t_SL g156126 (.A(n_7219),
    .B(n_10621),
    .C(n_1470),
    .Y(n_2727));
 NOR3xp33_ASAP7_75t_SL g156127 (.A(n_2490),
    .B(n_1887),
    .C(n_2470),
    .Y(n_2933));
 NOR3xp33_ASAP7_75t_SL g156128 (.A(n_2491),
    .B(n_1888),
    .C(n_2496),
    .Y(n_2932));
 NOR3xp33_ASAP7_75t_SL g156129 (.A(n_2492),
    .B(n_1885),
    .C(n_2471),
    .Y(n_2931));
 NAND4xp25_ASAP7_75t_SL g156132 (.A(n_10628),
    .B(n_1483),
    .C(n_7202),
    .D(n_2282),
    .Y(n_2724));
 NAND3xp33_ASAP7_75t_SL g156137 (.A(n_2419),
    .B(n_10624),
    .C(n_7215),
    .Y(n_2721));
 NAND3xp33_ASAP7_75t_SL g156139 (.A(n_10631),
    .B(n_17388),
    .C(n_7212),
    .Y(n_2719));
 NAND3xp33_ASAP7_75t_SL g156143 (.A(n_2413),
    .B(n_10633),
    .C(n_7209),
    .Y(n_2716));
 NAND3xp33_ASAP7_75t_SL g156144 (.A(n_2420),
    .B(n_10617),
    .C(n_7208),
    .Y(n_2715));
 NAND3xp33_ASAP7_75t_SL g156146 (.A(n_10623),
    .B(n_2416),
    .C(n_7206),
    .Y(n_2713));
 NAND3xp33_ASAP7_75t_SL g156147 (.A(n_10636),
    .B(n_47793),
    .C(n_7216),
    .Y(n_2712));
 A2O1A1Ixp33_ASAP7_75t_SL g156157 (.A1(u2_res_cnt[3]),
    .A2(n_31397),
    .B(n_13347),
    .C(u2_sync_resume),
    .Y(n_2817));
 NAND4xp25_ASAP7_75t_SL g156158 (.A(n_7222),
    .B(n_10615),
    .C(n_7167),
    .D(n_6583),
    .Y(n_2977));
 NOR2xp33_ASAP7_75t_SL g156161 (.A(n_29657),
    .B(n_24635),
    .Y(n_2985));
 NOR2xp33_ASAP7_75t_SL g156162 (.A(n_2775),
    .B(n_509),
    .Y(n_2984));
 NOR2xp33_ASAP7_75t_SL g156163 (.A(n_34540),
    .B(n_2773),
    .Y(n_2983));
 OAI31xp33_ASAP7_75t_SL g156167 (.A1(oc1_cfg[4]),
    .A2(o4_status[0]),
    .A3(o4_status[1]),
    .B(n_2951),
    .Y(n_2980));
 OAI21xp5_ASAP7_75t_SL g156172 (.A1(n_21776),
    .A2(u26_ac97_rst_104),
    .B(n_76054),
    .Y(n_2955));
 INVxp33_ASAP7_75t_R g156627 (.A(valid_s1),
    .Y(n_2571));
 INVxp67_ASAP7_75t_SL g156631 (.A(n_2951),
    .Y(n_4040));
 INVx1_ASAP7_75t_SL g156632 (.A(o4_empty),
    .Y(n_2951));
 INVxp67_ASAP7_75t_SL g156633 (.A(n_2990),
    .Y(n_4042));
 INVx1_ASAP7_75t_SL g156634 (.A(o7_empty),
    .Y(n_2990));
 INVxp67_ASAP7_75t_SL g156635 (.A(n_2950),
    .Y(n_3937));
 INVx1_ASAP7_75t_SL g156636 (.A(o6_empty),
    .Y(n_2950));
 INVx1_ASAP7_75t_SL g156640 (.A(o9_empty),
    .Y(n_2964));
 INVx1_ASAP7_75t_L g156642 (.A(n_2952),
    .Y(n_2953));
 HB1xp67_ASAP7_75t_SL g156643 (.A(in_valid_s[1]),
    .Y(n_2952));
 INVxp33_ASAP7_75t_R g156644 (.A(u1_sr[6]),
    .Y(n_4230));
 INVxp33_ASAP7_75t_R g156645 (.A(out_le[0]),
    .Y(n_5296));
 INVxp33_ASAP7_75t_R g156646 (.A(out_le[2]),
    .Y(n_5336));
 INVxp33_ASAP7_75t_R g156648 (.A(out_le[5]),
    .Y(n_5333));
 INVx5_ASAP7_75t_SL g156665_dup166718 (.A(n_11125),
    .Y(n_11128));
 AND2x2_ASAP7_75t_R g156687 (.A(u15_crac_we_r),
    .B(crac_out[31]),
    .Y(n_2947));
 NAND2xp33_ASAP7_75t_R g156688 (.A(out_slt9[0]),
    .B(n_9345),
    .Y(n_2277));
 O2A1O1Ixp33_ASAP7_75t_SL g156701 (.A1(i3_re),
    .A2(n_13035),
    .B(n_2306),
    .C(n_8186),
    .Y(n_2708));
 O2A1O1Ixp33_ASAP7_75t_SL g156703 (.A1(i6_re),
    .A2(n_13027),
    .B(n_2304),
    .C(n_19),
    .Y(n_2706));
 OAI211xp5_ASAP7_75t_SL g156706 (.A1(n_63),
    .A2(n_10613),
    .B(n_1475),
    .C(n_7168),
    .Y(n_2657));
 OAI211xp5_ASAP7_75t_SL g156707 (.A1(n_218),
    .A2(n_10613),
    .B(n_1488),
    .C(n_7172),
    .Y(n_2655));
 NAND3xp33_ASAP7_75t_L g156710 (.A(n_2369),
    .B(n_7218),
    .C(n_1329),
    .Y(n_2653));
 AOI221xp5_ASAP7_75t_R g156711 (.A1(n_2020),
    .A2(u2_cnt[7]),
    .B1(n_2021),
    .B2(n_2119),
    .C(n_2465),
    .Y(n_2567));
 NAND2xp5_ASAP7_75t_SL g156712 (.A(n_35476),
    .B(u2_sync_resume),
    .Y(n_2652));
 AOI21xp33_ASAP7_75t_R g156713 (.A1(i4_re),
    .A2(i4_empty),
    .B(ic1_int_set[1]),
    .Y(n_2566));
 AOI21xp33_ASAP7_75t_R g156714 (.A1(i6_re),
    .A2(i6_empty),
    .B(ic2_int_set[1]),
    .Y(n_2565));
 AOI21xp33_ASAP7_75t_R g156715 (.A1(i3_re),
    .A2(i3_empty),
    .B(ic0_int_set[1]),
    .Y(n_2564));
 AOI211xp5_ASAP7_75t_R g156718 (.A1(n_2330),
    .A2(u2_cnt[6]),
    .B(n_2217),
    .C(n_2467),
    .Y(n_2560));
 AOI22xp33_ASAP7_75t_R g156719 (.A1(u1_sr[0]),
    .A2(n_10735),
    .B1(in_slt3[0]),
    .B2(n_10761),
    .Y(n_2275));
 AOI22xp33_ASAP7_75t_R g156720 (.A1(u1_sr[1]),
    .A2(out_le[3]),
    .B1(in_slt3[1]),
    .B2(n_5338),
    .Y(n_2274));
 AOI22xp33_ASAP7_75t_R g156721 (.A1(u1_sr[2]),
    .A2(out_le[3]),
    .B1(in_slt3[2]),
    .B2(n_5338),
    .Y(n_2651));
 AOI22xp33_ASAP7_75t_R g156722 (.A1(u1_sr[3]),
    .A2(n_10735),
    .B1(in_slt3[3]),
    .B2(n_10761),
    .Y(n_2948));
 AOI22xp33_ASAP7_75t_R g156723 (.A1(u1_sr[4]),
    .A2(out_le[3]),
    .B1(in_slt3[4]),
    .B2(n_5338),
    .Y(n_3948));
 AOI22xp33_ASAP7_75t_R g156724 (.A1(u1_sr[4]),
    .A2(out_le[4]),
    .B1(in_slt4[4]),
    .B2(n_5341),
    .Y(n_3947));
 AOI22xp5_ASAP7_75t_SL g156728 (.A1(n_43468),
    .A2(n_1649),
    .B1(n_2237),
    .B2(n_1861),
    .Y(n_2702));
 AND2x4_ASAP7_75t_SL g156760_169534 (.A(n_69795),
    .B(n_14385),
    .Y(n_14386));
 OR2x2_ASAP7_75t_SL g156762_dup165229_dup187967 (.A(n_35904),
    .B(n_26050),
    .Y(n_35909));
 OR2x6_ASAP7_75t_SL g156762_dup166760_dup187969 (.A(n_26050),
    .B(n_35904),
    .Y(n_35911));
 OR2x6_ASAP7_75t_SL g156762_dup187968 (.A(n_26050),
    .B(n_35904),
    .Y(n_35910));
 AND3x4_ASAP7_75t_SL g156764 (.A(n_232),
    .B(n_11124),
    .C(o6_we),
    .Y(n_2836));
 OR2x6_ASAP7_75t_SL g156770_dup214508 (.A(n_69796),
    .B(n_29352),
    .Y(n_67568));
 OR2x2_ASAP7_75t_L g156772_dup165220_dup (.A(n_24367),
    .B(n_11124),
    .Y(n_11135));
 OR2x6_ASAP7_75t_SL g156772_dup166716 (.A(n_24367),
    .B(n_11124),
    .Y(n_11125));
 OR2x2_ASAP7_75t_SL g156773_dup165222_dup (.A(n_70621),
    .B(n_64192),
    .Y(n_11204));
 AOI22xp33_ASAP7_75t_SL g156870 (.A1(n_2743),
    .A2(u8_wp[0]),
    .B1(n_78931),
    .B2(o9_we),
    .Y(n_2775));
 AOI22xp33_ASAP7_75t_SL g156872 (.A1(n_40418),
    .A2(n_2748),
    .B1(n_24373),
    .B2(o3_we),
    .Y(n_2773));
 INVxp33_ASAP7_75t_R g156876 (.A(in_valid_s1[1]),
    .Y(n_2557));
 INVxp33_ASAP7_75t_R g156877 (.A(in_valid[0]),
    .Y(n_2442));
 INVxp33_ASAP7_75t_R g156878 (.A(valid),
    .Y(n_2190));
 INVxp33_ASAP7_75t_R g156879 (.A(in_valid[2]),
    .Y(n_2271));
 INVxp33_ASAP7_75t_R g156882 (.A(n_12142),
    .Y(n_2767));
 INVxp33_ASAP7_75t_R g156892 (.A(u1_sr[5]),
    .Y(n_4003));
 INVxp33_ASAP7_75t_R g156893 (.A(out_le[1]),
    .Y(n_5284));
 INVx3_ASAP7_75t_SL g156894 (.A(n_47786),
    .Y(n_3415));
 INVx3_ASAP7_75t_SL g156895 (.A(n_47786),
    .Y(n_3425));
 BUFx12f_ASAP7_75t_SL g156896 (.A(n_47786),
    .Y(n_3420));
 INVx3_ASAP7_75t_SL g156902 (.A(n_43534),
    .Y(n_3386));
 INVx3_ASAP7_75t_SL g156903 (.A(n_43534),
    .Y(n_3365));
 INVx3_ASAP7_75t_SL g156906 (.A(n_19383),
    .Y(n_3453));
 INVx3_ASAP7_75t_SL g156907 (.A(n_19383),
    .Y(n_3460));
 BUFx6f_ASAP7_75t_SL g156908 (.A(n_19383),
    .Y(n_3454));
 BUFx6f_ASAP7_75t_SL g156909 (.A(n_19383),
    .Y(n_3461));
 INVxp33_ASAP7_75t_R g156919 (.A(ld),
    .Y(n_5529));
 INVxp33_ASAP7_75t_R g156920 (.A(n_9394),
    .Y(n_5532));
 INVxp33_ASAP7_75t_R g156921 (.A(n_9395),
    .Y(n_5522));
 OAI221xp5_ASAP7_75t_SL g156929 (.A1(n_1739),
    .A2(n_23655),
    .B1(n_57084),
    .B2(n_4339),
    .C(n_2434),
    .Y(n_2435));
 OAI221xp5_ASAP7_75t_SL g156931 (.A1(n_40904),
    .A2(n_23655),
    .B1(n_4341),
    .B2(n_57084),
    .C(n_2432),
    .Y(n_2433));
 NOR2xp33_ASAP7_75t_SL g156936 (.A(n_1503),
    .B(n_8306),
    .Y(n_2647));
 NOR2xp33_ASAP7_75t_SL g156937 (.A(n_2645),
    .B(n_8306),
    .Y(n_2646));
 NOR2xp33_ASAP7_75t_SL g156938 (.A(n_1376),
    .B(n_8306),
    .Y(n_2644));
 OAI221xp5_ASAP7_75t_SL g156940 (.A1(n_65298),
    .A2(n_2428),
    .B1(n_64715),
    .B2(n_2427),
    .C(n_19687),
    .Y(n_2429));
 NOR2xp33_ASAP7_75t_SL g156941 (.A(n_1496),
    .B(n_8306),
    .Y(n_2643));
 NOR2xp33_ASAP7_75t_SL g156942 (.A(n_1494),
    .B(n_8306),
    .Y(n_2642));
 NOR2xp33_ASAP7_75t_SL g156943 (.A(n_2640),
    .B(n_8306),
    .Y(n_2641));
 NOR2xp33_ASAP7_75t_SL g156944 (.A(n_25293),
    .B(n_8306),
    .Y(n_2639));
 NOR2xp33_ASAP7_75t_SL g156945 (.A(n_1379),
    .B(n_8306),
    .Y(n_2660));
 NOR2xp33_ASAP7_75t_SL g156957 (.A(n_1501),
    .B(n_8306),
    .Y(n_2624));
 NOR2xp33_ASAP7_75t_SL g156958 (.A(n_88),
    .B(n_8306),
    .Y(n_2623));
 NOR2xp33_ASAP7_75t_SL g156962 (.A(n_143),
    .B(n_8306),
    .Y(n_2620));
 NOR2xp33_ASAP7_75t_SL g156963 (.A(n_12),
    .B(n_8306),
    .Y(n_2619));
 NOR2xp33_ASAP7_75t_SL g156968 (.A(n_19),
    .B(n_8306),
    .Y(n_2650));
 O2A1O1Ixp33_ASAP7_75t_R g156969 (.A1(u4_wp[2]),
    .A2(n_65325),
    .B(n_368),
    .C(n_24632),
    .Y(n_2696));
 O2A1O1Ixp33_ASAP7_75t_R g156970 (.A1(u5_wp[2]),
    .A2(n_455),
    .B(n_456),
    .C(n_2746),
    .Y(n_2695));
 O2A1O1Ixp33_ASAP7_75t_R g156971 (.A1(u6_wp[2]),
    .A2(n_2693),
    .B(n_369),
    .C(n_50109),
    .Y(n_2694));
 O2A1O1Ixp33_ASAP7_75t_R g156972 (.A1(u7_wp[2]),
    .A2(n_2691),
    .B(n_464),
    .C(n_2752),
    .Y(n_2692));
 O2A1O1Ixp33_ASAP7_75t_R g156974 (.A1(u3_wp[2]),
    .A2(n_2687),
    .B(n_469),
    .C(n_2748),
    .Y(n_2688));
 NOR2xp33_ASAP7_75t_SL g156975 (.A(n_431),
    .B(n_8306),
    .Y(n_2595));
 NOR2xp33_ASAP7_75t_SL g156976 (.A(n_330),
    .B(n_8306),
    .Y(n_2573));
 NOR2xp33_ASAP7_75t_SL g156977 (.A(n_423),
    .B(n_8306),
    .Y(n_2611));
 NOR2xp33_ASAP7_75t_SL g156978 (.A(n_50546),
    .B(n_8306),
    .Y(n_2610));
 NOR2xp33_ASAP7_75t_SL g156979 (.A(n_435),
    .B(n_8306),
    .Y(n_2609));
 NOR2xp33_ASAP7_75t_SL g156980 (.A(n_50452),
    .B(n_8306),
    .Y(n_2608));
 AOI221xp5_ASAP7_75t_SL g156981 (.A1(n_7084),
    .A2(u13_intm_r[2]),
    .B1(i4_dout[2]),
    .B2(n_8173),
    .C(n_10878),
    .Y(n_2420));
 AOI221xp5_ASAP7_75t_SL g156982 (.A1(n_7082),
    .A2(u13_intm_r[12]),
    .B1(i4_dout[12]),
    .B2(n_8174),
    .C(n_10871),
    .Y(n_2419));
 AOI221xp5_ASAP7_75t_SL g156983 (.A1(n_7082),
    .A2(u13_intm_r[0]),
    .B1(i4_dout[0]),
    .B2(n_8174),
    .C(n_10881),
    .Y(n_2418));
 AOI221xp5_ASAP7_75t_SL g156984 (.A1(n_7083),
    .A2(u13_intm_r[7]),
    .B1(i4_dout[7]),
    .B2(n_8174),
    .C(n_10887),
    .Y(n_2416));
 AOI221xp5_ASAP7_75t_SL g156986 (.A1(n_7082),
    .A2(n_307),
    .B1(i4_dout[4]),
    .B2(n_8174),
    .C(n_10882),
    .Y(n_2413));
 OAI31xp33_ASAP7_75t_SL g156993 (.A1(ic0_cfg[4]),
    .A2(i3_status[0]),
    .A3(i3_status[1]),
    .B(n_2226),
    .Y(n_2546));
 OAI31xp33_ASAP7_75t_SL g156995 (.A1(ic2_cfg[4]),
    .A2(i6_status[0]),
    .A3(i6_status[1]),
    .B(n_2227),
    .Y(n_2544));
 AOI22xp5_ASAP7_75t_SL g157 (.A1(\u8_mem[3] [10]),
    .A2(n_78273),
    .B1(n_79178),
    .B2(\u8_mem[2] [10]),
    .Y(n_71350));
 NAND3xp33_ASAP7_75t_SL g157003 (.A(n_2685),
    .B(n_1797),
    .C(n_2298),
    .Y(n_2686));
 OAI211xp5_ASAP7_75t_SL g157006 (.A1(n_13734),
    .A2(n_4343),
    .B(n_1436),
    .C(n_2263),
    .Y(n_2603));
 OAI211xp5_ASAP7_75t_SL g157010 (.A1(n_4318),
    .A2(n_4316),
    .B(n_1456),
    .C(n_52979),
    .Y(n_2598));
 NAND4xp25_ASAP7_75t_SL g157015 (.A(n_28893),
    .B(n_8128),
    .C(n_1749),
    .D(n_77397),
    .Y(n_2539));
 OAI221xp5_ASAP7_75t_SL g157028 (.A1(n_34649),
    .A2(n_2428),
    .B1(n_2384),
    .B2(n_64715),
    .C(n_56871),
    .Y(n_2385));
 O2A1O1Ixp33_ASAP7_75t_SL g157063 (.A1(oc1_cfg[4]),
    .A2(o4_status[0]),
    .B(o4_status[1]),
    .C(oc1_cfg[5]),
    .Y(n_2522));
 O2A1O1Ixp33_ASAP7_75t_SL g157065 (.A1(oc4_cfg[4]),
    .A2(o8_status[0]),
    .B(o8_status[1]),
    .C(oc4_cfg[5]),
    .Y(n_2520));
 O2A1O1Ixp33_ASAP7_75t_SL g157067 (.A1(ic0_cfg[4]),
    .A2(i3_status[0]),
    .B(i3_status[1]),
    .C(ic0_cfg[5]),
    .Y(n_2373));
 O2A1O1Ixp33_ASAP7_75t_L g157069 (.A1(ic2_cfg[4]),
    .A2(i6_status[0]),
    .B(i6_status[1]),
    .C(ic2_cfg[5]),
    .Y(n_2371));
 NAND5xp2_ASAP7_75t_R g157070 (.A(n_1535),
    .B(n_1903),
    .C(n_1914),
    .D(u2_cnt[3]),
    .E(u2_cnt[7]),
    .Y(n_1915));
 NAND2xp5_ASAP7_75t_SL g157071 (.A(n_28811),
    .B(u2_sync_resume),
    .Y(n_2519));
 AOI22xp5_ASAP7_75t_R g157073 (.A1(n_14933),
    .A2(i6_dout[31]),
    .B1(n_8173),
    .B2(i4_dout[31]),
    .Y(n_2369));
 OAI22xp5_ASAP7_75t_SL g157074 (.A1(n_65895),
    .A2(n_7170),
    .B1(n_6956),
    .B2(n_2517),
    .Y(n_2518));
 OAI22xp5_ASAP7_75t_SL g157075 (.A1(n_2203),
    .A2(n_7170),
    .B1(n_212),
    .B2(n_6956),
    .Y(n_2516));
 OAI211xp5_ASAP7_75t_SL g157078 (.A1(n_34649),
    .A2(n_15100),
    .B(n_7523),
    .C(n_2511),
    .Y(n_2513));
 OAI211xp5_ASAP7_75t_SL g157080 (.A1(n_5674),
    .A2(n_46227),
    .B(n_20760),
    .C(n_2230),
    .Y(n_2594));
 NAND4xp25_ASAP7_75t_SL g157082 (.A(n_1426),
    .B(n_2362),
    .C(n_1411),
    .D(n_36769),
    .Y(n_2363));
 OAI211xp5_ASAP7_75t_SL g157084 (.A1(n_65298),
    .A2(n_15100),
    .B(n_2508),
    .C(n_65054),
    .Y(n_2509));
 NAND4xp25_ASAP7_75t_SL g157094 (.A(n_28246),
    .B(n_1400),
    .C(n_1420),
    .D(n_78040),
    .Y(n_2350));
 OAI211xp5_ASAP7_75t_SL g157098 (.A1(n_15100),
    .A2(n_34434),
    .B(n_2143),
    .C(n_2540),
    .Y(n_2541));
 NAND4xp25_ASAP7_75t_SL g157103 (.A(n_1440),
    .B(n_2446),
    .C(n_1390),
    .D(n_2059),
    .Y(n_2447));
 NAND4xp25_ASAP7_75t_SL g157107 (.A(n_2053),
    .B(n_2014),
    .C(n_1434),
    .D(n_1387),
    .Y(n_2348));
 NOR5xp2_ASAP7_75t_SL g157115 (.A(n_509),
    .B(n_14763),
    .C(n_2743),
    .D(n_78931),
    .E(u8_wp[2]),
    .Y(n_2744));
 OR3x1_ASAP7_75t_R g157116 (.A(n_1894),
    .B(u2_cnt[5]),
    .C(u2_cnt[3]),
    .Y(n_2129));
 OR5x1_ASAP7_75t_R g157118 (.A(n_1044),
    .B(n_517),
    .C(n_181),
    .D(n_35645),
    .E(n_37457),
    .Y(n_1913));
 NAND2xp5_ASAP7_75t_SL g157127 (.A(n_19008),
    .B(n_2265),
    .Y(n_2492));
 NAND2xp5_ASAP7_75t_SL g157128 (.A(n_1484),
    .B(n_2266),
    .Y(n_2491));
 NAND2xp5_ASAP7_75t_SL g157129 (.A(n_1490),
    .B(n_2268),
    .Y(n_2490));
 NAND4xp25_ASAP7_75t_SL g157137 (.A(n_35466),
    .B(n_34102),
    .C(n_1812),
    .D(n_1755),
    .Y(n_2337));
 OAI211xp5_ASAP7_75t_SL g157139 (.A1(n_8113),
    .A2(n_4540),
    .B(n_2232),
    .C(n_7806),
    .Y(n_2584));
 OAI211xp5_ASAP7_75t_SL g157144 (.A1(n_15079),
    .A2(n_8113),
    .B(n_2234),
    .C(n_2578),
    .Y(n_2579));
 O2A1O1Ixp33_ASAP7_75t_R g157146 (.A1(n_1841),
    .A2(u2_cnt[5]),
    .B(n_2330),
    .C(n_2465),
    .Y(n_2331));
 NAND3xp33_ASAP7_75t_R g157153 (.A(n_1895),
    .B(u2_cnt[5]),
    .C(u2_cnt[3]),
    .Y(n_2223));
 AOI22xp33_ASAP7_75t_R g157156 (.A1(u1_sr[0]),
    .A2(n_10709),
    .B1(in_slt4[0]),
    .B2(n_10787),
    .Y(n_2479));
 AOI22xp33_ASAP7_75t_R g157157 (.A1(u1_sr[2]),
    .A2(out_le[4]),
    .B1(in_slt4[2]),
    .B2(n_5341),
    .Y(n_2576));
 AOI22xp33_ASAP7_75t_R g157158 (.A1(u1_sr[3]),
    .A2(n_10709),
    .B1(in_slt4[3]),
    .B2(n_10787),
    .Y(n_2941));
 AOI22xp33_ASAP7_75t_R g157159 (.A1(u1_sr[1]),
    .A2(out_le[4]),
    .B1(in_slt4[1]),
    .B2(n_5341),
    .Y(n_2478));
 OAI21xp33_ASAP7_75t_SL g157163 (.A1(n_8340),
    .A2(n_2206),
    .B(n_2256),
    .Y(n_2477));
 OAI21xp33_ASAP7_75t_SL g157164 (.A1(n_2205),
    .A2(n_8340),
    .B(n_2261),
    .Y(n_2475));
 OAI21xp5_ASAP7_75t_SL g157166 (.A1(n_2179),
    .A2(n_8340),
    .B(n_2278),
    .Y(n_2473));
 OAI21xp5_ASAP7_75t_SL g157183 (.A1(n_2208),
    .A2(n_8340),
    .B(n_7176),
    .Y(n_2471));
 OAI21xp5_ASAP7_75t_SL g157184 (.A1(n_2207),
    .A2(n_8340),
    .B(n_7173),
    .Y(n_2496));
 OAI21xp5_ASAP7_75t_SL g157185 (.A1(n_2180),
    .A2(n_8340),
    .B(n_7171),
    .Y(n_2470));
 AND3x4_ASAP7_75t_SL g157188 (.A(n_2664),
    .B(n_2663),
    .C(o8_we),
    .Y(n_3188));
 AND3x4_ASAP7_75t_SL g157189 (.A(n_2664),
    .B(n_2663),
    .C(o8_we),
    .Y(n_2737));
 AND3x4_ASAP7_75t_SL g157193 (.A(n_24805),
    .B(n_24804),
    .C(o3_we),
    .Y(n_2735));
 AND3x4_ASAP7_75t_SL g157194 (.A(n_169),
    .B(n_2669),
    .C(o6_we),
    .Y(n_3285));
 AND3x4_ASAP7_75t_SL g157195 (.A(n_231),
    .B(o6_we),
    .C(n_2669),
    .Y(n_2734));
 AND3x4_ASAP7_75t_SL g157196 (.A(n_78931),
    .B(o9_we),
    .C(n_64814),
    .Y(n_3320));
 AND3x4_ASAP7_75t_SL g157197 (.A(n_78931),
    .B(o9_we),
    .C(n_64814),
    .Y(n_2733));
 INVxp33_ASAP7_75t_R g157198 (.A(in_valid[1]),
    .Y(n_2222));
 INVxp33_ASAP7_75t_R g157199 (.A(u1_sr[4]),
    .Y(n_2974));
 INVx1_ASAP7_75t_L g157202 (.A(o8_we),
    .Y(n_2752));
 INVx1_ASAP7_75t_L g157203 (.A(o6_we),
    .Y(n_2746));
 INVx1_ASAP7_75t_L g157204 (.A(o9_we),
    .Y(n_2743));
 INVxp67_ASAP7_75t_SL g157205 (.A(o3_we),
    .Y(n_2748));
 INVxp33_ASAP7_75t_R g157207 (.A(out_le[3]),
    .Y(n_5338));
 NAND2xp5_ASAP7_75t_L g157212 (.A(i4_dout[22]),
    .B(n_8173),
    .Y(n_2268));
 NAND2xp5_ASAP7_75t_L g157214 (.A(i4_dout[21]),
    .B(n_8173),
    .Y(n_2266));
 NAND2xp5_ASAP7_75t_SL g157215 (.A(n_8173),
    .B(i4_dout[20]),
    .Y(n_2265));
 NAND2xp33_ASAP7_75t_R g157220 (.A(i4_dout[1]),
    .B(n_8173),
    .Y(n_2281));
 NAND2xp33_ASAP7_75t_R g157221 (.A(i4_dout[17]),
    .B(n_8173),
    .Y(n_2282));
 NAND2xp5_ASAP7_75t_L g157223 (.A(n_8173),
    .B(i4_dout[27]),
    .Y(n_2273));
 NAND2xp5_ASAP7_75t_SL g157224 (.A(n_8174),
    .B(i4_dout[28]),
    .Y(n_2278));
 NOR2xp33_ASAP7_75t_R g157226 (.A(u2_bit_clk_e),
    .B(n_258),
    .Y(n_2237));
 NAND2xp5_ASAP7_75t_SL g157270 (.A(n_8174),
    .B(i4_dout[26]),
    .Y(n_2261));
 NAND2xp5_ASAP7_75t_L g157275 (.A(n_8174),
    .B(i4_dout[25]),
    .Y(n_2256));
 XOR2xp5_ASAP7_75t_SL g157279 (.A(n_16),
    .B(n_43604),
    .Y(n_2124));
 NAND2xp33_ASAP7_75t_SL g157280 (.A(n_13035),
    .B(i3_re),
    .Y(n_2306));
 NAND2xp33_ASAP7_75t_SL g157281 (.A(n_13027),
    .B(i6_re),
    .Y(n_2304));
 AOI222xp33_ASAP7_75t_SL g157285 (.A1(n_36528),
    .A2(n_67490),
    .B1(\u8_mem[0] [29]),
    .B2(n_27133),
    .C1(\u8_mem[1] [29]),
    .C2(n_27134),
    .Y(n_2254));
 AO21x1_ASAP7_75t_R g157286 (.A1(n_1903),
    .A2(n_1083),
    .B(n_2119),
    .Y(n_1904));
 NOR2xp33_ASAP7_75t_R g157287 (.A(u2_cnt[6]),
    .B(n_2330),
    .Y(n_2217));
 AOI311xp33_ASAP7_75t_R g157289 (.A1(u2_cnt[4]),
    .A2(u2_cnt[5]),
    .A3(n_1082),
    .B(u2_cnt[7]),
    .C(u2_cnt[6]),
    .Y(n_1651));
 OAI21xp5_ASAP7_75t_SL g157290 (.A1(n_42621),
    .A2(n_18885),
    .B(n_31561),
    .Y(n_2216));
 NAND5xp2_ASAP7_75t_R g157291 (.A(n_1336),
    .B(n_633),
    .C(n_1903),
    .D(n_1192),
    .E(n_2288),
    .Y(n_1337));
 NOR3xp33_ASAP7_75t_R g157293 (.A(n_13758),
    .B(n_8186),
    .C(i3_re),
    .Y(n_2452));
 NOR3xp33_ASAP7_75t_R g157294 (.A(n_19),
    .B(n_13764),
    .C(i6_re),
    .Y(n_2453));
 AND3x1_ASAP7_75t_R g157295 (.A(n_2119),
    .B(n_1330),
    .C(n_588),
    .Y(n_2120));
 NAND2xp5_ASAP7_75t_SL g157296 (.A(n_59764),
    .B(u2_sync_resume),
    .Y(n_2251));
 NAND5xp2_ASAP7_75t_R g157297 (.A(n_1336),
    .B(n_1193),
    .C(u2_cnt[5]),
    .D(n_1192),
    .E(u2_cnt[2]),
    .Y(n_1194));
 OAI21xp33_ASAP7_75t_SL g157298 (.A1(n_1343),
    .A2(n_321),
    .B(n_2286),
    .Y(n_2302));
 AND3x1_ASAP7_75t_SL g157299 (.A(u13_csr[1]),
    .B(n_7196),
    .C(n_8336),
    .Y(n_2118));
 AOI222xp33_ASAP7_75t_SL g157306 (.A1(n_47551),
    .A2(n_66199),
    .B1(n_24512),
    .B2(\u3_mem[0] [28]),
    .C1(n_24513),
    .C2(\u3_mem[1] [28]),
    .Y(n_2298));
 AOI221xp5_ASAP7_75t_SL g157307 (.A1(n_24512),
    .A2(\u3_mem[0] [29]),
    .B1(n_47551),
    .B2(n_2168),
    .C(n_1296),
    .Y(n_2247));
 AOI221x1_ASAP7_75t_SL g157316 (.A1(n_24512),
    .A2(\u3_mem[0] [24]),
    .B1(n_47551),
    .B2(n_40287),
    .C(n_1286),
    .Y(n_2238));
 AOI222xp33_ASAP7_75t_SL g157317 (.A1(n_36528),
    .A2(n_16458),
    .B1(\u8_mem[0] [27]),
    .B2(n_27133),
    .C1(\u8_mem[1] [27]),
    .C2(n_27134),
    .Y(n_2263));
 AOI222xp33_ASAP7_75t_SL g157318 (.A1(n_36528),
    .A2(n_70887),
    .B1(\u8_mem[0] [28]),
    .B2(n_27133),
    .C1(\u8_mem[1] [28]),
    .C2(n_27134),
    .Y(n_2236));
 AND2x4_ASAP7_75t_SL g157327_dup (.A(n_7084),
    .B(rf_we),
    .Y(n_6748));
 INVxp67_ASAP7_75t_R g157331 (.A(i3_dout[20]),
    .Y(n_2208));
 INVxp67_ASAP7_75t_R g157332 (.A(i3_dout[21]),
    .Y(n_2207));
 INVxp67_ASAP7_75t_R g157333 (.A(i3_dout[22]),
    .Y(n_2180));
 INVxp33_ASAP7_75t_R g157334 (.A(i3_dout[25]),
    .Y(n_2206));
 INVxp33_ASAP7_75t_R g157335 (.A(i3_dout[26]),
    .Y(n_2205));
 INVxp67_ASAP7_75t_R g157337 (.A(i3_dout[28]),
    .Y(n_2179));
 INVx1_ASAP7_75t_L g157338 (.A(i4_dout[23]),
    .Y(n_2235));
 INVxp67_ASAP7_75t_R g157339 (.A(i6_dout[29]),
    .Y(n_2203));
 INVxp33_ASAP7_75t_R g157341 (.A(n_2020),
    .Y(n_2021));
 INVx1_ASAP7_75t_SL g157343 (.A(i3_full),
    .Y(n_2226));
 INVx1_ASAP7_75t_L g157345 (.A(u2_bit_clk_e),
    .Y(n_2286));
 INVx1_ASAP7_75t_SL g157347 (.A(i6_full),
    .Y(n_2227));
 INVxp33_ASAP7_75t_R g157348 (.A(n_2228),
    .Y(n_3908));
 INVx1_ASAP7_75t_L g157349 (.A(i4_full),
    .Y(n_2228));
 INVxp33_ASAP7_75t_R g157350 (.A(u1_sr[3]),
    .Y(n_2684));
 INVxp33_ASAP7_75t_R g157353 (.A(out_le[4]),
    .Y(n_5341));
 NAND2xp5_ASAP7_75t_SL g157433 (.A(n_37200),
    .B(n_21015),
    .Y(n_2195));
 NAND2xp5_ASAP7_75t_SL g157454 (.A(n_37200),
    .B(n_36969),
    .Y(n_2193));
 NAND2xp5_ASAP7_75t_SL g157462 (.A(n_47551),
    .B(n_50344),
    .Y(n_2191));
 NAND2xp5_ASAP7_75t_L g157463 (.A(n_47551),
    .B(n_48729),
    .Y(n_2224));
 NOR2xp33_ASAP7_75t_R g157464 (.A(n_2465),
    .B(n_2288),
    .Y(n_2289));
 NOR3xp33_ASAP7_75t_L g157465 (.A(n_1648),
    .B(n_1647),
    .C(n_362),
    .Y(n_1649));
 NAND2xp33_ASAP7_75t_R g157469 (.A(n_1645),
    .B(n_1841),
    .Y(n_2020));
 NAND2xp5_ASAP7_75t_SL g157477 (.A(n_7570),
    .B(n_573),
    .Y(n_2685));
 NAND2xp5_ASAP7_75t_SL g157479 (.A(n_2188),
    .B(n_53003),
    .Y(n_2486));
 NAND2xp5_ASAP7_75t_SL g157480 (.A(n_644),
    .B(n_41637),
    .Y(n_2185));
 NAND2xp5_ASAP7_75t_L g157483 (.A(n_644),
    .B(n_31445),
    .Y(n_2183));
 AO21x1_ASAP7_75t_SL g157487 (.A1(n_1338),
    .A2(n_1346),
    .B(n_4548),
    .Y(n_2332));
 NAND2xp5_ASAP7_75t_SL g157493 (.A(n_34203),
    .B(n_78041),
    .Y(n_2362));
 NAND2xp5_ASAP7_75t_SL g157495 (.A(n_78041),
    .B(n_37355),
    .Y(n_2113));
 NAND2xp5_ASAP7_75t_SL g157500 (.A(n_49620),
    .B(n_50293),
    .Y(n_2503));
 INVxp33_ASAP7_75t_R g157512 (.A(n_1894),
    .Y(n_1895));
 O2A1O1Ixp33_ASAP7_75t_R g157513 (.A1(n_635),
    .A2(u2_cnt[4]),
    .B(n_1645),
    .C(u2_cnt[7]),
    .Y(n_1646));
 NAND2xp5_ASAP7_75t_SL g157516 (.A(n_37368),
    .B(n_78810),
    .Y(n_2108));
 NAND2xp5_ASAP7_75t_SL g157525 (.A(n_78810),
    .B(n_37355),
    .Y(n_2098));
 NAND2xp5_ASAP7_75t_SL g157529 (.A(n_78810),
    .B(n_46642),
    .Y(n_2092));
 NAND2xp5_ASAP7_75t_SL g157546 (.A(n_24350),
    .B(n_13547),
    .Y(n_2074));
 XOR2xp5_ASAP7_75t_L g157547 (.A(n_50088),
    .B(n_47540),
    .Y(n_2073));
 OAI21xp33_ASAP7_75t_SL g157551 (.A1(n_247),
    .A2(n_64715),
    .B(n_1917),
    .Y(n_2164));
 OAI21xp33_ASAP7_75t_SL g157554 (.A1(n_4028),
    .A2(n_640),
    .B(n_40421),
    .Y(n_2162));
 OAI21xp33_ASAP7_75t_SL g157559 (.A1(n_34),
    .A2(n_10613),
    .B(n_8246),
    .Y(n_1888));
 OAI21xp33_ASAP7_75t_L g157561 (.A1(n_75),
    .A2(n_10613),
    .B(n_6721),
    .Y(n_1887));
 OAI21xp5_ASAP7_75t_L g157566 (.A1(n_2),
    .A2(n_10613),
    .B(n_6616),
    .Y(n_1885));
 NAND2xp33_ASAP7_75t_L g157567 (.A(n_36528),
    .B(n_15491),
    .Y(n_2059));
 NAND2xp5_ASAP7_75t_SL g157569 (.A(n_36528),
    .B(n_65293),
    .Y(n_2057));
 AOI211xp5_ASAP7_75t_R g157570 (.A1(n_2290),
    .A2(u2_cnt[3]),
    .B(n_1284),
    .C(n_2467),
    .Y(n_2464));
 NAND2xp5_ASAP7_75t_L g157575 (.A(n_36528),
    .B(n_57289),
    .Y(n_2053));
 NAND2xp5_ASAP7_75t_SL g157577 (.A(n_65578),
    .B(n_36528),
    .Y(n_2052));
 AOI211xp5_ASAP7_75t_R g157579 (.A1(n_2288),
    .A2(u2_cnt[1]),
    .B(n_1193),
    .C(n_2465),
    .Y(n_2466));
 O2A1O1Ixp33_ASAP7_75t_R g157580 (.A1(n_655),
    .A2(u2_cnt[2]),
    .B(n_2290),
    .C(n_2467),
    .Y(n_2291));
 NAND5xp2_ASAP7_75t_R g157581 (.A(n_528),
    .B(n_1088),
    .C(n_1193),
    .D(n_1903),
    .E(u2_cnt[6]),
    .Y(n_1089));
 AOI221xp5_ASAP7_75t_R g157583 (.A1(n_736),
    .A2(u2_cnt[4]),
    .B1(n_737),
    .B2(n_1914),
    .C(n_2467),
    .Y(n_2468));
 NOR2xp33_ASAP7_75t_SL g157589 (.A(n_27061),
    .B(n_700),
    .Y(n_2155));
 NOR2xp33_ASAP7_75t_SL g157596 (.A(n_1808),
    .B(n_1775),
    .Y(n_2149));
 AOI221xp5_ASAP7_75t_SL g157597 (.A1(n_24512),
    .A2(\u3_mem[0] [31]),
    .B1(\u3_mem[1] [31]),
    .B2(n_24513),
    .C(n_1794),
    .Y(n_2230));
 NOR2xp33_ASAP7_75t_SL g157602 (.A(n_1768),
    .B(n_1965),
    .Y(n_2232));
 NOR2xp33_ASAP7_75t_SL g157605 (.A(n_1764),
    .B(n_1990),
    .Y(n_2234));
 NOR2xp67_ASAP7_75t_SL g157606 (.A(n_1785),
    .B(n_6232),
    .Y(n_2143));
 NAND2xp5_ASAP7_75t_SL g157628 (.A(n_14108),
    .B(n_1932),
    .Y(n_2578));
 OAI21xp5_ASAP7_75t_SL g157630 (.A1(n_29953),
    .A2(n_1310),
    .B(n_79203),
    .Y(n_2345));
 NAND2xp5_ASAP7_75t_L g157634 (.A(n_2013),
    .B(n_67490),
    .Y(n_2016));
 NAND3xp33_ASAP7_75t_R g157636 (.A(n_1535),
    .B(u2_cnt[4]),
    .C(n_2119),
    .Y(n_1894));
 NAND2xp5_ASAP7_75t_L g157637 (.A(n_2013),
    .B(n_70887),
    .Y(n_2014));
 NAND2xp5_ASAP7_75t_SL g157639 (.A(n_71352),
    .B(n_2013),
    .Y(n_2009));
 NAND2xp5_ASAP7_75t_SL g157640 (.A(n_65578),
    .B(n_2013),
    .Y(n_2446));
 NAND2xp5_ASAP7_75t_SL g157641 (.A(n_573),
    .B(n_46334),
    .Y(n_2174));
 NAND2xp5_ASAP7_75t_SL g157642 (.A(n_57289),
    .B(n_2013),
    .Y(n_2444));
 NAND2xp5_ASAP7_75t_SL g157643 (.A(n_79203),
    .B(n_15491),
    .Y(n_2434));
 NAND2xp5_ASAP7_75t_SL g157644 (.A(n_573),
    .B(n_50344),
    .Y(n_2176));
 NAND2xp5_ASAP7_75t_SL g157646 (.A(n_79193),
    .B(n_48974),
    .Y(n_2432));
 NAND2xp5_ASAP7_75t_SL g157649 (.A(n_34645),
    .B(n_666),
    .Y(n_2500));
 NAND2xp5_ASAP7_75t_SL g157653 (.A(n_1836),
    .B(n_666),
    .Y(n_2401));
 NAND2xp5_ASAP7_75t_SL g157654 (.A(n_1844),
    .B(n_666),
    .Y(n_2403));
 NAND2xp5_ASAP7_75t_SL g157655 (.A(n_50293),
    .B(n_1842),
    .Y(n_2540));
 NAND2xp5_ASAP7_75t_SL g157656 (.A(n_50293),
    .B(n_1840),
    .Y(n_2511));
 NAND2xp5_ASAP7_75t_SL g157659 (.A(n_28327),
    .B(n_78041),
    .Y(n_1999));
 NAND2xp5_ASAP7_75t_L g157662 (.A(n_50293),
    .B(n_1831),
    .Y(n_2508));
 NAND2xp33_ASAP7_75t_R g157670 (.A(u2_cnt[5]),
    .B(n_1841),
    .Y(n_2330));
 INVx1_ASAP7_75t_SL g157675 (.A(n_1836),
    .Y(n_2384));
 INVx1_ASAP7_75t_SL g157676 (.A(n_36107),
    .Y(n_2424));
 INVxp33_ASAP7_75t_SL g157677 (.A(n_49620),
    .Y(n_1872));
 INVx1_ASAP7_75t_L g157678 (.A(n_28370),
    .Y(n_4428));
 INVx1_ASAP7_75t_SL g157687 (.A(n_36383),
    .Y(n_2375));
 INVxp67_ASAP7_75t_SL g157688 (.A(n_1831),
    .Y(n_2498));
 INVxp67_ASAP7_75t_SL g157694 (.A(n_36525),
    .Y(n_1742));
 INVx1_ASAP7_75t_SL g157697 (.A(n_21015),
    .Y(n_4332));
 INVx1_ASAP7_75t_SL g157700 (.A(n_14108),
    .Y(n_2393));
 INVxp33_ASAP7_75t_SL g157701 (.A(n_59477),
    .Y(n_1739));
 INVxp67_ASAP7_75t_L g157709 (.A(n_34203),
    .Y(n_1853));
 INVxp67_ASAP7_75t_SL g157714 (.A(n_28327),
    .Y(n_4416));
 INVxp33_ASAP7_75t_SL g157717 (.A(n_26733),
    .Y(n_1847));
 INVx1_ASAP7_75t_SL g157718 (.A(n_13547),
    .Y(n_4568));
 INVxp33_ASAP7_75t_L g157723 (.A(n_53003),
    .Y(n_1955));
 INVx1_ASAP7_75t_SL g157725 (.A(n_1844),
    .Y(n_2427));
 INVxp33_ASAP7_75t_SL g157726 (.A(n_34645),
    .Y(n_1736));
 INVxp67_ASAP7_75t_SL g157727 (.A(n_34190),
    .Y(n_4422));
 INVxp33_ASAP7_75t_SL g157732 (.A(n_35407),
    .Y(n_1845));
 INVx1_ASAP7_75t_L g157735 (.A(n_47552),
    .Y(n_4381));
 INVxp67_ASAP7_75t_SL g157736 (.A(n_31107),
    .Y(n_4424));
 INVx1_ASAP7_75t_SL g157740 (.A(n_18709),
    .Y(n_4377));
 INVxp33_ASAP7_75t_SL g157741 (.A(n_57289),
    .Y(n_1846));
 INVxp33_ASAP7_75t_SL g157743 (.A(n_40287),
    .Y(n_1957));
 INVxp33_ASAP7_75t_SL g157744 (.A(n_48729),
    .Y(n_1959));
 INVx1_ASAP7_75t_SL g157747 (.A(n_1838),
    .Y(n_2440));
 INVxp67_ASAP7_75t_SL g157748 (.A(n_48974),
    .Y(n_1849));
 INVxp67_ASAP7_75t_SL g157749 (.A(n_31445),
    .Y(n_4324));
 INVx1_ASAP7_75t_SL g157751 (.A(n_50344),
    .Y(n_4357));
 INVxp67_ASAP7_75t_SL g157752 (.A(n_15491),
    .Y(n_1734));
 INVxp67_ASAP7_75t_L g157755 (.A(n_14017),
    .Y(n_1850));
 INVxp67_ASAP7_75t_SL g157758 (.A(n_46642),
    .Y(n_4426));
 INVx1_ASAP7_75t_L g157759 (.A(n_46334),
    .Y(n_4345));
 INVxp67_ASAP7_75t_SL g157760 (.A(n_65578),
    .Y(n_1852));
 INVxp67_ASAP7_75t_SL g157762 (.A(n_16458),
    .Y(n_4355));
 INVxp67_ASAP7_75t_SL g157763 (.A(n_70887),
    .Y(n_4353));
 INVxp67_ASAP7_75t_SL g157765 (.A(n_67490),
    .Y(n_4350));
 INVxp33_ASAP7_75t_R g157766 (.A(u1_sr[2]),
    .Y(n_2292));
 INVxp33_ASAP7_75t_R g157767 (.A(n_2138),
    .Y(n_2465));
 INVxp33_ASAP7_75t_R g157769 (.A(n_2467),
    .Y(n_2138));
 BUFx3_ASAP7_75t_SL g157770 (.A(u13_csr[1]),
    .Y(n_2467));
 NAND2xp5_ASAP7_75t_SL g157774 (.A(n_42621),
    .B(n_8175),
    .Y(n_1857));
 NAND2xp5_ASAP7_75t_SL g157776 (.A(n_21111),
    .B(n_11559),
    .Y(n_1635));
 NAND2xp5_ASAP7_75t_SL g157777 (.A(n_46260),
    .B(n_11585),
    .Y(n_1634));
 NAND2xp5_ASAP7_75t_SL g157778 (.A(n_21109),
    .B(n_11580),
    .Y(n_1633));
 NAND2xp5_ASAP7_75t_SL g157779 (.A(n_21096),
    .B(n_11555),
    .Y(n_1632));
 NAND2xp5_ASAP7_75t_SL g157780 (.A(n_21095),
    .B(n_11572),
    .Y(n_1631));
 NAND2xp5_ASAP7_75t_SL g157781 (.A(n_21119),
    .B(n_11560),
    .Y(n_1630));
 NAND2xp5_ASAP7_75t_SL g157782 (.A(n_32411),
    .B(n_11648),
    .Y(n_1629));
 NAND2xp5_ASAP7_75t_SL g157783 (.A(n_32385),
    .B(n_11622),
    .Y(n_1628));
 NAND2xp5_ASAP7_75t_SL g157784 (.A(n_32389),
    .B(n_11638),
    .Y(n_1627));
 NAND2xp5_ASAP7_75t_SL g157785 (.A(n_32387),
    .B(n_11650),
    .Y(n_1626));
 NAND2xp5_ASAP7_75t_SL g157786 (.A(n_32393),
    .B(n_11641),
    .Y(n_1625));
 NAND2xp5_ASAP7_75t_SL g157787 (.A(n_32402),
    .B(n_11642),
    .Y(n_1624));
 NAND2xp5_ASAP7_75t_SL g157788 (.A(n_32399),
    .B(n_11637),
    .Y(n_1623));
 NAND2xp5_ASAP7_75t_SL g157789 (.A(n_9703),
    .B(n_11636),
    .Y(n_1622));
 NAND2xp5_ASAP7_75t_SL g157790 (.A(n_32409),
    .B(n_11635),
    .Y(n_1621));
 NAND2xp5_ASAP7_75t_SL g157791 (.A(n_32395),
    .B(n_11644),
    .Y(n_1531));
 NAND2xp5_ASAP7_75t_SL g157792 (.A(n_32408),
    .B(n_11634),
    .Y(n_1620));
 NAND2xp5_ASAP7_75t_SL g157793 (.A(n_32384),
    .B(n_11621),
    .Y(n_1619));
 NAND2xp5_ASAP7_75t_SL g157794 (.A(n_32406),
    .B(n_11646),
    .Y(n_1618));
 NAND2xp5_ASAP7_75t_SL g157795 (.A(n_32404),
    .B(n_11645),
    .Y(n_1617));
 NAND2xp5_ASAP7_75t_SL g157796 (.A(n_9686),
    .B(n_11647),
    .Y(n_1616));
 NAND2xp5_ASAP7_75t_SL g157797 (.A(n_32386),
    .B(n_11620),
    .Y(n_1615));
 NAND2xp5_ASAP7_75t_SL g157798 (.A(n_32410),
    .B(n_11632),
    .Y(n_1614));
 NAND2xp5_ASAP7_75t_SL g157799 (.A(n_32383),
    .B(n_11619),
    .Y(n_1530));
 NAND2xp5_ASAP7_75t_SL g157800 (.A(n_32392),
    .B(n_11631),
    .Y(n_1613));
 NAND2xp5_ASAP7_75t_SL g157801 (.A(n_9682),
    .B(n_11649),
    .Y(n_1612));
 NAND2xp5_ASAP7_75t_SL g157802 (.A(n_32403),
    .B(n_11630),
    .Y(n_1611));
 NAND2xp5_ASAP7_75t_SL g157803 (.A(n_21094),
    .B(n_11564),
    .Y(n_1610));
 NAND2xp5_ASAP7_75t_SL g157804 (.A(n_32391),
    .B(n_11623),
    .Y(n_1609));
 NAND2xp5_ASAP7_75t_SL g157805 (.A(n_9701),
    .B(n_11629),
    .Y(n_1608));
 NAND2xp5_ASAP7_75t_SL g157806 (.A(n_32396),
    .B(n_11639),
    .Y(n_1607));
 NAND2xp5_ASAP7_75t_SL g157807 (.A(n_32394),
    .B(n_11628),
    .Y(n_1606));
 NAND2xp5_ASAP7_75t_SL g157808 (.A(n_32405),
    .B(n_11627),
    .Y(n_1605));
 NAND2xp5_ASAP7_75t_SL g157809 (.A(n_32407),
    .B(n_11626),
    .Y(n_1604));
 NAND2xp5_ASAP7_75t_SL g157810 (.A(n_32398),
    .B(n_11625),
    .Y(n_1603));
 NAND2xp5_ASAP7_75t_SL g157811 (.A(n_32388),
    .B(n_11624),
    .Y(n_1602));
 NAND2xp5_ASAP7_75t_SL g157812 (.A(n_32390),
    .B(n_11633),
    .Y(n_1601));
 NAND2xp5_ASAP7_75t_SL g157813 (.A(n_32400),
    .B(n_11640),
    .Y(n_1600));
 NAND2xp5_ASAP7_75t_SL g157814 (.A(n_21107),
    .B(n_11570),
    .Y(n_1599));
 NAND2xp5_ASAP7_75t_SL g157815 (.A(n_21103),
    .B(n_11576),
    .Y(n_1598));
 NAND2xp5_ASAP7_75t_SL g157816 (.A(n_21122),
    .B(n_11550),
    .Y(n_1597));
 NAND2xp5_ASAP7_75t_SL g157817 (.A(n_21098),
    .B(n_11566),
    .Y(n_1596));
 NAND2xp5_ASAP7_75t_SL g157818 (.A(n_21124),
    .B(n_11575),
    .Y(n_1595));
 NAND2xp5_ASAP7_75t_SL g157819 (.A(n_21112),
    .B(n_11579),
    .Y(n_1594));
 NAND2xp5_ASAP7_75t_SL g157820 (.A(n_21121),
    .B(n_11561),
    .Y(n_1593));
 NAND2xp5_ASAP7_75t_SL g157821 (.A(n_21118),
    .B(n_11558),
    .Y(n_1592));
 NAND2xp5_ASAP7_75t_SL g157822 (.A(n_21106),
    .B(n_11554),
    .Y(n_1591));
 NAND2xp5_ASAP7_75t_SL g157824 (.A(n_21114),
    .B(n_11578),
    .Y(n_1590));
 NAND2xp5_ASAP7_75t_SL g157825 (.A(n_46258),
    .B(n_11611),
    .Y(n_1589));
 NAND2xp5_ASAP7_75t_SL g157826 (.A(n_21099),
    .B(n_11577),
    .Y(n_1588));
 NAND2xp5_ASAP7_75t_SL g157827 (.A(n_21123),
    .B(n_11562),
    .Y(n_1587));
 NAND2xp5_ASAP7_75t_SL g157828 (.A(n_21120),
    .B(n_11567),
    .Y(n_1586));
 NAND2xp5_ASAP7_75t_SL g157829 (.A(n_46246),
    .B(n_11609),
    .Y(n_1585));
 NAND2xp5_ASAP7_75t_SL g157830 (.A(n_46253),
    .B(n_11589),
    .Y(n_1584));
 NAND2xp5_ASAP7_75t_SL g157831 (.A(n_46239),
    .B(n_11590),
    .Y(n_1583));
 NAND2xp5_ASAP7_75t_SL g157832 (.A(n_46241),
    .B(n_11612),
    .Y(n_1582));
 NAND2xp5_ASAP7_75t_SL g157833 (.A(n_46245),
    .B(n_11593),
    .Y(n_1581));
 NAND2xp5_ASAP7_75t_SL g157834 (.A(n_46250),
    .B(n_11608),
    .Y(n_1580));
 NAND2xp5_ASAP7_75t_SL g157835 (.A(n_46263),
    .B(n_11584),
    .Y(n_1579));
 NAND2xp5_ASAP7_75t_SL g157836 (.A(n_46243),
    .B(n_11594),
    .Y(n_1578));
 NAND2xp5_ASAP7_75t_SL g157837 (.A(n_46237),
    .B(n_11607),
    .Y(n_1577));
 NAND2xp5_ASAP7_75t_SL g157838 (.A(n_46240),
    .B(n_11597),
    .Y(n_1576));
 NAND2xp5_ASAP7_75t_SL g157839 (.A(n_46242),
    .B(n_11606),
    .Y(n_1575));
 NAND2xp5_ASAP7_75t_SL g157840 (.A(n_9663),
    .B(n_11592),
    .Y(n_1574));
 NAND2xp5_ASAP7_75t_SL g157841 (.A(n_21100),
    .B(n_11553),
    .Y(n_1573));
 NAND2xp5_ASAP7_75t_SL g157842 (.A(n_46251),
    .B(n_11615),
    .Y(n_1572));
 NAND2xp5_ASAP7_75t_SL g157843 (.A(n_46236),
    .B(n_11588),
    .Y(n_1571));
 NAND2xp5_ASAP7_75t_SL g157844 (.A(n_9654),
    .B(n_11613),
    .Y(n_1570));
 NAND2xp5_ASAP7_75t_SL g157845 (.A(n_46254),
    .B(n_11602),
    .Y(n_1569));
 NAND2xp5_ASAP7_75t_SL g157846 (.A(n_46259),
    .B(n_11605),
    .Y(n_1568));
 NAND2xp5_ASAP7_75t_SL g157847 (.A(n_46244),
    .B(n_11599),
    .Y(n_1567));
 NAND2xp5_ASAP7_75t_SL g157848 (.A(n_46262),
    .B(n_11587),
    .Y(n_1566));
 NAND2xp5_ASAP7_75t_SL g157849 (.A(n_46247),
    .B(n_11603),
    .Y(n_1565));
 NAND2xp5_ASAP7_75t_SL g157850 (.A(n_46249),
    .B(n_11595),
    .Y(n_1564));
 NAND2xp5_ASAP7_75t_SL g157851 (.A(n_9650),
    .B(n_11596),
    .Y(n_1563));
 NAND2xp5_ASAP7_75t_SL g157852 (.A(n_46257),
    .B(n_11614),
    .Y(n_1660));
 NAND2xp5_ASAP7_75t_SL g157853 (.A(n_46256),
    .B(n_11610),
    .Y(n_1561));
 NAND2xp5_ASAP7_75t_SL g157854 (.A(n_21116),
    .B(n_11569),
    .Y(n_1560));
 NAND2xp5_ASAP7_75t_SL g157855 (.A(n_46261),
    .B(n_11586),
    .Y(n_1559));
 NAND3xp33_ASAP7_75t_SL g157856 (.A(n_27257),
    .B(n_28955),
    .C(n_1058),
    .Y(n_1558));
 NAND2xp5_ASAP7_75t_SL g157857 (.A(n_46248),
    .B(n_11600),
    .Y(n_1555));
 NAND2xp5_ASAP7_75t_SL g157858 (.A(n_21108),
    .B(n_11557),
    .Y(n_1554));
 NAND2xp5_ASAP7_75t_SL g157859 (.A(n_46252),
    .B(n_11604),
    .Y(n_1553));
 NAND2xp5_ASAP7_75t_SL g157860 (.A(n_21102),
    .B(n_11552),
    .Y(n_1552));
 NAND2xp5_ASAP7_75t_SL g157861 (.A(n_21110),
    .B(n_11565),
    .Y(n_1551));
 NAND2xp5_ASAP7_75t_SL g157862 (.A(n_46255),
    .B(n_11591),
    .Y(n_1550));
 NAND2xp5_ASAP7_75t_SL g157863 (.A(n_21117),
    .B(n_11573),
    .Y(n_1549));
 NAND2xp5_ASAP7_75t_SL g157864 (.A(n_9665),
    .B(n_11598),
    .Y(n_1548));
 NAND2xp5_ASAP7_75t_L g157865 (.A(n_468),
    .B(n_597),
    .Y(n_778));
 NAND2xp5_ASAP7_75t_SL g157866 (.A(n_32401),
    .B(n_11643),
    .Y(n_1547));
 NAND2xp5_ASAP7_75t_SL g157867 (.A(n_21104),
    .B(n_11574),
    .Y(n_1546));
 NAND2xp5_ASAP7_75t_SL g157868 (.A(n_21113),
    .B(n_11571),
    .Y(n_1545));
 NAND2xp5_ASAP7_75t_SL g157869 (.A(n_21101),
    .B(n_11556),
    .Y(n_1544));
 NAND2xp5_ASAP7_75t_SL g157871 (.A(n_21097),
    .B(n_11551),
    .Y(n_1540));
 NAND2xp5_ASAP7_75t_SL g157874 (.A(n_21105),
    .B(n_11563),
    .Y(n_1637));
 NAND2xp33_ASAP7_75t_SL g157875 (.A(n_1306),
    .B(u2_to_cnt[4]),
    .Y(n_1861));
 NAND2xp5_ASAP7_75t_SL g157892 (.A(n_51053),
    .B(n_19496),
    .Y(n_1836));
 AND2x2_ASAP7_75t_SL g157898 (.A(n_56863),
    .B(n_31900),
    .Y(n_4316));
 NAND2xp5_ASAP7_75t_SL g157899 (.A(n_1261),
    .B(n_33790),
    .Y(n_1968));
 NAND2xp5_ASAP7_75t_SL g157906 (.A(n_19506),
    .B(n_51047),
    .Y(n_1831));
 AND2x2_ASAP7_75t_SL g157907 (.A(n_7411),
    .B(n_6065),
    .Y(n_4405));
 NAND2x1_ASAP7_75t_SL g157913 (.A(n_1033),
    .B(n_798),
    .Y(n_1828));
 AND2x2_ASAP7_75t_SL g157921 (.A(n_1145),
    .B(n_1040),
    .Y(n_4540));
 AND2x2_ASAP7_75t_SL g157945 (.A(n_51038),
    .B(n_6301),
    .Y(n_4448));
 NAND2x1_ASAP7_75t_SL g157947 (.A(n_33789),
    .B(n_7410),
    .Y(n_4515));
 NAND2xp5_ASAP7_75t_SL g157948 (.A(n_19504),
    .B(n_51046),
    .Y(n_1840));
 NAND2xp5_ASAP7_75t_SL g157950 (.A(n_19505),
    .B(n_51049),
    .Y(n_1842));
 NAND2xp5_ASAP7_75t_SL g157951 (.A(n_51040),
    .B(n_19497),
    .Y(n_1844));
 NAND2xp5_ASAP7_75t_SL g157970 (.A(n_51482),
    .B(n_7542),
    .Y(n_1723));
 NAND2xp5_ASAP7_75t_SL g157971 (.A(n_51495),
    .B(n_7543),
    .Y(n_1838));
 AND2x2_ASAP7_75t_SL g157975 (.A(n_13989),
    .B(n_51486),
    .Y(n_4341));
 AND2x2_ASAP7_75t_SL g157978 (.A(n_51489),
    .B(n_7541),
    .Y(n_4339));
 AND2x2_ASAP7_75t_SL g157991 (.A(n_56849),
    .B(n_7881),
    .Y(n_4320));
 AOI22xp5_ASAP7_75t_SL g158 (.A1(\u8_mem[0] [10]),
    .A2(n_59474),
    .B1(\u8_mem[1] [10]),
    .B2(n_78274),
    .Y(n_71351));
 INVx1_ASAP7_75t_L g158000 (.A(n_35550),
    .Y(n_4343));
 INVxp67_ASAP7_75t_SL g158003 (.A(n_2168),
    .Y(n_4346));
 NAND2xp5_ASAP7_75t_SL g158006 (.A(n_21115),
    .B(n_11568),
    .Y(n_1519));
 NAND2xp5_ASAP7_75t_SL g158008 (.A(n_46238),
    .B(n_11601),
    .Y(n_1516));
 NAND4xp25_ASAP7_75t_SL g158009 (.A(n_490),
    .B(n_443),
    .C(n_461),
    .D(n_454),
    .Y(n_1086));
 NAND4xp25_ASAP7_75t_SL g158011 (.A(n_442),
    .B(n_451),
    .C(n_462),
    .D(n_467),
    .Y(n_1084));
 A2O1A1Ixp33_ASAP7_75t_R g158013 (.A1(u2_cnt[1]),
    .A2(n_1088),
    .B(u2_cnt[4]),
    .C(u2_cnt[6]),
    .Y(n_1330));
 NOR4xp25_ASAP7_75t_R g158015 (.A(n_1661),
    .B(u12_we2),
    .C(wb_addr_i[5]),
    .D(wb_addr_i[6]),
    .Y(n_1869));
 NOR3xp33_ASAP7_75t_R g158017 (.A(n_1082),
    .B(u2_cnt[6]),
    .C(u2_cnt[4]),
    .Y(n_1083));
 NAND3xp33_ASAP7_75t_R g158018 (.A(n_1336),
    .B(n_714),
    .C(n_1645),
    .Y(n_1510));
 AOI22xp33_ASAP7_75t_L g158036 (.A1(oc2_cfg[6]),
    .A2(n_8212),
    .B1(u13_intm_r[22]),
    .B2(n_7082),
    .Y(n_1490));
 OAI21xp5_ASAP7_75t_SL g158038 (.A1(n_6960),
    .A2(n_72),
    .B(n_1287),
    .Y(n_1896));
 AOI22xp33_ASAP7_75t_L g158039 (.A1(crac_out[31]),
    .A2(n_22851),
    .B1(n_6961),
    .B2(u13_occ0_r[31]),
    .Y(n_1329));
 AOI22xp5_ASAP7_75t_SL g158040 (.A1(oc3_cfg[2]),
    .A2(n_8212),
    .B1(u13_intm_r[26]),
    .B2(n_7082),
    .Y(n_1488));
 AOI22xp33_ASAP7_75t_L g158044 (.A1(oc2_cfg[5]),
    .A2(n_8212),
    .B1(u13_intm_r[21]),
    .B2(n_7082),
    .Y(n_1484));
 AOI22xp33_ASAP7_75t_L g158045 (.A1(oc2_cfg[1]),
    .A2(n_6961),
    .B1(u13_intm_r[17]),
    .B2(n_7083),
    .Y(n_1483));
 AOI22xp33_ASAP7_75t_SL g158052 (.A1(oc3_cfg[1]),
    .A2(n_8212),
    .B1(u13_intm_r[25]),
    .B2(n_7082),
    .Y(n_1475));
 AOI22xp33_ASAP7_75t_L g158057 (.A1(oc3_cfg[0]),
    .A2(n_6961),
    .B1(n_227),
    .B2(n_7084),
    .Y(n_1470));
 OAI22xp33_ASAP7_75t_SL g158065 (.A1(n_1372),
    .A2(u7_rp[0]),
    .B1(n_419),
    .B2(n_29364),
    .Y(n_1917));
 OAI21xp33_ASAP7_75t_SL g158070 (.A1(n_59339),
    .A2(n_69),
    .B(n_1288),
    .Y(n_1816));
 OAI22xp33_ASAP7_75t_SL g158071 (.A1(n_17623),
    .A2(n_24),
    .B1(n_23530),
    .B2(n_137),
    .Y(n_1965));
 AOI22xp33_ASAP7_75t_R g158072 (.A1(\u5_mem[2] [22]),
    .A2(n_1459),
    .B1(\u5_mem[3] [22]),
    .B2(n_56865),
    .Y(n_1461));
 AOI22xp33_ASAP7_75t_R g158073 (.A1(\u5_mem[2] [23]),
    .A2(n_1459),
    .B1(\u5_mem[3] [23]),
    .B2(n_56865),
    .Y(n_1460));
 AOI22xp33_ASAP7_75t_L g158074 (.A1(\u5_mem[2] [24]),
    .A2(n_1459),
    .B1(\u5_mem[3] [24]),
    .B2(n_56865),
    .Y(n_1457));
 AOI22xp33_ASAP7_75t_R g158075 (.A1(\u5_mem[2] [25]),
    .A2(n_1459),
    .B1(\u5_mem[3] [25]),
    .B2(n_56865),
    .Y(n_1456));
 AOI22xp5_ASAP7_75t_R g158076 (.A1(\u5_mem[2] [27]),
    .A2(n_1459),
    .B1(\u5_mem[3] [27]),
    .B2(n_56865),
    .Y(n_1455));
 AOI22xp33_ASAP7_75t_L g158081 (.A1(\u4_mem[2] [29]),
    .A2(n_17624),
    .B1(\u4_mem[3] [29]),
    .B2(n_23531),
    .Y(n_1812));
 AOI22xp33_ASAP7_75t_SL g158082 (.A1(\u4_mem[2] [24]),
    .A2(n_17624),
    .B1(\u4_mem[3] [24]),
    .B2(n_23531),
    .Y(n_1809));
 AOI22xp33_ASAP7_75t_L g158083 (.A1(\u5_mem[2] [26]),
    .A2(n_1459),
    .B1(\u5_mem[3] [26]),
    .B2(n_56865),
    .Y(n_1452));
 OAI21xp5_ASAP7_75t_SL g158084 (.A1(n_59339),
    .A2(n_154),
    .B(n_1297),
    .Y(n_1808));
 AOI22xp33_ASAP7_75t_L g158085 (.A1(\u4_mem[2] [27]),
    .A2(n_17624),
    .B1(\u4_mem[3] [27]),
    .B2(n_23531),
    .Y(n_1807));
 OAI22xp33_ASAP7_75t_SL g158087 (.A1(n_62),
    .A2(n_17623),
    .B1(n_23530),
    .B2(n_160),
    .Y(n_1972));
 AOI22xp33_ASAP7_75t_L g158088 (.A1(\u4_mem[2] [22]),
    .A2(n_17624),
    .B1(\u4_mem[3] [22]),
    .B2(n_23531),
    .Y(n_1805));
 OAI22xp33_ASAP7_75t_SL g158090 (.A1(n_111),
    .A2(n_17623),
    .B1(n_23530),
    .B2(n_156),
    .Y(n_1990));
 AOI22xp33_ASAP7_75t_L g158091 (.A1(\u4_mem[2] [31]),
    .A2(n_17624),
    .B1(\u4_mem[3] [31]),
    .B2(n_23531),
    .Y(n_1803));
 AOI22xp33_ASAP7_75t_SL g158092 (.A1(\u4_mem[2] [26]),
    .A2(n_17624),
    .B1(\u4_mem[3] [26]),
    .B2(n_23531),
    .Y(n_1802));
 AOI22xp5_ASAP7_75t_SL g158093 (.A1(\u3_mem[2] [26]),
    .A2(n_77398),
    .B1(\u3_mem[3] [26]),
    .B2(n_22062),
    .Y(n_1801));
 AOI22xp33_ASAP7_75t_L g158095 (.A1(n_77398),
    .A2(\u3_mem[2] [28]),
    .B1(\u3_mem[3] [28]),
    .B2(n_22062),
    .Y(n_1797));
 OAI22xp5_ASAP7_75t_SL g158098 (.A1(n_1783),
    .A2(n_48),
    .B1(n_1782),
    .B2(n_20),
    .Y(n_1794));
 OAI22xp5_ASAP7_75t_SL g158101 (.A1(n_65029),
    .A2(n_84),
    .B1(n_67),
    .B2(n_59256),
    .Y(n_1793));
 OAI22xp5_ASAP7_75t_SL g158103 (.A1(n_65029),
    .A2(n_93),
    .B1(n_71),
    .B2(n_59256),
    .Y(n_1789));
 OAI22xp5_ASAP7_75t_SL g158104 (.A1(n_65029),
    .A2(n_123),
    .B1(n_161),
    .B2(n_59256),
    .Y(n_1788));
 OAI22xp5_ASAP7_75t_SL g158108 (.A1(n_65029),
    .A2(n_55),
    .B1(n_74),
    .B2(n_59256),
    .Y(n_1785));
 AOI22xp33_ASAP7_75t_SL g158111 (.A1(\u8_mem[2] [20]),
    .A2(n_51488),
    .B1(\u8_mem[3] [20]),
    .B2(n_14001),
    .Y(n_1444));
 OAI22xp33_ASAP7_75t_SL g158113 (.A1(n_1783),
    .A2(n_52),
    .B1(n_1782),
    .B2(n_79),
    .Y(n_1784));
 OAI22xp33_ASAP7_75t_L g158114 (.A1(n_1783),
    .A2(n_118),
    .B1(n_1782),
    .B2(n_8),
    .Y(n_1781));
 AOI22xp5_ASAP7_75t_SL g158115 (.A1(\u3_mem[2] [22]),
    .A2(n_77398),
    .B1(\u3_mem[3] [22]),
    .B2(n_22062),
    .Y(n_1780));
 AOI22xp33_ASAP7_75t_SL g158116 (.A1(\u8_mem[2] [21]),
    .A2(n_51488),
    .B1(\u8_mem[3] [21]),
    .B2(n_14001),
    .Y(n_1440));
 AOI22xp5_ASAP7_75t_SL g158117 (.A1(\u3_mem[2] [23]),
    .A2(n_77398),
    .B1(\u3_mem[3] [23]),
    .B2(n_22062),
    .Y(n_1779));
 AOI22xp33_ASAP7_75t_L g158118 (.A1(\u8_mem[2] [22]),
    .A2(n_51488),
    .B1(n_14001),
    .B2(\u8_mem[3] [22]),
    .Y(n_1439));
 AOI22xp33_ASAP7_75t_L g158120 (.A1(\u8_mem[2] [25]),
    .A2(n_51488),
    .B1(\u8_mem[3] [25]),
    .B2(n_14001),
    .Y(n_1437));
 AOI22xp33_ASAP7_75t_R g158122 (.A1(\u8_mem[2] [27]),
    .A2(n_51488),
    .B1(\u8_mem[3] [27]),
    .B2(n_14001),
    .Y(n_1436));
 AOI22xp33_ASAP7_75t_L g158123 (.A1(\u8_mem[2] [28]),
    .A2(n_51488),
    .B1(\u8_mem[3] [28]),
    .B2(n_14001),
    .Y(n_1435));
 AOI22xp33_ASAP7_75t_L g158124 (.A1(\u8_mem[2] [24]),
    .A2(n_51488),
    .B1(\u8_mem[3] [24]),
    .B2(n_14001),
    .Y(n_1434));
 AOI22xp33_ASAP7_75t_L g158125 (.A1(\u8_mem[2] [29]),
    .A2(n_51488),
    .B1(\u8_mem[3] [29]),
    .B2(n_14001),
    .Y(n_1433));
 AOI22xp33_ASAP7_75t_SL g158126 (.A1(\u8_mem[2] [30]),
    .A2(n_51488),
    .B1(\u8_mem[3] [30]),
    .B2(n_14001),
    .Y(n_1432));
 AOI22xp5_ASAP7_75t_SL g158128 (.A1(n_77398),
    .A2(\u3_mem[2] [25]),
    .B1(\u3_mem[3] [25]),
    .B2(n_22062),
    .Y(n_1777));
 AOI22xp33_ASAP7_75t_L g158129 (.A1(\u6_mem[1] [23]),
    .A2(n_48415),
    .B1(\u6_mem[3] [23]),
    .B2(n_17704),
    .Y(n_1430));
 AOI22xp33_ASAP7_75t_SL g158131 (.A1(\u6_mem[1] [20]),
    .A2(n_48415),
    .B1(\u6_mem[3] [20]),
    .B2(n_17704),
    .Y(n_1426));
 AOI22xp33_ASAP7_75t_L g158135 (.A1(\u6_mem[1] [28]),
    .A2(n_48415),
    .B1(\u6_mem[3] [28]),
    .B2(n_17704),
    .Y(n_1422));
 AOI22xp33_ASAP7_75t_L g158136 (.A1(\u6_mem[1] [30]),
    .A2(n_48415),
    .B1(\u6_mem[3] [30]),
    .B2(n_17704),
    .Y(n_1421));
 AOI22xp33_ASAP7_75t_L g158137 (.A1(\u6_mem[1] [31]),
    .A2(n_48415),
    .B1(\u6_mem[3] [31]),
    .B2(n_17704),
    .Y(n_1420));
 AOI22xp33_ASAP7_75t_L g158139 (.A1(n_48415),
    .A2(\u6_mem[1] [22]),
    .B1(\u6_mem[3] [22]),
    .B2(n_17704),
    .Y(n_1418));
 OAI22xp33_ASAP7_75t_SL g158142 (.A1(n_89),
    .A2(n_64994),
    .B1(n_7),
    .B2(n_64993),
    .Y(n_1775));
 AOI22xp33_ASAP7_75t_SL g158144 (.A1(n_64793),
    .A2(\u5_mem[0] [23]),
    .B1(n_6071),
    .B2(\u5_mem[1] [23]),
    .Y(n_1992));
 OAI22xp5_ASAP7_75t_SL g158148 (.A1(n_9),
    .A2(n_64994),
    .B1(n_3),
    .B2(n_64993),
    .Y(n_1770));
 OAI22xp5_ASAP7_75t_SL g158149 (.A1(n_51),
    .A2(n_64994),
    .B1(n_149),
    .B2(n_64993),
    .Y(n_1769));
 OAI22xp33_ASAP7_75t_SL g158152 (.A1(n_21),
    .A2(n_36011),
    .B1(n_58),
    .B2(n_1762),
    .Y(n_1768));
 AOI22xp33_ASAP7_75t_SL g158153 (.A1(\u4_mem[0] [27]),
    .A2(n_1766),
    .B1(\u4_mem[1] [27]),
    .B2(n_1765),
    .Y(n_1767));
 OAI22xp33_ASAP7_75t_SL g158154 (.A1(n_66),
    .A2(n_36011),
    .B1(n_37),
    .B2(n_1762),
    .Y(n_1764));
 OAI22xp33_ASAP7_75t_SL g158156 (.A1(n_94),
    .A2(n_36011),
    .B1(n_144),
    .B2(n_1762),
    .Y(n_1760));
 AOI22xp33_ASAP7_75t_SL g158159 (.A1(\u4_mem[0] [22]),
    .A2(n_1766),
    .B1(\u4_mem[1] [22]),
    .B2(n_1765),
    .Y(n_1757));
 AOI22xp33_ASAP7_75t_SL g158161 (.A1(\u4_mem[0] [29]),
    .A2(n_1766),
    .B1(\u4_mem[1] [29]),
    .B2(n_1765),
    .Y(n_1755));
 AOI22xp33_ASAP7_75t_SL g158162 (.A1(\u4_mem[0] [24]),
    .A2(n_1766),
    .B1(\u4_mem[1] [24]),
    .B2(n_1765),
    .Y(n_1754));
 AOI22xp5_ASAP7_75t_SL g158163 (.A1(\u4_mem[0] [31]),
    .A2(n_1766),
    .B1(\u4_mem[1] [31]),
    .B2(n_1765),
    .Y(n_1753));
 OAI22xp33_ASAP7_75t_L g158164 (.A1(n_64994),
    .A2(n_90),
    .B1(n_134),
    .B2(n_64993),
    .Y(n_1752));
 AOI22xp33_ASAP7_75t_L g158165 (.A1(\u3_mem[0] [26]),
    .A2(n_24512),
    .B1(\u3_mem[1] [26]),
    .B2(n_24513),
    .Y(n_1751));
 AOI22xp5_ASAP7_75t_L g158167 (.A1(\u3_mem[0] [30]),
    .A2(n_24512),
    .B1(\u3_mem[1] [30]),
    .B2(n_24513),
    .Y(n_1749));
 AOI22xp33_ASAP7_75t_L g158171 (.A1(\u6_mem[0] [20]),
    .A2(n_79305),
    .B1(\u6_mem[2] [20]),
    .B2(n_79306),
    .Y(n_1411));
 AOI22xp33_ASAP7_75t_SL g158174 (.A1(n_79305),
    .A2(\u6_mem[0] [23]),
    .B1(\u6_mem[2] [23]),
    .B2(n_79306),
    .Y(n_1406));
 AOI22xp33_ASAP7_75t_L g158177 (.A1(\u6_mem[0] [27]),
    .A2(n_79305),
    .B1(\u6_mem[2] [27]),
    .B2(n_79306),
    .Y(n_1403));
 AOI22xp33_ASAP7_75t_SL g158179 (.A1(\u6_mem[0] [30]),
    .A2(n_79305),
    .B1(\u6_mem[2] [30]),
    .B2(n_79306),
    .Y(n_1401));
 AOI22xp33_ASAP7_75t_SL g158180 (.A1(n_79305),
    .A2(\u6_mem[0] [31]),
    .B1(\u6_mem[2] [31]),
    .B2(n_79306),
    .Y(n_1400));
 AOI22xp33_ASAP7_75t_SL g158189 (.A1(\u3_mem[0] [22]),
    .A2(n_24512),
    .B1(\u3_mem[1] [22]),
    .B2(n_24513),
    .Y(n_1747));
 AOI22xp33_ASAP7_75t_L g158192 (.A1(\u8_mem[0] [20]),
    .A2(n_27133),
    .B1(\u8_mem[1] [20]),
    .B2(n_27134),
    .Y(n_1391));
 AOI22xp33_ASAP7_75t_R g158193 (.A1(\u8_mem[0] [21]),
    .A2(n_27133),
    .B1(\u8_mem[1] [21]),
    .B2(n_27134),
    .Y(n_1390));
 AOI22xp33_ASAP7_75t_L g158194 (.A1(\u8_mem[0] [22]),
    .A2(n_27133),
    .B1(\u8_mem[1] [22]),
    .B2(n_27134),
    .Y(n_1389));
 AOI22xp33_ASAP7_75t_SL g158195 (.A1(\u3_mem[0] [23]),
    .A2(n_24512),
    .B1(\u3_mem[1] [23]),
    .B2(n_24513),
    .Y(n_1745));
 AOI22xp33_ASAP7_75t_L g158197 (.A1(\u8_mem[0] [24]),
    .A2(n_27133),
    .B1(\u8_mem[1] [24]),
    .B2(n_27134),
    .Y(n_1387));
 AOI22xp33_ASAP7_75t_L g158198 (.A1(\u8_mem[0] [25]),
    .A2(n_27133),
    .B1(\u8_mem[1] [25]),
    .B2(n_27134),
    .Y(n_1386));
 AOI22xp33_ASAP7_75t_L g158201 (.A1(\u3_mem[0] [25]),
    .A2(n_24512),
    .B1(n_24513),
    .B2(\u3_mem[1] [25]),
    .Y(n_1744));
 NOR3xp33_ASAP7_75t_R g158216 (.A(n_2290),
    .B(n_1914),
    .C(n_634),
    .Y(n_1841));
 NAND2x1_ASAP7_75t_SL g158227 (.A(n_33793),
    .B(n_7563),
    .Y(n_2168));
 INVx1_ASAP7_75t_SL g158231 (.A(n_7544),
    .Y(n_1310));
 INVx1_ASAP7_75t_SL g158233 (.A(n_23529),
    .Y(n_1892));
 INVxp67_ASAP7_75t_SL g158235 (.A(n_1648),
    .Y(n_1306));
 INVxp67_ASAP7_75t_SL g158238 (.A(n_2458),
    .Y(n_1113));
 INVxp67_ASAP7_75t_SL g158239 (.A(n_19578),
    .Y(n_1343));
 INVxp33_ASAP7_75t_R g158243 (.A(u1_sr[1]),
    .Y(n_2136));
 INVx5_ASAP7_75t_SL g158250_dup (.A(n_10613),
    .Y(n_10626));
 AOI22xp5_ASAP7_75t_SL g158266 (.A1(\u4_mem[0] [19]),
    .A2(n_58959),
    .B1(\u4_mem[1] [19]),
    .B2(n_50709),
    .Y(n_1338));
 NAND2xp5_ASAP7_75t_L g158283 (.A(\u5_mem[3] [21]),
    .B(n_56865),
    .Y(n_1297));
 NOR2xp33_ASAP7_75t_R g158284 (.A(n_53),
    .B(n_1285),
    .Y(n_1296));
 NOR3xp33_ASAP7_75t_R g158288 (.A(n_47541),
    .B(n_19009),
    .C(n_24726),
    .Y(n_1292));
 NOR2xp33_ASAP7_75t_L g158289 (.A(n_178),
    .B(n_1289),
    .Y(n_1290));
 NAND2xp5_ASAP7_75t_R g158292 (.A(\u5_mem[3] [20]),
    .B(n_56865),
    .Y(n_1288));
 NAND2xp5_ASAP7_75t_SL g158293 (.A(n_7086),
    .B(u13_intm_r[1]),
    .Y(n_1287));
 NOR2xp33_ASAP7_75t_L g158294 (.A(n_22),
    .B(n_1285),
    .Y(n_1286));
 NOR2xp33_ASAP7_75t_L g158297 (.A(n_366),
    .B(n_1058),
    .Y(n_1059));
 NOR2xp33_ASAP7_75t_R g158299 (.A(u2_cnt[3]),
    .B(n_2290),
    .Y(n_1284));
 AOI22xp5_ASAP7_75t_SL g158301 (.A1(\u4_mem[0] [5]),
    .A2(n_58959),
    .B1(\u4_mem[1] [5]),
    .B2(n_50709),
    .Y(n_1054));
 AOI31xp33_ASAP7_75t_SL g158302 (.A1(n_274),
    .A2(n_186),
    .A3(n_73),
    .B(u14_u7_en_out_l2),
    .Y(n_709));
 AOI31xp33_ASAP7_75t_SL g158303 (.A1(n_285),
    .A2(n_265),
    .A3(n_113),
    .B(u14_u6_en_out_l2),
    .Y(n_710));
 AOI211xp5_ASAP7_75t_SL g158306 (.A1(oc3_cfg[1]),
    .A2(in_slt1[7]),
    .B(n_57965),
    .C(n_389),
    .Y(n_1051));
 OR4x1_ASAP7_75t_R g158311 (.A(out_slt0[14]),
    .B(out_slt0[13]),
    .C(n_62918),
    .D(n_1042),
    .Y(n_1044));
 AOI22xp5_ASAP7_75t_SL g158312 (.A1(n_58959),
    .A2(\u4_mem[0] [16]),
    .B1(\u4_mem[1] [16]),
    .B2(n_50709),
    .Y(n_1041));
 AOI22xp5_ASAP7_75t_SL g158313 (.A1(\u4_mem[0] [4]),
    .A2(n_58959),
    .B1(\u4_mem[1] [4]),
    .B2(n_50709),
    .Y(n_1040));
 AOI22xp5_ASAP7_75t_SL g158321 (.A1(n_58959),
    .A2(\u4_mem[0] [17]),
    .B1(n_50709),
    .B2(\u4_mem[1] [17]),
    .Y(n_1033));
 AOI22xp5_ASAP7_75t_SL g158322 (.A1(n_58959),
    .A2(\u4_mem[0] [7]),
    .B1(\u4_mem[1] [7]),
    .B2(n_50709),
    .Y(n_1032));
 AOI22xp5_ASAP7_75t_SL g158346 (.A1(n_58959),
    .A2(\u4_mem[0] [6]),
    .B1(\u4_mem[1] [6]),
    .B2(n_50709),
    .Y(n_1017));
 AOI222xp33_ASAP7_75t_SL g158362 (.A1(u13_intm_r[28]),
    .A2(u13_ints_r[28]),
    .B1(u13_intm_r[21]),
    .B2(u13_ints_r[21]),
    .C1(u13_intm_r[0]),
    .C2(u13_ints_r[0]),
    .Y(n_597));
 NAND3xp33_ASAP7_75t_R g158372 (.A(n_528),
    .B(n_1903),
    .C(n_1192),
    .Y(n_529));
 NOR2xp33_ASAP7_75t_R g158464 (.A(u2_cnt[6]),
    .B(n_713),
    .Y(n_1535));
 XNOR2xp5_ASAP7_75t_SL g158466 (.A(n_7656),
    .B(n_267),
    .Y(n_2462));
 NAND2xp5_ASAP7_75t_SL g158469 (.A(n_696),
    .B(n_178),
    .Y(n_1648));
 XNOR2xp5_ASAP7_75t_SL g158472 (.A(n_18897),
    .B(n_18745),
    .Y(n_2458));
 OAI221xp5_ASAP7_75t_SL g158474 (.A1(n_1679),
    .A2(n_34480),
    .B1(n_34484),
    .B2(n_1705),
    .C(n_13247),
    .Y(n_4849));
 OAI221xp5_ASAP7_75t_SL g158477 (.A1(n_1679),
    .A2(n_14313),
    .B1(n_1705),
    .B2(n_21709),
    .C(n_10942),
    .Y(n_4851));
 OAI21xp5_ASAP7_75t_SL g158479 (.A1(n_26831),
    .A2(n_1534),
    .B(n_1528),
    .Y(n_4710));
 OAI21xp5_ASAP7_75t_SL g158516 (.A1(n_26859),
    .A2(n_1534),
    .B(n_1527),
    .Y(n_4712));
 NAND2x1_ASAP7_75t_SL g158517 (.A(n_603),
    .B(u12_we1),
    .Y(n_1661));
 OAI221xp5_ASAP7_75t_SL g158521 (.A1(n_1679),
    .A2(n_36288),
    .B1(n_1705),
    .B2(n_14309),
    .C(n_10943),
    .Y(n_4956));
 OAI221xp5_ASAP7_75t_SL g158527 (.A1(n_1679),
    .A2(n_21705),
    .B1(n_21697),
    .B2(n_1705),
    .C(n_10944),
    .Y(n_4877));
 OAI21xp5_ASAP7_75t_SL g158530 (.A1(n_34480),
    .A2(n_10937),
    .B(n_729),
    .Y(n_4881));
 OAI221xp5_ASAP7_75t_SL g158532 (.A1(n_1679),
    .A2(n_14309),
    .B1(n_1705),
    .B2(n_21705),
    .C(n_13237),
    .Y(n_4869));
 AOI22xp5_ASAP7_75t_SL g158559 (.A1(\u5_mem[0] [0]),
    .A2(n_53101),
    .B1(\u5_mem[2] [0]),
    .B2(n_65643),
    .Y(n_1153));
 AOI22xp5_ASAP7_75t_SL g158576 (.A1(n_58959),
    .A2(\u4_mem[0] [0]),
    .B1(\u4_mem[2] [0]),
    .B2(n_35632),
    .Y(n_933));
 AOI22xp33_ASAP7_75t_SL g158611 (.A1(n_2687),
    .A2(n_71972),
    .B1(u3_rp[3]),
    .B2(n_450),
    .Y(n_908));
 AOI22xp33_ASAP7_75t_SL g158713 (.A1(n_50388),
    .A2(\u3_mem[2] [15]),
    .B1(n_71972),
    .B2(\u3_mem[3] [15]),
    .Y(n_1261));
 AOI22xp5_ASAP7_75t_SL g158721 (.A1(\u4_mem[1] [2]),
    .A2(n_50709),
    .B1(\u4_mem[3] [2]),
    .B2(n_30078),
    .Y(n_811));
 AOI22xp33_ASAP7_75t_SL g158725 (.A1(n_50388),
    .A2(\u3_mem[2] [16]),
    .B1(n_71972),
    .B2(\u3_mem[3] [16]),
    .Y(n_1259));
 AOI22xp5_ASAP7_75t_SL g158728 (.A1(n_35632),
    .A2(\u4_mem[2] [15]),
    .B1(\u4_mem[3] [15]),
    .B2(n_30078),
    .Y(n_805));
 AOI22xp33_ASAP7_75t_SL g158734 (.A1(\u4_mem[2] [5]),
    .A2(n_35632),
    .B1(\u4_mem[3] [5]),
    .B2(n_30078),
    .Y(n_801));
 AOI22xp5_ASAP7_75t_SL g158738 (.A1(\u4_mem[2] [17]),
    .A2(n_35632),
    .B1(\u4_mem[3] [17]),
    .B2(n_30078),
    .Y(n_798));
 AO22x1_ASAP7_75t_SL g158753 (.A1(n_35632),
    .A2(\u4_mem[2] [18]),
    .B1(\u4_mem[3] [18]),
    .B2(n_30078),
    .Y(n_1643));
 AOI22xp5_ASAP7_75t_SL g158758 (.A1(\u4_mem[1] [12]),
    .A2(n_50709),
    .B1(\u4_mem[3] [12]),
    .B2(n_30078),
    .Y(n_782));
 AOI22xp5_ASAP7_75t_SL g158760 (.A1(\u4_mem[2] [19]),
    .A2(n_35632),
    .B1(\u4_mem[3] [19]),
    .B2(n_30078),
    .Y(n_1346));
 AOI22xp5_ASAP7_75t_SL g158768 (.A1(\u4_mem[1] [3]),
    .A2(n_50709),
    .B1(\u4_mem[3] [3]),
    .B2(n_30078),
    .Y(n_775));
 AOI22xp33_ASAP7_75t_SL g158771 (.A1(\u4_mem[2] [4]),
    .A2(n_35632),
    .B1(n_30078),
    .B2(\u4_mem[3] [4]),
    .Y(n_1145));
 AOI22xp5_ASAP7_75t_SL g158775 (.A1(n_35632),
    .A2(\u4_mem[2] [6]),
    .B1(\u4_mem[3] [6]),
    .B2(n_30078),
    .Y(n_769));
 AOI22xp5_ASAP7_75t_SL g158782 (.A1(\u4_mem[1] [14]),
    .A2(n_50709),
    .B1(\u4_mem[3] [14]),
    .B2(n_30078),
    .Y(n_1175));
 AOI22xp5_ASAP7_75t_SL g158784 (.A1(n_35632),
    .A2(\u4_mem[2] [7]),
    .B1(\u4_mem[3] [7]),
    .B2(n_30078),
    .Y(n_761));
 AOI22xp5_ASAP7_75t_SL g158786 (.A1(\u4_mem[1] [0]),
    .A2(n_50709),
    .B1(\u4_mem[3] [0]),
    .B2(n_30078),
    .Y(n_759));
 AOI22xp33_ASAP7_75t_SL g158789 (.A1(\u3_mem[1] [4]),
    .A2(n_43317),
    .B1(\u3_mem[3] [4]),
    .B2(n_71972),
    .Y(n_1244));
 AOI22xp5_ASAP7_75t_SL g158792 (.A1(\u4_mem[1] [10]),
    .A2(n_50709),
    .B1(\u4_mem[3] [10]),
    .B2(n_30078),
    .Y(n_1177));
 AOI22xp33_ASAP7_75t_SL g158795 (.A1(\u3_mem[1] [18]),
    .A2(n_43317),
    .B1(\u3_mem[3] [18]),
    .B2(n_71972),
    .Y(n_1863));
 AOI22xp5_ASAP7_75t_SL g158796 (.A1(n_43317),
    .A2(\u3_mem[1] [7]),
    .B1(\u3_mem[3] [7]),
    .B2(n_71972),
    .Y(n_1241));
 AOI22xp5_ASAP7_75t_SL g158803 (.A1(\u4_mem[2] [8]),
    .A2(n_35632),
    .B1(\u4_mem[3] [8]),
    .B2(n_30078),
    .Y(n_752));
 AOI22xp5_ASAP7_75t_SL g158819 (.A1(\u4_mem[1] [1]),
    .A2(n_50709),
    .B1(\u4_mem[3] [1]),
    .B2(n_30078),
    .Y(n_742));
 OAI22xp5_ASAP7_75t_SL g158829 (.A1(n_14313),
    .A2(n_10937),
    .B1(n_1680),
    .B2(n_1679),
    .Y(n_4883));
 OAI22xp5_ASAP7_75t_SL g158831 (.A1(n_14301),
    .A2(n_48648),
    .B1(n_1677),
    .B2(n_50458),
    .Y(n_5211));
 INVxp33_ASAP7_75t_R g158832 (.A(n_713),
    .Y(n_714));
 INVxp33_ASAP7_75t_R g158833 (.A(n_736),
    .Y(n_737));
 INVxp67_ASAP7_75t_L g158834 (.A(n_696),
    .Y(n_1289));
 INVxp33_ASAP7_75t_R g158836 (.A(u1_sr[0]),
    .Y(n_1231));
 INVxp33_ASAP7_75t_R g158842 (.A(n_7084),
    .Y(n_1186));
 NOR2xp33_ASAP7_75t_R g158846 (.A(n_40417),
    .B(n_640),
    .Y(n_1229));
 AND2x2_ASAP7_75t_R g158847 (.A(n_19010),
    .B(n_47541),
    .Y(n_720));
 NOR2xp33_ASAP7_75t_R g158848 (.A(n_19010),
    .B(n_47541),
    .Y(n_719));
 NAND2xp5_ASAP7_75t_L g158849 (.A(u10_din_tmp1[10]),
    .B(n_24336),
    .Y(n_1228));
 NOR2xp33_ASAP7_75t_R g158854 (.A(u2_to_cnt[2]),
    .B(n_705),
    .Y(n_706));
 NAND2xp5_ASAP7_75t_SL g158862 (.A(u10_din_tmp1[7]),
    .B(n_24336),
    .Y(n_1358));
 NAND2xp5_ASAP7_75t_SL g158877 (.A(u10_din_tmp1[14]),
    .B(n_24336),
    .Y(n_1214));
 NAND2xp5_ASAP7_75t_SL g158878 (.A(n_24336),
    .B(u10_din_tmp1[12]),
    .Y(n_1209));
 NAND2xp5_ASAP7_75t_SL g158879 (.A(u10_din_tmp1[15]),
    .B(n_24336),
    .Y(n_1208));
 NAND2xp5_ASAP7_75t_L g158886 (.A(\u7_mem[0] [4]),
    .B(n_49129),
    .Y(n_672));
 NAND2xp5_ASAP7_75t_SL g158890 (.A(u10_din_tmp1[13]),
    .B(n_24336),
    .Y(n_1201));
 NAND2xp33_ASAP7_75t_R g158894 (.A(n_633),
    .B(u2_cnt[0]),
    .Y(n_713));
 NAND2xp33_ASAP7_75t_R g158895 (.A(n_655),
    .B(n_1088),
    .Y(n_736));
 NAND2xp5_ASAP7_75t_SL g158901 (.A(n_71972),
    .B(u3_rp[0]),
    .Y(n_616));
 NOR2xp67_ASAP7_75t_SL g158902 (.A(n_183),
    .B(n_347),
    .Y(n_696));
 NOR2x1_ASAP7_75t_L g158905 (.A(n_21878),
    .B(n_1365),
    .Y(n_4665));
 NOR2x1_ASAP7_75t_L g158906 (.A(n_1680),
    .B(n_10937),
    .Y(n_4919));
 NOR2x1_ASAP7_75t_L g158907 (.A(n_21646),
    .B(n_10937),
    .Y(n_4907));
 NOR2xp67_ASAP7_75t_SL g158908 (.A(n_26807),
    .B(n_1534),
    .Y(n_4695));
 NOR2x1_ASAP7_75t_R g158909 (.A(n_1704),
    .B(n_10937),
    .Y(n_4911));
 NOR2xp67_ASAP7_75t_L g158910 (.A(n_36288),
    .B(n_10937),
    .Y(n_4905));
 NOR2x1_ASAP7_75t_L g158911 (.A(n_1681),
    .B(n_10937),
    .Y(n_4915));
 NOR2x1_ASAP7_75t_R g158912 (.A(n_21631),
    .B(n_10937),
    .Y(n_4901));
 NOR2xp67_ASAP7_75t_SL g158913 (.A(n_21709),
    .B(n_10937),
    .Y(n_4899));
 NOR2xp67_ASAP7_75t_SL g158915 (.A(n_34500),
    .B(n_48637),
    .Y(n_5177));
 NOR2xp67_ASAP7_75t_SL g158916 (.A(n_26819),
    .B(n_1534),
    .Y(n_4667));
 NOR2x1_ASAP7_75t_L g158918 (.A(n_26823),
    .B(n_1365),
    .Y(n_4671));
 NOR2x1_ASAP7_75t_L g158922 (.A(n_26827),
    .B(n_1365),
    .Y(n_4675));
 NOR2xp67_ASAP7_75t_SL g158924 (.A(n_11693),
    .B(n_1365),
    .Y(n_4691));
 NOR2x1_ASAP7_75t_R g158926 (.A(n_34492),
    .B(n_48648),
    .Y(n_5173));
 NOR2x1_ASAP7_75t_L g158927 (.A(n_14309),
    .B(n_10937),
    .Y(n_4909));
 NOR2x1_ASAP7_75t_L g158929 (.A(n_21697),
    .B(n_10937),
    .Y(n_4917));
 NAND2xp33_ASAP7_75t_R g158930 (.A(u2_cnt[2]),
    .B(n_655),
    .Y(n_2290));
 NOR2xp67_ASAP7_75t_SL g158931 (.A(n_24886),
    .B(n_48637),
    .Y(n_5181));
 NOR2x1_ASAP7_75t_R g158932 (.A(n_21638),
    .B(n_10937),
    .Y(n_4903));
 NOR2x1_ASAP7_75t_L g158933 (.A(n_21705),
    .B(n_10937),
    .Y(n_4913));
 NOR2xp67_ASAP7_75t_SL g158934 (.A(n_26815),
    .B(n_1534),
    .Y(n_4673));
 NOR2xp67_ASAP7_75t_SL g158935 (.A(n_1699),
    .B(n_1365),
    .Y(n_4689));
 NOR2xp67_ASAP7_75t_SL g158936 (.A(n_48052),
    .B(n_48637),
    .Y(n_5171));
 NOR2x1_ASAP7_75t_SL g158937 (.A(n_26811),
    .B(n_1534),
    .Y(n_4693));
 NOR2xp67_ASAP7_75t_SL g158938 (.A(n_1714),
    .B(n_48637),
    .Y(n_5185));
 NOR2xp67_ASAP7_75t_SL g158939 (.A(n_14288),
    .B(n_1365),
    .Y(n_4661));
 NOR2xp67_ASAP7_75t_SL g158940 (.A(n_21669),
    .B(n_1365),
    .Y(n_4663));
 INVxp67_ASAP7_75t_SL g158944 (.A(n_28955),
    .Y(n_707));
 INVxp67_ASAP7_75t_SL g158946 (.A(n_24738),
    .Y(n_703));
 INVxp33_ASAP7_75t_R g158947 (.A(n_26254),
    .Y(n_670));
 INVx1_ASAP7_75t_L g158948 (.A(n_18886),
    .Y(n_603));
 INVx1_ASAP7_75t_SL g158960 (.A(n_29364),
    .Y(n_1372));
 INVxp33_ASAP7_75t_R g158963 (.A(n_7196),
    .Y(n_700));
 INVx3_ASAP7_75t_SL g158969 (.A(n_36011),
    .Y(n_1766));
 NAND4xp25_ASAP7_75t_SL g158982 (.A(n_162),
    .B(n_1919),
    .C(u2_res_cnt[0]),
    .D(u2_res_cnt[2]),
    .Y(n_607));
 NAND2xp33_ASAP7_75t_R g158984 (.A(n_634),
    .B(n_633),
    .Y(n_635));
 AOI22xp5_ASAP7_75t_R g158985 (.A1(u13_intm_r[20]),
    .A2(u13_ints_r[20]),
    .B1(u13_intm_r[17]),
    .B2(u13_ints_r[17]),
    .Y(n_468));
 AOI22xp5_ASAP7_75t_SL g158986 (.A1(u13_intm_r[22]),
    .A2(u13_ints_r[22]),
    .B1(u13_intm_r[19]),
    .B2(u13_ints_r[19]),
    .Y(n_490));
 AOI22xp5_ASAP7_75t_SL g158988 (.A1(u13_intm_r[2]),
    .A2(u13_ints_r[2]),
    .B1(u13_intm_r[1]),
    .B2(u13_ints_r[1]),
    .Y(n_442));
 AOI22xp33_ASAP7_75t_SL g158989 (.A1(u13_intm_r[11]),
    .A2(u13_ints_r[11]),
    .B1(u13_intm_r[10]),
    .B2(u13_ints_r[10]),
    .Y(n_467));
 AOI22xp33_ASAP7_75t_SL g158990 (.A1(u13_intm_r[12]),
    .A2(u13_ints_r[12]),
    .B1(u13_intm_r[9]),
    .B2(u13_ints_r[9]),
    .Y(n_462));
 AOI22xp33_ASAP7_75t_SL g158991 (.A1(u13_intm_r[13]),
    .A2(u13_ints_r[13]),
    .B1(u13_intm_r[8]),
    .B2(u13_ints_r[8]),
    .Y(n_445));
 AOI22xp33_ASAP7_75t_SL g158992 (.A1(in_slt6[17]),
    .A2(n_728),
    .B1(in_slt6[19]),
    .B2(n_1361),
    .Y(n_729));
 AOI22xp33_ASAP7_75t_SL g158994 (.A1(u13_intm_r[23]),
    .A2(u13_ints_r[23]),
    .B1(u13_intm_r[18]),
    .B2(u13_ints_r[18]),
    .Y(n_454));
 AOI22xp5_ASAP7_75t_SL g158995 (.A1(u13_intm_r[27]),
    .A2(u13_ints_r[27]),
    .B1(u13_intm_r[26]),
    .B2(u13_ints_r[26]),
    .Y(n_443));
 AOI22xp33_ASAP7_75t_SL g158996 (.A1(u13_intm_r[25]),
    .A2(u13_ints_r[25]),
    .B1(u13_intm_r[24]),
    .B2(u13_ints_r[24]),
    .Y(n_461));
 AOI22xp5_ASAP7_75t_SL g158997 (.A1(in_slt4[16]),
    .A2(n_1667),
    .B1(in_slt4[18]),
    .B2(n_1666),
    .Y(n_1527));
 AOI22xp5_ASAP7_75t_SL g158998 (.A1(in_slt4[17]),
    .A2(n_1667),
    .B1(in_slt4[19]),
    .B2(n_1666),
    .Y(n_1528));
 AOI22xp5_ASAP7_75t_SL g159 (.A1(\u6_mem[3] [9]),
    .A2(n_41152),
    .B1(\u6_mem[2] [9]),
    .B2(n_77853),
    .Y(n_12106));
 AOI22xp33_ASAP7_75t_SL g159000 (.A1(in_slt6[16]),
    .A2(n_728),
    .B1(in_slt6[18]),
    .B2(n_1361),
    .Y(n_744));
 AOI22xp5_ASAP7_75t_SL g159001 (.A1(u13_intm_r[16]),
    .A2(u13_ints_r[16]),
    .B1(u13_intm_r[4]),
    .B2(u13_ints_r[4]),
    .Y(n_451));
 AOI22xp33_ASAP7_75t_SL g159002 (.A1(u13_intm_r[7]),
    .A2(u13_ints_r[7]),
    .B1(u13_intm_r[6]),
    .B2(u13_ints_r[6]),
    .Y(n_363));
 AOI22xp33_ASAP7_75t_SL g159003 (.A1(u13_intm_r[5]),
    .A2(u13_ints_r[5]),
    .B1(u13_intm_r[3]),
    .B2(u13_ints_r[3]),
    .Y(n_452));
 AOI21xp33_ASAP7_75t_R g159011 (.A1(u15_rdd3),
    .A2(crac_rd_done),
    .B(n_39),
    .Y(n_460));
 NOR2xp33_ASAP7_75t_R g159022 (.A(n_634),
    .B(n_633),
    .Y(n_1082));
 OAI22xp5_ASAP7_75t_SL g159025 (.A1(u11_wp[3]),
    .A2(n_506),
    .B1(u11_rp[2]),
    .B2(n_105),
    .Y(n_1058));
 AND2x2_ASAP7_75t_R g159034 (.A(n_634),
    .B(n_528),
    .Y(n_1336));
 NAND2xp5_ASAP7_75t_SL g159055 (.A(n_695),
    .B(n_71972),
    .Y(n_1782));
 AND2x4_ASAP7_75t_SL g159059_dup212431 (.A(n_53365),
    .B(n_49129),
    .Y(n_65055));
 AND2x4_ASAP7_75t_SL g159064 (.A(n_65643),
    .B(n_7668),
    .Y(n_1459));
 OR2x2_ASAP7_75t_SL g159065 (.A(n_640),
    .B(n_7564),
    .Y(n_1783));
 NAND2x1_ASAP7_75t_SL g159070 (.A(n_36008),
    .B(n_50709),
    .Y(n_1762));
 AND2x2_ASAP7_75t_SL g159071 (.A(n_36008),
    .B(n_50709),
    .Y(n_1765));
 AND2x2_ASAP7_75t_SL g159072 (.A(n_31888),
    .B(n_7668),
    .Y(n_2002));
 OR2x2_ASAP7_75t_SL g159073 (.A(n_640),
    .B(n_7567),
    .Y(n_1285));
 INVxp33_ASAP7_75t_R g159082 (.A(u1_sdata_in_r),
    .Y(n_560));
 HB1xp67_ASAP7_75t_SL g159085 (.A(n_347),
    .Y(n_705));
 INVxp33_ASAP7_75t_R g159086 (.A(u2_bit_clk_r),
    .Y(n_806));
 INVx1_ASAP7_75t_SL g159088 (.A(n_70325),
    .Y(n_624));
 NAND2xp33_ASAP7_75t_R g159145 (.A(u10_wp[3]),
    .B(n_557),
    .Y(n_1029));
 NAND2xp5_ASAP7_75t_SL g159146 (.A(n_28954),
    .B(n_225),
    .Y(n_625));
 NAND2xp33_ASAP7_75t_R g159147 (.A(u9_wp[3]),
    .B(n_521),
    .Y(n_786));
 NAND2xp5_ASAP7_75t_L g159149 (.A(in_slt1[11]),
    .B(oc0_cfg[1]),
    .Y(n_269));
 NOR2xp33_ASAP7_75t_SL g159152 (.A(u26_ps_cnt[3]),
    .B(u26_ps_cnt[2]),
    .Y(n_278));
 NOR2xp33_ASAP7_75t_R g159153 (.A(u14_u4_full_empty_r),
    .B(n_4075),
    .Y(n_491));
 NOR2xp33_ASAP7_75t_R g159154 (.A(u14_u0_full_empty_r),
    .B(n_4075),
    .Y(n_390));
 OR2x2_ASAP7_75t_L g159156 (.A(u14_u3_full_empty_r),
    .B(n_4075),
    .Y(n_389));
 OR2x2_ASAP7_75t_L g159157 (.A(u14_u1_full_empty_r),
    .B(n_4075),
    .Y(n_388));
 NOR2xp33_ASAP7_75t_R g159158 (.A(u14_u5_full_empty_r),
    .B(n_4075),
    .Y(n_387));
 NOR2xp33_ASAP7_75t_R g159159 (.A(dma_ack_i[7]),
    .B(n_15),
    .Y(n_487));
 NOR2xp33_ASAP7_75t_R g159161 (.A(dma_ack_i[8]),
    .B(n_108),
    .Y(n_391));
 NOR2x1_ASAP7_75t_SL g159173 (.A(u14_u1_en_out_l2),
    .B(n_256),
    .Y(n_519));
 NAND2xp5_ASAP7_75t_SL g159177 (.A(u2_to_cnt[0]),
    .B(u2_to_cnt[1]),
    .Y(n_347));
 NOR2xp33_ASAP7_75t_R g159178 (.A(n_147),
    .B(n_634),
    .Y(n_1088));
 NOR2xp33_ASAP7_75t_R g159181 (.A(n_148),
    .B(n_2288),
    .Y(n_655));
 NAND2x1_ASAP7_75t_SL g159183 (.A(out_slt0[8]),
    .B(n_31579),
    .Y(n_3468));
 NAND2xp33_ASAP7_75t_R g159185_dup163779 (.A(wb_addr_i[5]),
    .B(n_6552),
    .Y(n_7231));
 NOR2xp33_ASAP7_75t_R g159186 (.A(u2_cnt[2]),
    .B(u2_cnt[1]),
    .Y(n_633));
 INVx1_ASAP7_75t_L g159223 (.A(n_522),
    .Y(n_523));
 INVxp33_ASAP7_75t_R g159233 (.A(n_1645),
    .Y(n_588));
 INVx1_ASAP7_75t_L g159239 (.A(n_7668),
    .Y(n_589));
 INVxp67_ASAP7_75t_R g159242 (.A(n_695),
    .Y(n_2523));
 INVx2_ASAP7_75t_SL g159247 (.A(n_640),
    .Y(n_695));
 INVxp67_ASAP7_75t_SL g159266 (.A(n_71972),
    .Y(n_450));
 BUFx4f_ASAP7_75t_SL g159280_dup168589 (.A(n_20426),
    .Y(n_13236));
 INVx4_ASAP7_75t_SL g159288 (.A(n_24336),
    .Y(n_1365));
 INVx4_ASAP7_75t_SL g159291 (.A(n_24336),
    .Y(n_1534));
 NAND2xp5_ASAP7_75t_R g159293 (.A(u5_wp[2]),
    .B(n_455),
    .Y(n_456));
 NOR2xp33_ASAP7_75t_R g159295 (.A(crac_wr),
    .B(u15_crac_rd),
    .Y(n_280));
 NAND2x1_ASAP7_75t_L g159297 (.A(n_24737),
    .B(n_203),
    .Y(n_4276));
 NOR2xp33_ASAP7_75t_SL g159301 (.A(oc4_cfg[2]),
    .B(n_70326),
    .Y(n_370));
 NAND2xp33_ASAP7_75t_L g159302 (.A(oc3_cfg[0]),
    .B(n_155),
    .Y(n_459));
 NAND2xp33_ASAP7_75t_R g159303 (.A(u11_wp[3]),
    .B(n_659),
    .Y(n_660));
 NAND2xp5_ASAP7_75t_SL g159304 (.A(u3_wp[2]),
    .B(n_2687),
    .Y(n_469));
 NAND2xp5_ASAP7_75t_SL g159305 (.A(u8_wp[2]),
    .B(n_2689),
    .Y(n_463));
 NAND2xp5_ASAP7_75t_SL g159306 (.A(u6_wp[2]),
    .B(n_2693),
    .Y(n_369));
 NAND2xp5_ASAP7_75t_SL g159307 (.A(n_24737),
    .B(n_259),
    .Y(n_522));
 NAND2xp5_ASAP7_75t_L g159308 (.A(u7_wp[2]),
    .B(n_2691),
    .Y(n_464));
 NAND2xp5_ASAP7_75t_SL g159309 (.A(u4_wp[2]),
    .B(n_65325),
    .Y(n_368));
 NAND2xp5_ASAP7_75t_SL g159311 (.A(n_19616),
    .B(u5_rp[0]),
    .Y(n_273));
 NAND2xp33_ASAP7_75t_SL g159313 (.A(n_64714),
    .B(u7_rp[0]),
    .Y(n_267));
 NOR2xp33_ASAP7_75t_R g159319 (.A(u2_cnt[7]),
    .B(u2_cnt[4]),
    .Y(n_528));
 NOR2xp33_ASAP7_75t_R g159320 (.A(u2_cnt[1]),
    .B(n_2288),
    .Y(n_1193));
 NOR2xp33_ASAP7_75t_R g159327 (.A(n_1192),
    .B(n_1903),
    .Y(n_1645));
 OR2x2_ASAP7_75t_SL g159332 (.A(n_417),
    .B(oc0_cfg[3]),
    .Y(n_640));
 AND2x2_ASAP7_75t_SL g159333 (.A(u8_rp[0]),
    .B(n_253),
    .Y(n_636));
 OR2x2_ASAP7_75t_SL g159343 (.A(u4_rp[1]),
    .B(u4_rp[2]),
    .Y(n_415));
 AND2x4_ASAP7_75t_SL g159365 (.A(u11_rp[0]),
    .B(n_13764),
    .Y(n_1167));
 AND2x4_ASAP7_75t_SL g159366 (.A(u9_rp[0]),
    .B(n_13758),
    .Y(n_1171));
 NOR2x1_ASAP7_75t_SL g159374 (.A(n_336),
    .B(n_275),
    .Y(n_684));
 INVxp67_ASAP7_75t_R g159376 (.A(crac_din[8]),
    .Y(n_99));
 INVxp33_ASAP7_75t_R g159378 (.A(\u7_mem[2] [23]),
    .Y(n_93));
 INVxp33_ASAP7_75t_R g159379 (.A(u15_rdd2),
    .Y(n_39));
 INVxp33_ASAP7_75t_R g159381 (.A(crac_din[11]),
    .Y(n_130));
 INVxp67_ASAP7_75t_L g159383 (.A(crac_din[6]),
    .Y(n_49));
 INVxp33_ASAP7_75t_R g159384 (.A(crac_din[3]),
    .Y(n_42));
 INVx1_ASAP7_75t_L g159385 (.A(crac_din[4]),
    .Y(n_158));
 INVxp33_ASAP7_75t_R g159386 (.A(\u4_mem[3] [28]),
    .Y(n_156));
 INVxp67_ASAP7_75t_L g159387 (.A(u13_occ1_r[7]),
    .Y(n_133));
 INVx1_ASAP7_75t_SL g159389 (.A(u13_occ0_r[7]),
    .Y(n_41));
 INVx1_ASAP7_75t_SL g159390 (.A(u13_occ0_r[15]),
    .Y(n_97));
 INVxp67_ASAP7_75t_SL g159392 (.A(crac_din[13]),
    .Y(n_47));
 INVxp67_ASAP7_75t_L g159393 (.A(u13_occ1_r[15]),
    .Y(n_81));
 INVxp67_ASAP7_75t_R g159394 (.A(\u5_mem[1] [29]),
    .Y(n_149));
 INVx1_ASAP7_75t_L g159396 (.A(crac_din[7]),
    .Y(n_153));
 INVxp33_ASAP7_75t_R g159398 (.A(\u5_mem[0] [20]),
    .Y(n_90));
 INVx1_ASAP7_75t_L g159399 (.A(u13_icc_r[7]),
    .Y(n_1496));
 INVx1_ASAP7_75t_SL g159401 (.A(crac_din[2]),
    .Y(n_95));
 INVxp67_ASAP7_75t_R g159402 (.A(u13_icc_r[23]),
    .Y(n_12));
 INVx1_ASAP7_75t_R g159403 (.A(crac_din[12]),
    .Y(n_76));
 INVxp33_ASAP7_75t_R g159406 (.A(\u4_mem[0] [28]),
    .Y(n_66));
 INVx1_ASAP7_75t_L g159407 (.A(u13_icc_r[15]),
    .Y(n_1494));
 INVxp67_ASAP7_75t_R g159409 (.A(\u4_mem[1] [25]),
    .Y(n_104));
 INVxp67_ASAP7_75t_L g159411 (.A(crac_din[1]),
    .Y(n_157));
 INVxp33_ASAP7_75t_R g159412 (.A(\u5_mem[1] [28]),
    .Y(n_3));
 INVxp67_ASAP7_75t_L g159413 (.A(crac_din[15]),
    .Y(n_152));
 INVxp67_ASAP7_75t_R g159414 (.A(crac_din[0]),
    .Y(n_65));
 INVxp33_ASAP7_75t_R g159421 (.A(u12_wb_ack_o_745),
    .Y(n_31561));
 INVxp33_ASAP7_75t_R g159423 (.A(\u4_mem[1] [28]),
    .Y(n_37));
 INVxp67_ASAP7_75t_L g159426 (.A(u14_u1_en_out_l2),
    .Y(n_43));
 INVxp67_ASAP7_75t_R g159427 (.A(\u7_mem[3] [23]),
    .Y(n_71));
 INVxp67_ASAP7_75t_R g159429 (.A(\u7_mem[3] [24]),
    .Y(n_67));
 INVxp67_ASAP7_75t_R g159431 (.A(\u7_mem[3] [26]),
    .Y(n_6));
 INVxp33_ASAP7_75t_R g159432 (.A(\u4_mem[1] [20]),
    .Y(n_58));
 INVxp33_ASAP7_75t_R g159433 (.A(\u4_mem[2] [20]),
    .Y(n_24));
 INVxp33_ASAP7_75t_R g159434 (.A(\u4_mem[3] [21]),
    .Y(n_160));
 INVxp33_ASAP7_75t_R g159435 (.A(\u7_mem[2] [21]),
    .Y(n_123));
 INVxp67_ASAP7_75t_R g159436 (.A(\u7_mem[3] [22]),
    .Y(n_74));
 INVxp33_ASAP7_75t_R g159438 (.A(\u4_mem[0] [21]),
    .Y(n_94));
 INVxp67_ASAP7_75t_SL g159441 (.A(oc5_cfg[5]),
    .Y(n_59));
 INVx1_ASAP7_75t_L g159442 (.A(oc3_cfg[6]),
    .Y(n_2517));
 INVx1_ASAP7_75t_L g159444 (.A(ic0_cfg[5]),
    .Y(n_1503));
 INVx1_ASAP7_75t_SL g159445 (.A(u2_res_cnt[3]),
    .Y(n_162));
 HB1xp67_ASAP7_75t_L g159447 (.A(u13_ints_r[18]),
    .Y(n_2048));
 INVxp33_ASAP7_75t_L g159449 (.A(ic2_cfg[4]),
    .Y(n_88));
 INVx1_ASAP7_75t_SL g159450 (.A(ic2_cfg[1]),
    .Y(n_2640));
 INVxp33_ASAP7_75t_L g159451 (.A(ic2_cfg[5]),
    .Y(n_143));
 INVxp67_ASAP7_75t_R g159453 (.A(crac_out[19]),
    .Y(n_1319));
 INVxp33_ASAP7_75t_R g159454 (.A(n_289),
    .Y(n_290));
 INVxp67_ASAP7_75t_SL g159455 (.A(u13_intm_r[11]),
    .Y(n_289));
 HB1xp67_ASAP7_75t_L g159457 (.A(u13_intm_r[19]),
    .Y(n_291));
 HB1xp67_ASAP7_75t_L g159458 (.A(u13_ints_r[9]),
    .Y(n_2031));
 INVx1_ASAP7_75t_SL g159459 (.A(oc5_cfg[6]),
    .Y(n_1381));
 INVxp67_ASAP7_75t_R g159463 (.A(oc3_cfg[5]),
    .Y(n_212));
 HB1xp67_ASAP7_75t_SL g159464 (.A(u13_ints_r[5]),
    .Y(n_2106));
 HB1xp67_ASAP7_75t_SL g159465 (.A(u13_ints_r[11]),
    .Y(n_2065));
 INVx1_ASAP7_75t_L g159466 (.A(ic1_cfg[5]),
    .Y(n_1379));
 INVxp67_ASAP7_75t_R g159467 (.A(n_218),
    .Y(n_219));
 INVxp67_ASAP7_75t_R g159468 (.A(u13_ints_r[26]),
    .Y(n_218));
 INVx1_ASAP7_75t_SL g159470 (.A(u14_u7_en_out_l2),
    .Y(n_220));
 INVx1_ASAP7_75t_SL g159472 (.A(u14_u8_en_out_l2),
    .Y(n_295));
 INVxp67_ASAP7_75t_L g159475 (.A(crac_out[18]),
    .Y(n_1325));
 HB1xp67_ASAP7_75t_SL g159476 (.A(u13_ints_r[1]),
    .Y(n_2063));
 INVxp67_ASAP7_75t_SL g159477 (.A(oc0_cfg[1]),
    .Y(n_72));
 INVxp33_ASAP7_75t_R g159478 (.A(n_257),
    .Y(n_356));
 INVx1_ASAP7_75t_L g159480 (.A(oc0_cfg[6]),
    .Y(n_257));
 HB1xp67_ASAP7_75t_R g159481 (.A(u13_intm_r[6]),
    .Y(n_310));
 HB1xp67_ASAP7_75t_R g159483 (.A(u13_intm_r[10]),
    .Y(n_211));
 HB1xp67_ASAP7_75t_R g159485 (.A(oc1_cfg[4]),
    .Y(n_139));
 INVxp67_ASAP7_75t_SL g159486 (.A(oc1_cfg[4]),
    .Y(n_57));
 HB1xp67_ASAP7_75t_SL g159487 (.A(u13_ints_r[8]),
    .Y(n_2095));
 HB1xp67_ASAP7_75t_SL g159488 (.A(u13_ints_r[24]),
    .Y(n_2024));
 HB1xp67_ASAP7_75t_R g159490 (.A(u26_ps_cnt[5]),
    .Y(n_303));
 HB1xp67_ASAP7_75t_R g159492 (.A(u13_ints_r[3]),
    .Y(n_2038));
 INVxp67_ASAP7_75t_SL g159495 (.A(ic1_cfg[4]),
    .Y(n_1501));
 INVxp33_ASAP7_75t_R g159496 (.A(u13_ints_r[25]),
    .Y(n_63));
 HB1xp67_ASAP7_75t_SL g159498 (.A(u13_ints_r[14]),
    .Y(n_2130));
 HB1xp67_ASAP7_75t_SL g159500 (.A(u13_intm_r[8]),
    .Y(n_301));
 INVx1_ASAP7_75t_SL g159501 (.A(crac_out[17]),
    .Y(n_1322));
 INVx1_ASAP7_75t_SL g159502 (.A(n_31227),
    .Y(n_306));
 INVxp33_ASAP7_75t_R g159504 (.A(u13_ints_r[21]),
    .Y(n_34));
 HB1xp67_ASAP7_75t_SL g159506 (.A(u13_intm_r[18]),
    .Y(n_223));
 HB1xp67_ASAP7_75t_SL g159507 (.A(u13_ints_r[4]),
    .Y(n_2036));
 HB1xp67_ASAP7_75t_L g159510 (.A(u13_ints_r[23]),
    .Y(n_2678));
 INVx1_ASAP7_75t_SL g159511 (.A(ic1_cfg[1]),
    .Y(n_2645));
 INVxp33_ASAP7_75t_R g159512 (.A(u13_ints_r[27]),
    .Y(n_14));
 INVxp33_ASAP7_75t_R g159514 (.A(u13_ints_r[22]),
    .Y(n_75));
 HB1xp67_ASAP7_75t_SL g159517 (.A(u13_intm_r[4]),
    .Y(n_307));
 INVxp67_ASAP7_75t_SL g159518 (.A(ic0_cfg[4]),
    .Y(n_1376));
 HB1xp67_ASAP7_75t_L g159519 (.A(u13_ints_r[6]),
    .Y(n_2034));
 INVxp67_ASAP7_75t_R g159521 (.A(n_262),
    .Y(n_357));
 INVx1_ASAP7_75t_SL g159522 (.A(oc1_cfg[1]),
    .Y(n_262));
 INVxp33_ASAP7_75t_R g159527 (.A(u13_ints_r[16]),
    .Y(n_68));
 INVxp33_ASAP7_75t_R g159528 (.A(n_293),
    .Y(n_294));
 INVxp67_ASAP7_75t_SL g159529 (.A(oc5_cfg[4]),
    .Y(n_293));
 HB1xp67_ASAP7_75t_L g159531 (.A(u13_ints_r[10]),
    .Y(n_2029));
 HB1xp67_ASAP7_75t_SL g159533 (.A(u13_intm_r[23]),
    .Y(n_312));
 INVxp33_ASAP7_75t_R g159534 (.A(n_14906),
    .Y(n_360));
 INVxp67_ASAP7_75t_R g159537 (.A(u13_ints_r[28]),
    .Y(n_40));
 HB1xp67_ASAP7_75t_R g159538 (.A(u13_intm_r[9]),
    .Y(n_206));
 INVxp33_ASAP7_75t_R g159540 (.A(n_316),
    .Y(n_317));
 INVxp67_ASAP7_75t_SL g159541 (.A(u13_intm_r[3]),
    .Y(n_316));
 HB1xp67_ASAP7_75t_SL g159543 (.A(u13_intm_r[24]),
    .Y(n_227));
 HB1xp67_ASAP7_75t_R g159544 (.A(u13_intm_r[13]),
    .Y(n_319));
 INVxp33_ASAP7_75t_SL g159547 (.A(u13_ints_r[20]),
    .Y(n_2));
 INVxp67_ASAP7_75t_SL g159548 (.A(oc4_cfg[5]),
    .Y(n_103));
 INVxp33_ASAP7_75t_L g159549 (.A(n_258),
    .Y(n_362));
 INVx1_ASAP7_75t_SL g159551 (.A(u2_to_cnt[5]),
    .Y(n_258));
 INVxp33_ASAP7_75t_R g159552 (.A(n_229),
    .Y(n_230));
 INVxp67_ASAP7_75t_SL g159553 (.A(oc4_cfg[4]),
    .Y(n_229));
 HB1xp67_ASAP7_75t_L g159554 (.A(u13_ints_r[2]),
    .Y(n_2079));
 HB1xp67_ASAP7_75t_SL g159560 (.A(u2_to_cnt[3]),
    .Y(n_178));
 INVx1_ASAP7_75t_R g159561 (.A(u10_wp[3]),
    .Y(n_132));
 INVxp67_ASAP7_75t_R g159562 (.A(u2_res_cnt[2]),
    .Y(n_1));
 INVx1_ASAP7_75t_R g159570 (.A(u2_res_cnt[0]),
    .Y(n_1920));
 HB1xp67_ASAP7_75t_SL g159571 (.A(u2_to_cnt[1]),
    .Y(n_146));
 INVx1_ASAP7_75t_SL g159572 (.A(u11_rp[2]),
    .Y(n_506));
 INVx2_ASAP7_75t_L g159574 (.A(u2_res_cnt[1]),
    .Y(n_1919));
 INVxp67_ASAP7_75t_R g159575 (.A(crac_wr),
    .Y(n_23));
 INVx1_ASAP7_75t_SL g159578 (.A(u26_ps_cnt[1]),
    .Y(n_171));
 INVxp67_ASAP7_75t_SL g159585 (.A(u2_to_cnt[4]),
    .Y(n_1647));
 INVx1_ASAP7_75t_R g159586 (.A(u11_wp[3]),
    .Y(n_105));
 INVxp67_ASAP7_75t_SL g159590 (.A(u2_to_cnt[2]),
    .Y(n_183));
 HB1xp67_ASAP7_75t_SL g159594 (.A(n_184),
    .Y(n_339));
 INVx1_ASAP7_75t_L g159595 (.A(u26_cnt[0]),
    .Y(n_184));
 INVx1_ASAP7_75t_SL g159596 (.A(u2_to_cnt[0]),
    .Y(n_5));
 INVxp67_ASAP7_75t_SL g159598 (.A(u2_to_cnt[0]),
    .Y(n_321));
 HB1xp67_ASAP7_75t_L g159601 (.A(out_slt0[8]),
    .Y(n_181));
 INVxp67_ASAP7_75t_R g159604 (.A(n_256),
    .Y(n_517));
 INVx1_ASAP7_75t_SL g159607 (.A(out_slt0[11]),
    .Y(n_256));
 INVxp67_ASAP7_75t_SL g159612 (.A(n_172),
    .Y(n_366));
 INVx1_ASAP7_75t_SL g159614 (.A(u11_wp[0]),
    .Y(n_172));
 INVxp33_ASAP7_75t_R g159616 (.A(u2_cnt[1]),
    .Y(n_148));
 INVxp67_ASAP7_75t_L g159618 (.A(n_401),
    .Y(n_402));
 HB1xp67_ASAP7_75t_SL g159619 (.A(n_73),
    .Y(n_401));
 INVx1_ASAP7_75t_SL g159620 (.A(u10_wp[0]),
    .Y(n_73));
 INVx1_ASAP7_75t_SL g159627 (.A(n_113),
    .Y(n_399));
 INVxp33_ASAP7_75t_R g159631 (.A(u2_cnt[2]),
    .Y(n_147));
 INVxp67_ASAP7_75t_SL g159635 (.A(u7_wp[2]),
    .Y(n_16));
 INVxp33_ASAP7_75t_R g159638 (.A(u2_cnt[0]),
    .Y(n_2288));
 INVx2_ASAP7_75t_SL g159640 (.A(n_432),
    .Y(n_477));
 INVx2_ASAP7_75t_L g159644 (.A(oc5_cfg[2]),
    .Y(n_432));
 INVx1_ASAP7_75t_SL g159645 (.A(u6_rp[3]),
    .Y(n_2693));
 INVxp67_ASAP7_75t_L g159651 (.A(oc3_cfg[2]),
    .Y(n_155));
 HB1xp67_ASAP7_75t_SL g159652 (.A(oc3_cfg[2]),
    .Y(n_4027));
 INVx2_ASAP7_75t_L g159655 (.A(u7_rp[3]),
    .Y(n_2691));
 INVx1_ASAP7_75t_SL g159659 (.A(u5_rp[3]),
    .Y(n_455));
 HB1xp67_ASAP7_75t_SL g159661 (.A(n_332),
    .Y(n_4028));
 INVxp67_ASAP7_75t_SL g159662 (.A(n_608),
    .Y(n_332));
 INVx1_ASAP7_75t_SL g159663 (.A(oc0_cfg[2]),
    .Y(n_608));
 INVx1_ASAP7_75t_L g159664 (.A(u3_rp[3]),
    .Y(n_2687));
 INVx1_ASAP7_75t_SL g159666 (.A(u8_rp[3]),
    .Y(n_2689));
 INVx1_ASAP7_75t_SL g159668 (.A(n_101),
    .Y(n_247));
 INVx1_ASAP7_75t_SL g159671 (.A(oc4_cfg[2]),
    .Y(n_101));
 INVx1_ASAP7_75t_R g159674 (.A(n_7766),
    .Y(n_396));
 INVx3_ASAP7_75t_SL g159682 (.A(u7_wp[0]),
    .Y(n_2663));
 INVx2_ASAP7_75t_SL g159683 (.A(u7_wp[0]),
    .Y(n_136));
 INVx2_ASAP7_75t_SL g159695 (.A(n_259),
    .Y(n_203));
 INVx2_ASAP7_75t_SL g159696 (.A(u9_wp[2]),
    .Y(n_259));
 INVxp33_ASAP7_75t_L g159700 (.A(n_340),
    .Y(n_532));
 HB1xp67_ASAP7_75t_SL g159702 (.A(u9_wp[2]),
    .Y(n_340));
 INVx1_ASAP7_75t_SL g159705 (.A(n_12275),
    .Y(n_488));
 INVx2_ASAP7_75t_SL g159713 (.A(u10_wp[2]),
    .Y(n_234));
 INVx1_ASAP7_75t_SL g159723 (.A(n_231),
    .Y(n_232));
 INVx2_ASAP7_75t_SL g159724 (.A(u5_wp[0]),
    .Y(n_231));
 INVxp67_ASAP7_75t_SL g159725 (.A(n_19617),
    .Y(n_374));
 INVx2_ASAP7_75t_L g159727 (.A(u5_wp[0]),
    .Y(n_169));
 INVx1_ASAP7_75t_L g159733 (.A(n_225),
    .Y(n_226));
 INVx1_ASAP7_75t_L g159737 (.A(u11_wp[2]),
    .Y(n_217));
 INVxp33_ASAP7_75t_R g159758 (.A(u2_cnt[7]),
    .Y(n_2119));
 INVx1_ASAP7_75t_SL g159761 (.A(n_26382),
    .Y(n_2669));
 INVxp67_ASAP7_75t_SL g159768 (.A(n_26382),
    .Y(n_379));
 INVxp67_ASAP7_75t_SL g159772 (.A(oc1_cfg[0]),
    .Y(n_201));
 BUFx2_ASAP7_75t_SL g159776 (.A(oc1_cfg[0]),
    .Y(n_195));
 INVxp33_ASAP7_75t_R g159787 (.A(u2_cnt[4]),
    .Y(n_1914));
 INVxp33_ASAP7_75t_R g159802 (.A(u2_cnt[3]),
    .Y(n_634));
 BUFx2_ASAP7_75t_SL g159813 (.A(u7_wp[1]),
    .Y(n_2664));
 INVxp67_ASAP7_75t_R g159825 (.A(n_48675),
    .Y(n_2454));
 INVxp67_ASAP7_75t_SL g159829 (.A(u3_wp[1]),
    .Y(n_190));
 INVx1_ASAP7_75t_SL g159835 (.A(n_331),
    .Y(n_2753));
 INVxp67_ASAP7_75t_SL g159836 (.A(n_70326),
    .Y(n_331));
 INVx1_ASAP7_75t_SL g159840 (.A(n_57965),
    .Y(n_198));
 INVxp67_ASAP7_75t_SL g159845 (.A(n_179),
    .Y(n_245));
 HB1xp67_ASAP7_75t_SL g159846 (.A(oc3_cfg[0]),
    .Y(n_179));
 INVxp33_ASAP7_75t_R g159847 (.A(u2_cnt[6]),
    .Y(n_1192));
 INVxp67_ASAP7_75t_R g159852 (.A(n_34540),
    .Y(n_552));
 INVx1_ASAP7_75t_R g159863 (.A(n_509),
    .Y(n_556));
 INVx2_ASAP7_75t_L g159864 (.A(n_47740),
    .Y(n_509));
 INVxp33_ASAP7_75t_R g159869 (.A(u2_cnt[5]),
    .Y(n_1903));
 INVx2_ASAP7_75t_SL g159871 (.A(n_4542),
    .Y(n_521));
 BUFx2_ASAP7_75t_SL g159873 (.A(n_8186),
    .Y(n_4542));
 HB1xp67_ASAP7_75t_R g159879 (.A(ic2_cfg[0]),
    .Y(n_2788));
 INVxp33_ASAP7_75t_L g159881 (.A(n_19),
    .Y(n_281));
 INVxp67_ASAP7_75t_L g159882 (.A(n_4390),
    .Y(n_659));
 HB1xp67_ASAP7_75t_SL g159884 (.A(n_19),
    .Y(n_4390));
 INVx1_ASAP7_75t_SL g159885 (.A(ic2_cfg[0]),
    .Y(n_19));
 INVx2_ASAP7_75t_SL g159887 (.A(n_17686),
    .Y(n_557));
 BUFx12f_ASAP7_75t_SL g159894 (.A(n_423),
    .Y(n_1705));
 INVx1_ASAP7_75t_L g159895 (.A(n_423),
    .Y(n_1361));
 INVxp67_ASAP7_75t_R g159896 (.A(n_423),
    .Y(n_1523));
 BUFx2_ASAP7_75t_SL g159897 (.A(n_166),
    .Y(n_423));
 INVxp67_ASAP7_75t_SL g159898 (.A(ic2_cfg[2]),
    .Y(n_166));
 HB1xp67_ASAP7_75t_SL g159903 (.A(n_264),
    .Y(n_329));
 INVx1_ASAP7_75t_L g159904 (.A(n_431),
    .Y(n_1692));
 HB1xp67_ASAP7_75t_SL g159906 (.A(n_264),
    .Y(n_431));
 INVxp67_ASAP7_75t_SL g159907 (.A(ic0_cfg[2]),
    .Y(n_264));
 INVxp67_ASAP7_75t_SL g159908 (.A(n_285),
    .Y(n_286));
 INVx1_ASAP7_75t_SL g159909 (.A(ic0_cfg[2]),
    .Y(n_285));
 INVx2_ASAP7_75t_L g159913 (.A(n_330),
    .Y(n_1666));
 BUFx3_ASAP7_75t_SL g159915 (.A(n_185),
    .Y(n_330));
 INVxp67_ASAP7_75t_SL g159916 (.A(ic1_cfg[2]),
    .Y(n_185));
 INVxp67_ASAP7_75t_SL g159917 (.A(n_274),
    .Y(n_275));
 INVx1_ASAP7_75t_SL g159918 (.A(ic1_cfg[2]),
    .Y(n_274));
 INVx3_ASAP7_75t_SL g159919 (.A(n_573),
    .Y(n_2524));
 INVx2_ASAP7_75t_SL g159934 (.A(oc0_cfg[3]),
    .Y(n_176));
 INVx1_ASAP7_75t_L g159957 (.A(n_2013),
    .Y(n_4362));
 BUFx2_ASAP7_75t_SL g159958 (.A(n_79193),
    .Y(n_2013));
 INVx1_ASAP7_75t_SL g159966 (.A(oc5_cfg[3]),
    .Y(n_253));
 INVx1_ASAP7_75t_SL g159974 (.A(n_2428),
    .Y(n_666));
 BUFx2_ASAP7_75t_SL g159976 (.A(n_52768),
    .Y(n_2428));
 INVx1_ASAP7_75t_SL g159985 (.A(n_2188),
    .Y(n_842));
 INVx1_ASAP7_75t_R g159993 (.A(n_644),
    .Y(n_725));
 BUFx2_ASAP7_75t_L g159996 (.A(n_512),
    .Y(n_644));
 INVx1_ASAP7_75t_SL g159997 (.A(n_7671),
    .Y(n_512));
 INVx1_ASAP7_75t_SL g159998 (.A(n_643),
    .Y(n_4318));
 INVx2_ASAP7_75t_SL g16 (.A(wb_addr_i[3]),
    .Y(n_8177));
 INVxp33_ASAP7_75t_R g160 (.A(wb_data_i[16]),
    .Y(n_65947));
 INVx2_ASAP7_75t_SL g160007 (.A(n_2596),
    .Y(n_643));
 INVx1_ASAP7_75t_SL g160018 (.A(n_186),
    .Y(n_336));
 INVx1_ASAP7_75t_SL g160019 (.A(ic1_cfg[3]),
    .Y(n_186));
 INVx1_ASAP7_75t_SL g160027 (.A(n_265),
    .Y(n_427));
 INVx1_ASAP7_75t_SL g160028 (.A(ic0_cfg[3]),
    .Y(n_265));
 INVx2_ASAP7_75t_SL g160033 (.A(n_4548),
    .Y(n_1932));
 INVxp67_ASAP7_75t_L g160045 (.A(n_435),
    .Y(n_1362));
 HB1xp67_ASAP7_75t_SL g160046 (.A(n_263),
    .Y(n_435));
 INVx2_ASAP7_75t_SL g160049 (.A(n_1679),
    .Y(n_728));
 INVxp67_ASAP7_75t_SL g160051 (.A(ic2_cfg[3]),
    .Y(n_263));
 INVxp33_ASAP7_75t_R g160060 (.A(wb_data_i[0]),
    .Y(n_128));
 INVxp33_ASAP7_75t_R g160061 (.A(wb_data_i[29]),
    .Y(n_44));
 INVxp33_ASAP7_75t_R g160062 (.A(wb_data_i[30]),
    .Y(n_140));
 INVxp33_ASAP7_75t_R g160063 (.A(wb_data_i[1]),
    .Y(n_64));
 INVxp33_ASAP7_75t_R g160064 (.A(sdata_pad_i),
    .Y(n_107));
 INVxp33_ASAP7_75t_R g160065 (.A(\u4_mem[0] [25]),
    .Y(n_106));
 INVxp33_ASAP7_75t_R g160066 (.A(\u5_mem[0] [29]),
    .Y(n_51));
 INVxp33_ASAP7_75t_R g160067 (.A(\u7_mem[2] [22]),
    .Y(n_55));
 INVxp33_ASAP7_75t_R g160068 (.A(\u4_mem[1] [21]),
    .Y(n_144));
 INVxp67_ASAP7_75t_R g160069 (.A(\u7_mem[3] [21]),
    .Y(n_161));
 INVxp33_ASAP7_75t_R g160072 (.A(\u3_mem[2] [20]),
    .Y(n_52));
 INVxp67_ASAP7_75t_R g160074 (.A(\u3_mem[1] [29]),
    .Y(n_53));
 INVxp67_ASAP7_75t_R g160075 (.A(\u5_mem[2] [21]),
    .Y(n_154));
 INVxp33_ASAP7_75t_R g160076 (.A(\u4_mem[2] [21]),
    .Y(n_62));
 INVxp33_ASAP7_75t_R g160077 (.A(\u5_mem[0] [21]),
    .Y(n_89));
 INVxp33_ASAP7_75t_R g160078 (.A(\u4_mem[2] [28]),
    .Y(n_111));
 INVxp67_ASAP7_75t_R g160079 (.A(\u5_mem[2] [20]),
    .Y(n_69));
 INVxp33_ASAP7_75t_R g160080 (.A(\u3_mem[1] [24]),
    .Y(n_22));
 INVxp67_ASAP7_75t_R g160081 (.A(\u7_mem[2] [26]),
    .Y(n_116));
 INVxp33_ASAP7_75t_R g160083 (.A(\u5_mem[0] [25]),
    .Y(n_70));
 INVxp67_ASAP7_75t_R g160084 (.A(\u7_mem[2] [24]),
    .Y(n_84));
 INVxp67_ASAP7_75t_R g160085 (.A(\u5_mem[0] [28]),
    .Y(n_9));
 INVxp33_ASAP7_75t_R g160086 (.A(\u4_mem[0] [20]),
    .Y(n_21));
 INVxp33_ASAP7_75t_R g160087 (.A(\u5_mem[2] [28]),
    .Y(n_56));
 INVxp33_ASAP7_75t_R g160088 (.A(\u3_mem[3] [31]),
    .Y(n_20));
 INVxp33_ASAP7_75t_R g160089 (.A(\u5_mem[1] [20]),
    .Y(n_134));
 INVxp33_ASAP7_75t_R g160090 (.A(\u3_mem[2] [31]),
    .Y(n_48));
 INVxp67_ASAP7_75t_R g160091 (.A(\u5_mem[1] [21]),
    .Y(n_7));
 INVxp33_ASAP7_75t_R g160092 (.A(\u3_mem[2] [21]),
    .Y(n_118));
 INVxp33_ASAP7_75t_R g160093 (.A(\u4_mem[3] [20]),
    .Y(n_137));
 INVxp33_ASAP7_75t_R g160095 (.A(\u3_mem[3] [20]),
    .Y(n_79));
 INVx2_ASAP7_75t_R g160097 (.A(wb_cyc_i),
    .Y(n_38));
 INVx2_ASAP7_75t_L g160098 (.A(wb_stb_i),
    .Y(n_0));
 INVxp33_ASAP7_75t_R g160099 (.A(\u5_mem[1] [25]),
    .Y(n_4));
 INVxp33_ASAP7_75t_R g160100 (.A(out_slt0[14]),
    .Y(n_112));
 INVx1_ASAP7_75t_R g160103 (.A(in_slt6[18]),
    .Y(n_1680));
 INVx1_ASAP7_75t_R g160110 (.A(in_slt6[16]),
    .Y(n_1681));
 INVx1_ASAP7_75t_L g160112 (.A(in_slt3[9]),
    .Y(n_1714));
 INVx1_ASAP7_75t_R g160131 (.A(in_slt3[11]),
    .Y(n_1820));
 INVx1_ASAP7_75t_R g160140 (.A(in_slt3[19]),
    .Y(n_1677));
 INVx1_ASAP7_75t_L g160142 (.A(in_slt4[19]),
    .Y(n_1699));
 INVx1_ASAP7_75t_R g160144 (.A(in_slt3[18]),
    .Y(n_1678));
 INVx1_ASAP7_75t_R g160145 (.A(in_slt6[4]),
    .Y(n_1707));
 INVx1_ASAP7_75t_R g160147 (.A(in_slt6[14]),
    .Y(n_1704));
 INVxp67_ASAP7_75t_L g160151 (.A(in_slt6[19]),
    .Y(n_1701));
 INVxp67_ASAP7_75t_R g160153 (.A(u8_rp[0]),
    .Y(n_497));
 INVx1_ASAP7_75t_SL g160155 (.A(u3_rp[0]),
    .Y(n_417));
 INVxp67_ASAP7_75t_R g160156 (.A(u6_rp[0]),
    .Y(n_678));
 INVxp67_ASAP7_75t_SL g160157 (.A(u7_rp[0]),
    .Y(n_419));
 INVx1_ASAP7_75t_L g160159 (.A(in_slt0[15]),
    .Y(n_4075));
 INVxp33_ASAP7_75t_R g160160 (.A(bit_clk_pad_i),
    .Y(n_434));
 INVxp33_ASAP7_75t_R g161 (.A(wb_data_i[17]),
    .Y(n_65950));
 NAND4xp25_ASAP7_75t_SL g162 (.A(n_2332),
    .B(n_2074),
    .C(n_1753),
    .D(n_1803),
    .Y(n_7588));
 XNOR2xp5_ASAP7_75t_SL g162472 (.A(n_18896),
    .B(n_18742),
    .Y(n_5845));
 XNOR2xp5_ASAP7_75t_SL g162473 (.A(n_50812),
    .B(n_58734),
    .Y(n_5846));
 XNOR2xp5_ASAP7_75t_SL g162474 (.A(n_24375),
    .B(n_48437),
    .Y(n_5847));
 XNOR2xp5_ASAP7_75t_SL g162475 (.A(n_19594),
    .B(n_14013),
    .Y(n_5848));
 XNOR2xp5_ASAP7_75t_R g162476 (.A(u4_rp[3]),
    .B(n_30078),
    .Y(n_5849));
 AOI22xp5_ASAP7_75t_SL g162672 (.A1(n_50341),
    .A2(\u3_mem[0] [16]),
    .B1(\u3_mem[1] [16]),
    .B2(n_43317),
    .Y(n_6044));
 AOI22xp5_ASAP7_75t_SL g162680 (.A1(n_50341),
    .A2(\u3_mem[0] [8]),
    .B1(\u3_mem[2] [8]),
    .B2(n_7562),
    .Y(n_6051));
 AOI22xp33_ASAP7_75t_SL g162693 (.A1(\u3_mem[0] [17]),
    .A2(n_43318),
    .B1(n_43317),
    .B2(\u3_mem[1] [17]),
    .Y(n_6065));
 AO22x1_ASAP7_75t_SL g162845 (.A1(n_65055),
    .A2(\u7_mem[0] [22]),
    .B1(\u7_mem[1] [22]),
    .B2(n_65056),
    .Y(n_6232));
 AOI22xp5_ASAP7_75t_SL g162904 (.A1(n_49129),
    .A2(\u7_mem[0] [12]),
    .B1(\u7_mem[1] [12]),
    .B2(n_49617),
    .Y(n_6295));
 AOI22xp5_ASAP7_75t_SL g162906 (.A1(n_49129),
    .A2(\u7_mem[0] [15]),
    .B1(n_49617),
    .B2(\u7_mem[1] [15]),
    .Y(n_6297));
 HB1xp67_ASAP7_75t_SL g162909 (.A(n_49617),
    .Y(n_6299));
 AOI22xp5_ASAP7_75t_SL g162910 (.A1(\u7_mem[0] [7]),
    .A2(n_49129),
    .B1(\u7_mem[1] [7]),
    .B2(n_49617),
    .Y(n_6301));
 AND2x2_ASAP7_75t_L g163 (.A(out_slt4[19]),
    .B(n_43087),
    .Y(n_7589));
 AOI22xp33_ASAP7_75t_SL g163172 (.A1(u13_icc_r[23]),
    .A2(n_6615),
    .B1(n_312),
    .B2(n_7083),
    .Y(n_6583));
 AOI22xp33_ASAP7_75t_SL g163204 (.A1(crac_out[20]),
    .A2(n_22851),
    .B1(ic2_cfg[4]),
    .B2(n_6615),
    .Y(n_6616));
 AOI22xp33_ASAP7_75t_L g163310 (.A1(crac_out[22]),
    .A2(n_10867),
    .B1(ic2_cfg[6]),
    .B2(n_6615),
    .Y(n_6721));
 AND2x4_ASAP7_75t_SL g163319 (.A(n_7084),
    .B(rf_we),
    .Y(n_6732));
 INVx3_ASAP7_75t_SL g163643 (.A(n_8321),
    .Y(n_7082));
 INVx2_ASAP7_75t_R g163644 (.A(n_8321),
    .Y(n_7083));
 INVxp67_ASAP7_75t_L g163646 (.A(n_32317),
    .Y(n_7086));
 NOR2xp33_ASAP7_75t_SL g163647 (.A(n_32317),
    .B(n_316),
    .Y(n_7087));
 OR2x6_ASAP7_75t_SL g163648_dup (.A(n_32318),
    .B(n_32317),
    .Y(n_32335));
 NOR2xp33_ASAP7_75t_SL g163649 (.A(n_32317),
    .B(n_289),
    .Y(n_7089));
 AOI22xp33_ASAP7_75t_SL g163689 (.A1(n_22851),
    .A2(crac_out[16]),
    .B1(n_8247),
    .B2(ic2_cfg[0]),
    .Y(n_7132));
 NOR2x1_ASAP7_75t_R g163703_dup (.A(wb_addr_i[4]),
    .B(wb_addr_i[2]),
    .Y(n_7195));
 AOI221xp5_ASAP7_75t_SL g163706 (.A1(i6_dout[11]),
    .A2(n_14933),
    .B1(i4_dout[11]),
    .B2(n_8174),
    .C(n_7089),
    .Y(n_7152));
 AOI22xp33_ASAP7_75t_L g163720 (.A1(i6_dout[23]),
    .A2(n_8338),
    .B1(u13_occ0_r[23]),
    .B2(n_6961),
    .Y(n_7167));
 NAND2xp5_ASAP7_75t_L g163721 (.A(n_8338),
    .B(i6_dout[25]),
    .Y(n_7168));
 NAND2xp5_ASAP7_75t_L g163722 (.A(n_8338),
    .B(i6_dout[27]),
    .Y(n_7169));
 INVx2_ASAP7_75t_L g163723 (.A(n_8338),
    .Y(n_7170));
 NAND2xp5_ASAP7_75t_L g163724 (.A(i6_dout[22]),
    .B(n_8338),
    .Y(n_7171));
 NAND2xp5_ASAP7_75t_L g163725 (.A(i6_dout[26]),
    .B(n_8338),
    .Y(n_7172));
 NAND2xp5_ASAP7_75t_L g163726 (.A(i6_dout[21]),
    .B(n_8338),
    .Y(n_7173));
 NAND2xp5_ASAP7_75t_L g163727 (.A(i6_dout[16]),
    .B(n_8338),
    .Y(n_7174));
 NAND2xp5_ASAP7_75t_L g163728 (.A(i6_dout[28]),
    .B(n_8338),
    .Y(n_7175));
 NAND2xp5_ASAP7_75t_L g163729 (.A(i6_dout[20]),
    .B(n_8338),
    .Y(n_7176));
 AND2x2_ASAP7_75t_SL g163746 (.A(n_7195),
    .B(n_8256),
    .Y(n_7196));
 AOI22xp5_ASAP7_75t_R g163752 (.A1(i6_dout[17]),
    .A2(n_8338),
    .B1(i3_dout[17]),
    .B2(n_8235),
    .Y(n_7202));
 AOI22xp5_ASAP7_75t_R g163754 (.A1(i6_dout[6]),
    .A2(n_8338),
    .B1(i3_dout[6]),
    .B2(n_8235),
    .Y(n_7204));
 AOI22xp5_ASAP7_75t_R g163756 (.A1(i6_dout[7]),
    .A2(n_14933),
    .B1(i3_dout[7]),
    .B2(n_8235),
    .Y(n_7206));
 AOI22xp5_ASAP7_75t_R g163757 (.A1(i6_dout[0]),
    .A2(n_14933),
    .B1(i3_dout[0]),
    .B2(n_8235),
    .Y(n_7207));
 AOI22xp5_ASAP7_75t_R g163758 (.A1(i6_dout[2]),
    .A2(n_14933),
    .B1(i3_dout[2]),
    .B2(n_8235),
    .Y(n_7208));
 AOI22xp5_ASAP7_75t_R g163759 (.A1(i6_dout[4]),
    .A2(n_14933),
    .B1(i3_dout[4]),
    .B2(n_8235),
    .Y(n_7209));
 AOI22xp5_ASAP7_75t_R g163762 (.A1(i6_dout[9]),
    .A2(n_14933),
    .B1(i3_dout[9]),
    .B2(n_8235),
    .Y(n_7212));
 AOI22xp5_ASAP7_75t_L g163764 (.A1(i6_dout[12]),
    .A2(n_14933),
    .B1(i3_dout[12]),
    .B2(n_8341),
    .Y(n_7215));
 AOI22xp5_ASAP7_75t_L g163765 (.A1(i6_dout[14]),
    .A2(n_14933),
    .B1(i3_dout[14]),
    .B2(n_8341),
    .Y(n_7216));
 NAND2xp5_ASAP7_75t_L g163767 (.A(n_8341),
    .B(i3_dout[31]),
    .Y(n_7218));
 AOI22xp33_ASAP7_75t_SL g163768 (.A1(n_8341),
    .A2(i3_dout[24]),
    .B1(n_8173),
    .B2(i4_dout[24]),
    .Y(n_7219));
 NAND2xp5_ASAP7_75t_SL g163770 (.A(n_8341),
    .B(n_42621),
    .Y(n_7221));
 NAND2xp5_ASAP7_75t_L g163771 (.A(i3_dout[23]),
    .B(n_8341),
    .Y(n_7222));
 AOI21xp5_ASAP7_75t_SL g163774 (.A1(n_8341),
    .A2(i3_dout[1]),
    .B(n_1896),
    .Y(n_7225));
 AOI221xp5_ASAP7_75t_SL g163775 (.A1(n_8341),
    .A2(i3_dout[30]),
    .B1(n_8175),
    .B2(i4_dout[30]),
    .C(n_2518),
    .Y(n_7226));
 AOI221xp5_ASAP7_75t_SL g163776 (.A1(n_8341),
    .A2(i3_dout[29]),
    .B1(n_8175),
    .B2(i4_dout[29]),
    .C(n_2516),
    .Y(n_7227));
 HB1xp67_ASAP7_75t_L g163815 (.A(n_78274),
    .Y(n_7335));
 HB1xp67_ASAP7_75t_SL g163886 (.A(n_50388),
    .Y(n_7408));
 AOI22xp5_ASAP7_75t_SL g163888 (.A1(n_50342),
    .A2(\u3_mem[2] [1]),
    .B1(\u3_mem[3] [1]),
    .B2(n_71972),
    .Y(n_7410));
 AOI22xp33_ASAP7_75t_SL g163890 (.A1(n_50342),
    .A2(\u3_mem[2] [17]),
    .B1(n_71972),
    .B2(\u3_mem[3] [17]),
    .Y(n_7411));
 AOI22xp5_ASAP7_75t_SL g163893 (.A1(\u3_mem[0] [18]),
    .A2(n_50341),
    .B1(\u3_mem[2] [18]),
    .B2(n_50342),
    .Y(n_7414));
 AOI22xp5_ASAP7_75t_SL g163896 (.A1(\u3_mem[0] [7]),
    .A2(n_43318),
    .B1(n_50342),
    .B2(\u3_mem[2] [7]),
    .Y(n_7417));
 AOI22xp33_ASAP7_75t_L g163897 (.A1(\u3_mem[0] [5]),
    .A2(n_43318),
    .B1(n_50388),
    .B2(\u3_mem[2] [5]),
    .Y(n_7418));
 AND2x2_ASAP7_75t_L g163907 (.A(out_slt4[7]),
    .B(n_43087),
    .Y(n_7502));
 OAI211xp5_ASAP7_75t_SL g163908 (.A1(n_59639),
    .A2(n_4316),
    .B(n_7510),
    .C(n_21027),
    .Y(n_7511));
 NOR2xp67_ASAP7_75t_SL g163909 (.A(n_1769),
    .B(n_59341),
    .Y(n_7510));
 NAND2xp5_ASAP7_75t_SL g163910 (.A(n_7859),
    .B(n_79206),
    .Y(n_7514));
 NOR2xp67_ASAP7_75t_SL g163916 (.A(n_1788),
    .B(n_7522),
    .Y(n_7523));
 AO22x1_ASAP7_75t_SL g163917 (.A1(n_65056),
    .A2(\u7_mem[1] [21]),
    .B1(\u7_mem[0] [21]),
    .B2(n_65055),
    .Y(n_7522));
 AND2x2_ASAP7_75t_R g163919 (.A(out_slt3[5]),
    .B(n_5024),
    .Y(n_7524));
 AOI211xp5_ASAP7_75t_SL g163920 (.A1(n_17492),
    .A2(n_25405),
    .B(n_4379),
    .C(n_7526),
    .Y(n_7527));
 AND2x2_ASAP7_75t_R g163921 (.A(out_slt3[7]),
    .B(n_5024),
    .Y(n_7526));
 AOI22xp5_ASAP7_75t_SL g163923 (.A1(\u8_mem[0] [15]),
    .A2(n_59474),
    .B1(\u8_mem[1] [15]),
    .B2(n_78274),
    .Y(n_7538));
 AOI22xp5_ASAP7_75t_SL g163929 (.A1(n_59474),
    .A2(\u8_mem[0] [17]),
    .B1(n_78274),
    .B2(\u8_mem[1] [17]),
    .Y(n_7541));
 AOI22xp33_ASAP7_75t_SL g163930 (.A1(\u8_mem[0] [2]),
    .A2(n_59474),
    .B1(n_78274),
    .B2(\u8_mem[1] [2]),
    .Y(n_7542));
 AOI22xp5_ASAP7_75t_SL g163931 (.A1(\u8_mem[0] [3]),
    .A2(n_59474),
    .B1(\u8_mem[1] [3]),
    .B2(n_78274),
    .Y(n_7543));
 AOI22xp5_ASAP7_75t_SL g163932 (.A1(\u8_mem[0] [18]),
    .A2(n_59474),
    .B1(\u8_mem[1] [18]),
    .B2(n_78274),
    .Y(n_7544));
 NOR2xp33_ASAP7_75t_R g163947 (.A(u3_rp[1]),
    .B(n_6249),
    .Y(n_7562));
 OR2x6_ASAP7_75t_SL g163948 (.A(n_6249),
    .B(u3_rp[1]),
    .Y(n_7564));
 AND2x2_ASAP7_75t_L g163987 (.A(out_slt4[13]),
    .B(n_43087),
    .Y(n_7725));
 AND2x2_ASAP7_75t_SL g163992 (.A(out_slt7[12]),
    .B(n_5062),
    .Y(n_7735));
 INVxp33_ASAP7_75t_R g164 (.A(wb_data_i[8]),
    .Y(n_65977));
 INVx1_ASAP7_75t_SL g164004 (.A(n_7753),
    .Y(n_7754));
 NAND2x1_ASAP7_75t_SL g164005 (.A(n_1017),
    .B(n_769),
    .Y(n_7753));
 NAND2xp5_ASAP7_75t_SL g164006 (.A(n_7753),
    .B(n_24350),
    .Y(n_7755));
 INVx1_ASAP7_75t_SL g164007 (.A(n_7753),
    .Y(n_7756));
 BUFx3_ASAP7_75t_SL g164013 (.A(n_4024),
    .Y(n_7766));
 OR2x2_ASAP7_75t_SL g164038 (.A(u5_rp[2]),
    .B(u5_rp[1]),
    .Y(n_7872));
 AOI22xp33_ASAP7_75t_SL g164047 (.A1(\u5_mem[0] [12]),
    .A2(n_65642),
    .B1(n_65643),
    .B2(\u5_mem[2] [12]),
    .Y(n_7881));
 AOI22xp5_ASAP7_75t_SL g164049 (.A1(\u5_mem[0] [18]),
    .A2(n_65642),
    .B1(\u5_mem[2] [18]),
    .B2(n_65643),
    .Y(n_7883));
 INVx3_ASAP7_75t_SL g164055 (.A(u8_rp[2]),
    .Y(n_7888));
 NAND2xp33_ASAP7_75t_SL g164088 (.A(n_425),
    .B(n_2168),
    .Y(n_7927));
 AOI22xp5_ASAP7_75t_SL g164094 (.A1(n_38365),
    .A2(n_7939),
    .B1(n_79104),
    .B2(n_7941),
    .Y(n_7942));
 OAI211xp5_ASAP7_75t_SL g164096 (.A1(n_65000),
    .A2(n_725),
    .B(n_4320),
    .C(n_66666),
    .Y(n_7939));
 NAND2x1_ASAP7_75t_SL g164102 (.A(n_1032),
    .B(n_761),
    .Y(n_7990));
 AOI211xp5_ASAP7_75t_SL g164104 (.A1(n_2598),
    .A2(n_79104),
    .B(n_66678),
    .C(n_38376),
    .Y(n_7997));
 AOI211xp5_ASAP7_75t_SL g164106 (.A1(n_79207),
    .A2(n_5091),
    .B(n_79199),
    .C(n_73312),
    .Y(n_7999));
 AOI211xp5_ASAP7_75t_SL g164111 (.A1(n_18711),
    .A2(n_25405),
    .B(n_4366),
    .C(n_8005),
    .Y(n_8006));
 AND2x2_ASAP7_75t_R g164112 (.A(out_slt3[11]),
    .B(n_4513),
    .Y(n_8005));
 AOI211xp5_ASAP7_75t_SL g164113 (.A1(n_47554),
    .A2(n_25405),
    .B(n_4373),
    .C(n_8007),
    .Y(n_8008));
 AND2x2_ASAP7_75t_R g164114 (.A(out_slt3[10]),
    .B(n_4513),
    .Y(n_8007));
 AND2x2_ASAP7_75t_SL g164212 (.A(n_933),
    .B(n_759),
    .Y(n_8111));
 NAND2xp5_ASAP7_75t_SL g164213 (.A(n_933),
    .B(n_759),
    .Y(n_8112));
 AOI211xp5_ASAP7_75t_SL g164218 (.A1(n_8117),
    .A2(n_25405),
    .B(n_4347),
    .C(n_8118),
    .Y(n_8119));
 NAND4xp25_ASAP7_75t_SL g164219 (.A(n_2224),
    .B(n_1777),
    .C(n_7927),
    .D(n_1744),
    .Y(n_8117));
 AND2x2_ASAP7_75t_R g164220 (.A(out_slt3[13]),
    .B(n_4513),
    .Y(n_8118));
 BUFx6f_ASAP7_75t_SL g164241 (.A(n_8301),
    .Y(n_8173));
 BUFx6f_ASAP7_75t_SL g164243 (.A(n_8301),
    .Y(n_8174));
 BUFx3_ASAP7_75t_SL g164244 (.A(n_8173),
    .Y(n_8175));
 BUFx3_ASAP7_75t_L g164246_dup (.A(n_75733),
    .Y(n_10924));
 AOI21xp5_ASAP7_75t_SL g164248 (.A1(n_14098),
    .A2(n_375),
    .B(n_8191),
    .Y(n_8192));
 AND3x1_ASAP7_75t_SL g164250 (.A(rf_we),
    .B(n_75733),
    .C(n_6615),
    .Y(n_8191));
 NOR2x1p5_ASAP7_75t_L g164251 (.A(wb_addr_i[4]),
    .B(n_8189),
    .Y(n_6615));
 BUFx3_ASAP7_75t_SL g164265 (.A(n_8308),
    .Y(n_8212));
 OR2x2_ASAP7_75t_SL g164270_dup176230 (.A(n_26255),
    .B(n_22267),
    .Y(n_22268));
 OR2x2_ASAP7_75t_SL g164270_dup_dup (.A(n_26255),
    .B(n_22267),
    .Y(n_22276));
 INVx2_ASAP7_75t_R g164274 (.A(wb_addr_i[4]),
    .Y(n_8228));
 INVx2_ASAP7_75t_SL g164277 (.A(n_8313),
    .Y(n_8232));
 AND2x4_ASAP7_75t_SL g164279 (.A(n_8234),
    .B(n_8232),
    .Y(n_8235));
 AND2x2_ASAP7_75t_SL g164280 (.A(wb_addr_i[5]),
    .B(n_6552),
    .Y(n_8234));
 OR2x2_ASAP7_75t_SL g164284_dup (.A(n_10563),
    .B(wb_addr_i[4]),
    .Y(n_10576));
 AOI22xp5_ASAP7_75t_L g164286 (.A1(n_10565),
    .A2(ic2_cfg[5]),
    .B1(n_10867),
    .B2(crac_out[21]),
    .Y(n_8246));
 NOR2x1_ASAP7_75t_SL g164288 (.A(wb_addr_i[4]),
    .B(n_8183),
    .Y(n_8247));
 INVx2_ASAP7_75t_SL g164289 (.A(wb_addr_i[3]),
    .Y(n_8256));
 INVx6_ASAP7_75t_SL g164296 (.A(wb_addr_i[4]),
    .Y(n_8262));
 NOR2xp67_ASAP7_75t_SL g164306 (.A(n_8278),
    .B(n_8279),
    .Y(n_8280));
 OAI21xp33_ASAP7_75t_SL g164307 (.A1(n_8340),
    .A2(n_65896),
    .B(n_2273),
    .Y(n_8278));
 OAI211xp5_ASAP7_75t_SL g164308 (.A1(n_10613),
    .A2(n_14),
    .B(n_24341),
    .C(n_7169),
    .Y(n_8279));
 INVx3_ASAP7_75t_SL g164316 (.A(n_8321),
    .Y(n_7084));
 NOR2x1p5_ASAP7_75t_SL g164319 (.A(n_8299),
    .B(n_8319),
    .Y(n_8301));
 NAND2x1p5_ASAP7_75t_SL g164320 (.A(wb_addr_i[2]),
    .B(wb_addr_i[4]),
    .Y(n_8299));
 AND2x4_ASAP7_75t_SL g164326 (.A(n_8247),
    .B(rf_we),
    .Y(n_8306));
 NOR3x2_ASAP7_75t_SL g164327 (.B(wb_addr_i[3]),
    .C(wb_addr_i[4]),
    .Y(n_8308),
    .A(n_8307));
 INVx3_ASAP7_75t_SL g164328 (.A(wb_addr_i[2]),
    .Y(n_8307));
 INVx4_ASAP7_75t_SL g164330 (.A(wb_addr_i[2]),
    .Y(n_8309));
 INVx4_ASAP7_75t_SL g164332 (.A(wb_addr_i[2]),
    .Y(n_8311));
 NAND3x2_ASAP7_75t_SL g164334 (.B(wb_addr_i[3]),
    .C(wb_addr_i[4]),
    .Y(n_8313),
    .A(n_8309));
 NOR2x1p5_ASAP7_75t_SL g164335 (.A(wb_addr_i[6]),
    .B(n_8314),
    .Y(n_8315));
 INVx2_ASAP7_75t_L g164336 (.A(wb_addr_i[5]),
    .Y(n_8314));
 NAND3x2_ASAP7_75t_SL g164337 (.B(wb_addr_i[5]),
    .C(wb_addr_i[3]),
    .Y(n_8319),
    .A(n_6552));
 NAND3x2_ASAP7_75t_SL g164339 (.B(wb_addr_i[4]),
    .C(wb_addr_i[2]),
    .Y(n_8321),
    .A(n_8320));
 INVx4_ASAP7_75t_L g164340 (.A(wb_addr_i[3]),
    .Y(n_8320));
 NOR2xp33_ASAP7_75t_SL g164347 (.A(n_8332),
    .B(n_2473),
    .Y(n_8333));
 OAI211xp5_ASAP7_75t_SL g164348 (.A1(n_10613),
    .A2(n_40),
    .B(n_7175),
    .C(n_24626),
    .Y(n_8332));
 NOR2x1_ASAP7_75t_SL g164350 (.A(wb_addr_i[5]),
    .B(n_6552),
    .Y(n_8334));
 AND3x4_ASAP7_75t_SL g164351 (.A(n_8337),
    .B(n_8256),
    .C(n_8238),
    .Y(n_8338));
 NOR2x1_ASAP7_75t_SL g164352 (.A(wb_addr_i[5]),
    .B(n_6552),
    .Y(n_8337));
 OAI211xp5_ASAP7_75t_SL g165 (.A1(n_64103),
    .A2(n_6144),
    .B(n_4098),
    .C(n_57733),
    .Y(n_16899));
 OR2x4_ASAP7_75t_SL g165153 (.A(n_11124),
    .B(n_24367),
    .Y(n_9476));
 NAND4xp75_ASAP7_75t_SL g165213 (.A(rf_we),
    .B(n_8256),
    .C(n_8262),
    .D(wb_addr_i[2]),
    .Y(n_9555));
 AOI22xp33_ASAP7_75t_SL g165288 (.A1(n_1167),
    .A2(\u11_mem[1] [26]),
    .B1(n_46233),
    .B2(\u11_mem[3] [26]),
    .Y(n_9650));
 AOI22xp33_ASAP7_75t_SL g165292 (.A1(n_1167),
    .A2(\u11_mem[1] [16]),
    .B1(n_46233),
    .B2(\u11_mem[3] [16]),
    .Y(n_9654));
 AOI22xp33_ASAP7_75t_SL g165300 (.A1(n_1167),
    .A2(\u11_mem[1] [13]),
    .B1(n_46233),
    .B2(\u11_mem[3] [13]),
    .Y(n_9663));
 AOI22xp33_ASAP7_75t_SL g165302 (.A1(n_1167),
    .A2(\u11_mem[1] [28]),
    .B1(n_46233),
    .B2(\u11_mem[3] [28]),
    .Y(n_9665));
 AOI22xp33_ASAP7_75t_SL g165319 (.A1(n_1171),
    .A2(\u9_mem[1] [19]),
    .B1(n_22780),
    .B2(\u9_mem[3] [19]),
    .Y(n_9682));
 AOI22xp33_ASAP7_75t_SL g165323 (.A1(n_1171),
    .A2(\u9_mem[1] [14]),
    .B1(n_22780),
    .B2(\u9_mem[3] [14]),
    .Y(n_9686));
 AOI22xp33_ASAP7_75t_SL g165337 (.A1(n_1171),
    .A2(\u9_mem[1] [22]),
    .B1(n_22780),
    .B2(\u9_mem[3] [22]),
    .Y(n_9701));
 AOI22xp33_ASAP7_75t_SL g165339 (.A1(n_1171),
    .A2(\u9_mem[1] [7]),
    .B1(n_22780),
    .B2(\u9_mem[3] [7]),
    .Y(n_9703));
 AOI22xp5_ASAP7_75t_SL g165344 (.A1(n_11128),
    .A2(n_66004),
    .B1(\u5_mem[3] [6]),
    .B2(n_9476),
    .Y(n_9711));
 AOI22xp5_ASAP7_75t_SL g165346 (.A1(n_3420),
    .A2(n_66004),
    .B1(\u6_mem[0] [6]),
    .B2(n_3425),
    .Y(n_9713));
 AOI22xp5_ASAP7_75t_SL g165350 (.A1(n_66004),
    .A2(n_32163),
    .B1(\u5_mem[1] [6]),
    .B2(n_13500),
    .Y(n_9717));
 AOI22xp5_ASAP7_75t_SL g165354 (.A1(n_66004),
    .A2(n_3461),
    .B1(\u8_mem[0] [6]),
    .B2(n_3460),
    .Y(n_9721));
 AOI22xp5_ASAP7_75t_SL g165355 (.A1(n_3320),
    .A2(n_32644),
    .B1(\u8_mem[2] [6]),
    .B2(n_16908),
    .Y(n_9722));
 AOI22xp5_ASAP7_75t_SL g165356 (.A1(n_3285),
    .A2(n_66005),
    .B1(\u5_mem[2] [6]),
    .B2(n_43020),
    .Y(n_9723));
 AOI22xp5_ASAP7_75t_SL g165359 (.A1(n_3188),
    .A2(n_32644),
    .B1(\u7_mem[2] [6]),
    .B2(n_13325),
    .Y(n_9726));
 AOI22xp5_ASAP7_75t_SL g165360 (.A1(n_24633),
    .A2(n_66005),
    .B1(\u4_mem[2] [6]),
    .B2(n_13304),
    .Y(n_9727));
 AOI21xp5_ASAP7_75t_SL g165364 (.A1(n_16797),
    .A2(n_66005),
    .B(n_26581),
    .Y(n_9731));
 AOI22xp5_ASAP7_75t_SL g165371 (.A1(n_11126),
    .A2(n_66032),
    .B1(\u5_mem[3] [14]),
    .B2(n_9476),
    .Y(n_9738));
 AOI22xp33_ASAP7_75t_SL g165375 (.A1(n_3420),
    .A2(n_28251),
    .B1(\u6_mem[0] [14]),
    .B2(n_3415),
    .Y(n_9742));
 AOI22xp5_ASAP7_75t_SL g165378 (.A1(n_66032),
    .A2(n_32164),
    .B1(\u5_mem[1] [14]),
    .B2(n_13508),
    .Y(n_9745));
 AOI22xp5_ASAP7_75t_SL g165380 (.A1(n_66032),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [14]),
    .Y(n_9747));
 AOI22xp5_ASAP7_75t_SL g165384 (.A1(n_3320),
    .A2(n_28251),
    .B1(\u8_mem[2] [14]),
    .B2(n_16900),
    .Y(n_9751));
 AOI22xp5_ASAP7_75t_SL g165385 (.A1(n_3285),
    .A2(n_28251),
    .B1(\u5_mem[2] [14]),
    .B2(n_43020),
    .Y(n_9752));
 AOI22xp5_ASAP7_75t_SL g165388 (.A1(n_3188),
    .A2(n_66032),
    .B1(\u7_mem[2] [14]),
    .B2(n_13333),
    .Y(n_9755));
 AOI22xp5_ASAP7_75t_SL g165389 (.A1(n_24633),
    .A2(n_28251),
    .B1(\u4_mem[2] [14]),
    .B2(n_13312),
    .Y(n_9756));
 AOI22xp5_ASAP7_75t_SL g165390 (.A1(n_66032),
    .A2(n_3454),
    .B1(\u8_mem[0] [14]),
    .B2(n_3453),
    .Y(n_9757));
 AOI21xp5_ASAP7_75t_SL g165393 (.A1(n_16797),
    .A2(n_28251),
    .B(n_2639),
    .Y(n_9760));
 AOI22xp5_ASAP7_75t_SL g165400 (.A1(n_28913),
    .A2(n_11128),
    .B1(\u5_mem[3] [15]),
    .B2(n_9476),
    .Y(n_9767));
 AOI22xp5_ASAP7_75t_SL g165405 (.A1(n_3420),
    .A2(n_28913),
    .B1(\u6_mem[0] [15]),
    .B2(n_3415),
    .Y(n_9772));
 AOI22xp5_ASAP7_75t_SL g165407 (.A1(n_28913),
    .A2(n_32163),
    .B1(\u5_mem[1] [15]),
    .B2(n_13508),
    .Y(n_9774));
 AOI22xp5_ASAP7_75t_SL g165409 (.A1(n_28913),
    .A2(n_14386),
    .B1(n_31741),
    .B2(\u6_mem[1] [15]),
    .Y(n_9776));
 AOI22xp5_ASAP7_75t_SL g165413 (.A1(n_3320),
    .A2(n_28913),
    .B1(\u8_mem[2] [15]),
    .B2(n_16908),
    .Y(n_9780));
 AOI22xp5_ASAP7_75t_SL g165414 (.A1(n_3285),
    .A2(n_28913),
    .B1(\u5_mem[2] [15]),
    .B2(n_43028),
    .Y(n_9781));
 AOI22xp5_ASAP7_75t_SL g165417 (.A1(n_3188),
    .A2(n_28913),
    .B1(\u7_mem[2] [15]),
    .B2(n_13333),
    .Y(n_9784));
 AOI22xp5_ASAP7_75t_SL g165418 (.A1(n_24633),
    .A2(n_28913),
    .B1(\u4_mem[2] [15]),
    .B2(n_13312),
    .Y(n_9785));
 AOI22xp5_ASAP7_75t_SL g165419 (.A1(n_28913),
    .A2(n_3461),
    .B1(\u8_mem[0] [15]),
    .B2(n_3453),
    .Y(n_9786));
 AOI21xp5_ASAP7_75t_SL g165423 (.A1(n_16797),
    .A2(n_65990),
    .B(n_2642),
    .Y(n_9790));
 AOI22xp5_ASAP7_75t_SL g165433 (.A1(n_11126),
    .A2(n_65969),
    .B1(\u5_mem[3] [7]),
    .B2(n_9476),
    .Y(n_9800));
 AOI22xp5_ASAP7_75t_SL g165435 (.A1(n_65969),
    .A2(n_3420),
    .B1(\u6_mem[0] [7]),
    .B2(n_3425),
    .Y(n_9802));
 AOI22xp5_ASAP7_75t_SL g165437 (.A1(n_65969),
    .A2(n_32163),
    .B1(\u5_mem[1] [7]),
    .B2(n_13508),
    .Y(n_9804));
 AOI22xp5_ASAP7_75t_SL g165441 (.A1(n_65969),
    .A2(n_3461),
    .B1(\u8_mem[0] [7]),
    .B2(n_3460),
    .Y(n_9808));
 AOI22xp5_ASAP7_75t_SL g165443 (.A1(n_3320),
    .A2(n_65969),
    .B1(\u8_mem[2] [7]),
    .B2(n_16900),
    .Y(n_9810));
 AOI22xp5_ASAP7_75t_SL g165444 (.A1(n_3285),
    .A2(n_17578),
    .B1(\u5_mem[2] [7]),
    .B2(n_43020),
    .Y(n_9811));
 AOI22xp5_ASAP7_75t_SL g165447 (.A1(n_3188),
    .A2(n_65969),
    .B1(\u7_mem[2] [7]),
    .B2(n_13333),
    .Y(n_9814));
 AOI22xp5_ASAP7_75t_SL g165448 (.A1(n_24633),
    .A2(n_17578),
    .B1(\u4_mem[2] [7]),
    .B2(n_13312),
    .Y(n_9815));
 AOI21xp5_ASAP7_75t_SL g165450 (.A1(n_16797),
    .A2(n_17578),
    .B(n_2643),
    .Y(n_9817));
 AOI22xp5_ASAP7_75t_SL g165461 (.A1(n_11128),
    .A2(n_28330),
    .B1(\u5_mem[3] [2]),
    .B2(n_9476),
    .Y(n_9828));
 AOI22xp5_ASAP7_75t_SL g165465 (.A1(n_3420),
    .A2(n_28330),
    .B1(\u6_mem[0] [2]),
    .B2(n_3425),
    .Y(n_9832));
 AOI22xp5_ASAP7_75t_SL g165467 (.A1(n_28330),
    .A2(n_32164),
    .B1(\u5_mem[1] [2]),
    .B2(n_13500),
    .Y(n_9834));
 AOI22xp5_ASAP7_75t_SL g165471 (.A1(n_28330),
    .A2(n_3454),
    .B1(\u8_mem[0] [2]),
    .B2(n_3460),
    .Y(n_9838));
 AOI22xp5_ASAP7_75t_SL g165473 (.A1(n_3320),
    .A2(n_28330),
    .B1(\u8_mem[2] [2]),
    .B2(n_16908),
    .Y(n_9840));
 AOI22xp5_ASAP7_75t_SL g165474 (.A1(n_3285),
    .A2(n_66000),
    .B1(\u5_mem[2] [2]),
    .B2(n_43028),
    .Y(n_9841));
 AOI22xp5_ASAP7_75t_SL g165476 (.A1(n_3188),
    .A2(n_66000),
    .B1(\u7_mem[2] [2]),
    .B2(n_13325),
    .Y(n_9843));
 AOI22xp5_ASAP7_75t_SL g165477 (.A1(n_24633),
    .A2(n_28330),
    .B1(\u4_mem[2] [2]),
    .B2(n_13304),
    .Y(n_9844));
 AOI21xp5_ASAP7_75t_SL g165482 (.A1(n_16797),
    .A2(n_66000),
    .B(n_2595),
    .Y(n_9849));
 AOI22xp5_ASAP7_75t_SL g165490 (.A1(n_11128),
    .A2(n_66855),
    .B1(\u5_mem[3] [3]),
    .B2(n_9476),
    .Y(n_9857));
 AOI22xp5_ASAP7_75t_SL g165493 (.A1(n_3420),
    .A2(n_15867),
    .B1(\u6_mem[0] [3]),
    .B2(n_3415),
    .Y(n_9860));
 AOI22xp5_ASAP7_75t_SL g165496 (.A1(n_66855),
    .A2(n_32163),
    .B1(\u5_mem[1] [3]),
    .B2(n_13500),
    .Y(n_9863));
 AOI22xp5_ASAP7_75t_SL g165500 (.A1(n_66855),
    .A2(n_3461),
    .B1(\u8_mem[0] [3]),
    .B2(n_3460),
    .Y(n_9867));
 AOI22xp5_ASAP7_75t_SL g165502 (.A1(n_3320),
    .A2(n_66855),
    .B1(\u8_mem[2] [3]),
    .B2(n_16908),
    .Y(n_9869));
 AOI22xp5_ASAP7_75t_SL g165503 (.A1(n_3285),
    .A2(n_15867),
    .B1(\u5_mem[2] [3]),
    .B2(n_43028),
    .Y(n_9870));
 AOI22xp5_ASAP7_75t_SL g165506 (.A1(n_3188),
    .A2(n_66856),
    .B1(\u7_mem[2] [3]),
    .B2(n_13333),
    .Y(n_9873));
 AOI22xp5_ASAP7_75t_SL g165507 (.A1(n_24633),
    .A2(n_15867),
    .B1(\u4_mem[2] [3]),
    .B2(n_13304),
    .Y(n_9874));
 AOI21xp5_ASAP7_75t_SL g165510 (.A1(n_16797),
    .A2(n_66856),
    .B(n_2608),
    .Y(n_9877));
 AOI22xp5_ASAP7_75t_SL g165519 (.A1(n_11126),
    .A2(n_28240),
    .B1(\u5_mem[3] [8]),
    .B2(n_9476),
    .Y(n_9886));
 AOI22xp5_ASAP7_75t_SL g165522 (.A1(n_3420),
    .A2(n_65980),
    .B1(\u6_mem[0] [8]),
    .B2(n_3415),
    .Y(n_9889));
 AOI22xp5_ASAP7_75t_SL g165525 (.A1(n_28240),
    .A2(n_32163),
    .B1(\u5_mem[1] [8]),
    .B2(n_13508),
    .Y(n_9892));
 AOI22xp5_ASAP7_75t_SL g165529 (.A1(n_28240),
    .A2(n_3461),
    .B1(\u8_mem[0] [8]),
    .B2(n_3453),
    .Y(n_9896));
 AOI22xp5_ASAP7_75t_SL g165531 (.A1(n_3320),
    .A2(n_28240),
    .B1(\u8_mem[2] [8]),
    .B2(n_16908),
    .Y(n_9898));
 AOI22xp5_ASAP7_75t_SL g165532 (.A1(n_3285),
    .A2(n_65980),
    .B1(\u5_mem[2] [8]),
    .B2(n_43020),
    .Y(n_9899));
 AOI22xp5_ASAP7_75t_SL g165535 (.A1(n_3188),
    .A2(n_28240),
    .B1(\u7_mem[2] [8]),
    .B2(n_13333),
    .Y(n_9902));
 AOI22xp33_ASAP7_75t_SL g165536 (.A1(n_24633),
    .A2(n_65980),
    .B1(\u4_mem[2] [8]),
    .B2(n_13312),
    .Y(n_9903));
 AOI21xp5_ASAP7_75t_SL g165540 (.A1(n_16797),
    .A2(n_65980),
    .B(n_17688),
    .Y(n_9907));
 AOI22xp5_ASAP7_75t_SL g165546 (.A1(n_11128),
    .A2(n_65975),
    .B1(\u5_mem[3] [10]),
    .B2(n_9476),
    .Y(n_9914));
 AOI22xp5_ASAP7_75t_SL g165555 (.A1(n_65975),
    .A2(n_14386),
    .B1(\u6_mem[1] [10]),
    .B2(n_31741),
    .Y(n_9922));
 AOI22xp33_ASAP7_75t_SL g165559 (.A1(n_3320),
    .A2(n_65975),
    .B1(\u8_mem[2] [10]),
    .B2(n_16908),
    .Y(n_9926));
 AOI22xp5_ASAP7_75t_SL g165563 (.A1(n_3188),
    .A2(n_65972),
    .B1(\u7_mem[2] [10]),
    .B2(n_13325),
    .Y(n_9930));
 AOI21xp5_ASAP7_75t_SL g165569 (.A1(n_16797),
    .A2(n_65975),
    .B(n_2573),
    .Y(n_9936));
 AOI22xp33_ASAP7_75t_SL g165574 (.A1(n_3420),
    .A2(n_79972),
    .B1(\u6_mem[0] [9]),
    .B2(n_3415),
    .Y(n_9941));
 AOI22xp5_ASAP7_75t_SL g165577 (.A1(n_11126),
    .A2(n_79972),
    .B1(\u5_mem[3] [9]),
    .B2(n_9476),
    .Y(n_9944));
 AOI22xp5_ASAP7_75t_SL g165582 (.A1(n_9942),
    .A2(n_32164),
    .B1(\u5_mem[1] [9]),
    .B2(n_13508),
    .Y(n_9949));
 AOI22xp5_ASAP7_75t_SL g165587 (.A1(n_3320),
    .A2(n_79971),
    .B1(\u8_mem[2] [9]),
    .B2(n_16908),
    .Y(n_9954));
 AOI22xp5_ASAP7_75t_SL g165590 (.A1(n_3188),
    .A2(n_9942),
    .B1(\u7_mem[2] [9]),
    .B2(n_13325),
    .Y(n_9957));
 AOI22xp5_ASAP7_75t_SL g165591 (.A1(n_24633),
    .A2(n_79972),
    .B1(\u4_mem[2] [9]),
    .B2(n_13312),
    .Y(n_9958));
 AOI22xp5_ASAP7_75t_SL g165592 (.A1(n_9942),
    .A2(n_3461),
    .B1(\u8_mem[0] [9]),
    .B2(n_3460),
    .Y(n_9959));
 AOI22xp5_ASAP7_75t_SL g165593 (.A1(n_3285),
    .A2(n_79971),
    .B1(\u5_mem[2] [9]),
    .B2(n_43028),
    .Y(n_9960));
 AOI21xp5_ASAP7_75t_SL g165596 (.A1(n_16797),
    .A2(n_9942),
    .B(n_2646),
    .Y(n_9963));
 AOI22xp5_ASAP7_75t_SL g165633 (.A1(n_11128),
    .A2(n_10000),
    .B1(\u5_mem[3] [11]),
    .B2(n_9476),
    .Y(n_10001));
 AOI22xp5_ASAP7_75t_SL g165638 (.A1(n_3420),
    .A2(n_10000),
    .B1(\u6_mem[0] [11]),
    .B2(n_3415),
    .Y(n_10005));
 AOI22xp5_ASAP7_75t_SL g165640 (.A1(n_10000),
    .A2(n_32163),
    .B1(\u5_mem[1] [11]),
    .B2(n_13500),
    .Y(n_10007));
 AOI22xp5_ASAP7_75t_SL g165642 (.A1(n_10000),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [11]),
    .Y(n_10009));
 AOI22xp5_ASAP7_75t_SL g165646 (.A1(n_3320),
    .A2(n_10000),
    .B1(\u8_mem[2] [11]),
    .B2(n_16908),
    .Y(n_10013));
 AOI22xp5_ASAP7_75t_SL g165647 (.A1(n_3285),
    .A2(n_66842),
    .B1(\u5_mem[2] [11]),
    .B2(n_43028),
    .Y(n_10014));
 AOI22xp5_ASAP7_75t_SL g165650 (.A1(n_3188),
    .A2(n_10000),
    .B1(\u7_mem[2] [11]),
    .B2(n_13333),
    .Y(n_10017));
 AOI22xp5_ASAP7_75t_SL g165651 (.A1(n_24633),
    .A2(n_66842),
    .B1(\u4_mem[2] [11]),
    .B2(n_13312),
    .Y(n_10018));
 AOI22xp5_ASAP7_75t_SL g165652 (.A1(n_10000),
    .A2(n_3454),
    .B1(\u8_mem[0] [11]),
    .B2(n_3453),
    .Y(n_10019));
 AOI21xp5_ASAP7_75t_SL g165655 (.A1(n_16797),
    .A2(n_66843),
    .B(n_2610),
    .Y(n_10022));
 AOI22xp5_ASAP7_75t_SL g165662 (.A1(n_11126),
    .A2(n_65997),
    .B1(\u5_mem[3] [12]),
    .B2(n_9476),
    .Y(n_10030));
 AOI22xp5_ASAP7_75t_SL g165667 (.A1(n_3420),
    .A2(n_65997),
    .B1(\u6_mem[0] [12]),
    .B2(n_3415),
    .Y(n_10034));
 AOI22xp5_ASAP7_75t_SL g165669 (.A1(n_65997),
    .A2(n_32164),
    .B1(\u5_mem[1] [12]),
    .B2(n_13500),
    .Y(n_10036));
 AOI22xp5_ASAP7_75t_SL g165671 (.A1(n_65997),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [12]),
    .Y(n_10038));
 AOI22xp5_ASAP7_75t_SL g165675 (.A1(n_3320),
    .A2(n_65997),
    .B1(\u8_mem[2] [12]),
    .B2(n_16908),
    .Y(n_10042));
 AOI22xp5_ASAP7_75t_SL g165676 (.A1(n_3285),
    .A2(n_10026),
    .B1(\u5_mem[2] [12]),
    .B2(n_43028),
    .Y(n_10043));
 AOI22xp5_ASAP7_75t_SL g165679 (.A1(n_3188),
    .A2(n_65997),
    .B1(\u7_mem[2] [12]),
    .B2(n_13325),
    .Y(n_10046));
 AOI22xp5_ASAP7_75t_SL g165680 (.A1(n_24633),
    .A2(n_10026),
    .B1(\u4_mem[2] [12]),
    .B2(n_13304),
    .Y(n_10047));
 AOI22xp5_ASAP7_75t_SL g165681 (.A1(n_65997),
    .A2(n_3461),
    .B1(\u8_mem[0] [12]),
    .B2(n_3453),
    .Y(n_10048));
 AOI21xp5_ASAP7_75t_SL g165683 (.A1(n_16797),
    .A2(n_65997),
    .B(n_2624),
    .Y(n_10050));
 AOI22xp33_ASAP7_75t_SL g165690 (.A1(n_3420),
    .A2(n_66869),
    .B1(\u6_mem[0] [5]),
    .B2(n_3425),
    .Y(n_10057));
 AOI22xp5_ASAP7_75t_SL g165694 (.A1(n_11126),
    .A2(n_10058),
    .B1(\u5_mem[3] [5]),
    .B2(n_9476),
    .Y(n_10061));
 AOI22xp5_ASAP7_75t_SL g165698 (.A1(n_10058),
    .A2(n_32164),
    .B1(\u5_mem[1] [5]),
    .B2(n_13508),
    .Y(n_10065));
 AOI22xp5_ASAP7_75t_SL g165702 (.A1(n_10058),
    .A2(n_3461),
    .B1(\u8_mem[0] [5]),
    .B2(n_3453),
    .Y(n_10069));
 AOI22xp5_ASAP7_75t_SL g165704 (.A1(n_3320),
    .A2(n_10058),
    .B1(\u8_mem[2] [5]),
    .B2(n_16900),
    .Y(n_10071));
 AOI22xp5_ASAP7_75t_SL g165705 (.A1(n_3285),
    .A2(n_66869),
    .B1(\u5_mem[2] [5]),
    .B2(n_43028),
    .Y(n_10072));
 AOI22xp5_ASAP7_75t_SL g165708 (.A1(n_3188),
    .A2(n_10058),
    .B1(\u7_mem[2] [5]),
    .B2(n_13325),
    .Y(n_10075));
 AOI22xp5_ASAP7_75t_SL g165709 (.A1(n_24633),
    .A2(n_66869),
    .B1(\u4_mem[2] [5]),
    .B2(n_13312),
    .Y(n_10076));
 AOI21xp5_ASAP7_75t_SL g165712 (.A1(n_16797),
    .A2(n_10058),
    .B(n_2647),
    .Y(n_10079));
 AOI22xp5_ASAP7_75t_SL g165722 (.A1(n_11126),
    .A2(n_65955),
    .B1(\u5_mem[3] [13]),
    .B2(n_9476),
    .Y(n_10089));
 AOI22xp5_ASAP7_75t_SL g165725 (.A1(n_3420),
    .A2(n_35041),
    .B1(\u6_mem[0] [13]),
    .B2(n_3415),
    .Y(n_10092));
 AOI22xp5_ASAP7_75t_SL g165727 (.A1(n_35041),
    .A2(n_32164),
    .B1(\u5_mem[1] [13]),
    .B2(n_13500),
    .Y(n_10094));
 AOI22xp5_ASAP7_75t_SL g165732 (.A1(n_3320),
    .A2(n_65955),
    .B1(\u8_mem[2] [13]),
    .B2(n_16908),
    .Y(n_10099));
 AOI22xp5_ASAP7_75t_SL g165733 (.A1(n_3285),
    .A2(n_35041),
    .B1(\u5_mem[2] [13]),
    .B2(n_43020),
    .Y(n_10100));
 AOI22xp5_ASAP7_75t_SL g165736 (.A1(n_3188),
    .A2(n_65955),
    .B1(\u7_mem[2] [13]),
    .B2(n_13333),
    .Y(n_10103));
 AOI22xp5_ASAP7_75t_SL g165737 (.A1(n_24633),
    .A2(n_35041),
    .B1(\u4_mem[2] [13]),
    .B2(n_13312),
    .Y(n_10104));
 AOI22xp5_ASAP7_75t_SL g165738 (.A1(n_65955),
    .A2(n_3454),
    .B1(\u8_mem[0] [13]),
    .B2(n_3460),
    .Y(n_10105));
 AOI21xp5_ASAP7_75t_SL g165740 (.A1(n_16797),
    .A2(n_65955),
    .B(n_2660),
    .Y(n_10107));
 AOI22xp5_ASAP7_75t_SL g165752 (.A1(n_3420),
    .A2(n_28276),
    .B1(\u6_mem[0] [16]),
    .B2(n_3415),
    .Y(n_10119));
 AOI22xp5_ASAP7_75t_SL g165755 (.A1(n_65949),
    .A2(n_32164),
    .B1(\u5_mem[1] [16]),
    .B2(n_13508),
    .Y(n_10122));
 AOI22xp5_ASAP7_75t_SL g165757 (.A1(n_65949),
    .A2(n_14386),
    .B1(\u6_mem[1] [16]),
    .B2(n_22396),
    .Y(n_10124));
 AOI22xp5_ASAP7_75t_SL g165761 (.A1(n_3320),
    .A2(n_65949),
    .B1(\u8_mem[2] [16]),
    .B2(n_16908),
    .Y(n_10128));
 AOI22xp5_ASAP7_75t_SL g165762 (.A1(n_3285),
    .A2(n_28276),
    .B1(\u5_mem[2] [16]),
    .B2(n_43028),
    .Y(n_10129));
 AOI22xp5_ASAP7_75t_SL g165765 (.A1(n_3188),
    .A2(n_65949),
    .B1(\u7_mem[2] [16]),
    .B2(n_13325),
    .Y(n_10132));
 AOI22xp5_ASAP7_75t_SL g165766 (.A1(n_24633),
    .A2(n_28276),
    .B1(\u4_mem[2] [16]),
    .B2(n_13312),
    .Y(n_10133));
 AOI22xp5_ASAP7_75t_SL g165767 (.A1(n_65949),
    .A2(n_3454),
    .B1(\u8_mem[0] [16]),
    .B2(n_3460),
    .Y(n_10134));
 AOI21xp5_ASAP7_75t_SL g165771 (.A1(n_16797),
    .A2(n_65949),
    .B(n_2650),
    .Y(n_10138));
 AOI22xp5_ASAP7_75t_SL g165779 (.A1(n_3420),
    .A2(n_10143),
    .B1(\u6_mem[0] [17]),
    .B2(n_3415),
    .Y(n_10146));
 AOI22xp5_ASAP7_75t_SL g165784 (.A1(n_65952),
    .A2(n_32163),
    .B1(\u5_mem[1] [17]),
    .B2(n_13500),
    .Y(n_10151));
 AOI22xp5_ASAP7_75t_SL g165789 (.A1(n_3320),
    .A2(n_10143),
    .B1(\u8_mem[2] [17]),
    .B2(n_16908),
    .Y(n_10156));
 AOI22xp5_ASAP7_75t_SL g165790 (.A1(n_3285),
    .A2(n_65952),
    .B1(\u5_mem[2] [17]),
    .B2(n_43028),
    .Y(n_10157));
 AOI22xp33_ASAP7_75t_SL g165793 (.A1(n_3188),
    .A2(n_10143),
    .B1(\u7_mem[2] [17]),
    .B2(n_13325),
    .Y(n_10160));
 AOI22xp5_ASAP7_75t_SL g165794 (.A1(n_24633),
    .A2(n_65952),
    .B1(\u4_mem[2] [17]),
    .B2(n_13312),
    .Y(n_10161));
 AOI22xp5_ASAP7_75t_SL g165795 (.A1(n_10143),
    .A2(n_3454),
    .B1(\u8_mem[0] [17]),
    .B2(n_3453),
    .Y(n_10162));
 AOI21xp5_ASAP7_75t_SL g165798 (.A1(n_16797),
    .A2(n_65952),
    .B(n_2641),
    .Y(n_10165));
 AOI22xp5_ASAP7_75t_SL g165805 (.A1(n_3420),
    .A2(n_10194),
    .B1(\u6_mem[0] [18]),
    .B2(n_3425),
    .Y(n_10175));
 AOI22xp5_ASAP7_75t_SL g165807 (.A1(n_10194),
    .A2(n_32164),
    .B1(\u5_mem[1] [18]),
    .B2(n_13508),
    .Y(n_10177));
 AOI22xp5_ASAP7_75t_SL g165812 (.A1(n_3320),
    .A2(n_10171),
    .B1(\u8_mem[2] [18]),
    .B2(n_16908),
    .Y(n_10182));
 AOI22xp5_ASAP7_75t_SL g165813 (.A1(n_3285),
    .A2(n_10194),
    .B1(\u5_mem[2] [18]),
    .B2(n_43028),
    .Y(n_10183));
 AOI22xp5_ASAP7_75t_SL g165816 (.A1(n_3188),
    .A2(n_10171),
    .B1(\u7_mem[2] [18]),
    .B2(n_13325),
    .Y(n_10186));
 AOI22xp5_ASAP7_75t_SL g165817 (.A1(n_24633),
    .A2(n_10194),
    .B1(\u4_mem[2] [18]),
    .B2(n_13312),
    .Y(n_10187));
 AOI22xp5_ASAP7_75t_SL g165818 (.A1(n_10171),
    .A2(n_3454),
    .B1(\u8_mem[0] [18]),
    .B2(n_3460),
    .Y(n_10188));
 AOI21xp5_ASAP7_75t_SL g165822 (.A1(n_16797),
    .A2(n_10171),
    .B(n_2611),
    .Y(n_10192));
 AOI22xp5_ASAP7_75t_SL g165832 (.A1(n_3420),
    .A2(n_10196),
    .B1(\u6_mem[0] [19]),
    .B2(n_3425),
    .Y(n_10202));
 AOI22xp5_ASAP7_75t_SL g165833 (.A1(n_10198),
    .A2(n_73997),
    .B1(\u8_mem[1] [19]),
    .B2(n_73399),
    .Y(n_10203));
 AOI22xp5_ASAP7_75t_SL g165834 (.A1(n_10196),
    .A2(n_32164),
    .B1(\u5_mem[1] [19]),
    .B2(n_13508),
    .Y(n_10204));
 AOI22xp5_ASAP7_75t_SL g165839 (.A1(n_3320),
    .A2(n_10198),
    .B1(\u8_mem[2] [19]),
    .B2(n_16908),
    .Y(n_10209));
 AOI22xp5_ASAP7_75t_SL g165840 (.A1(n_3285),
    .A2(n_10196),
    .B1(\u5_mem[2] [19]),
    .B2(n_43028),
    .Y(n_10210));
 AOI22xp5_ASAP7_75t_SL g165843 (.A1(n_3188),
    .A2(n_10198),
    .B1(\u7_mem[2] [19]),
    .B2(n_13325),
    .Y(n_10213));
 AOI22xp5_ASAP7_75t_SL g165844 (.A1(n_24633),
    .A2(n_10196),
    .B1(\u4_mem[2] [19]),
    .B2(n_13312),
    .Y(n_10214));
 AOI22xp5_ASAP7_75t_SL g165845 (.A1(n_10198),
    .A2(n_3461),
    .B1(\u8_mem[0] [19]),
    .B2(n_3460),
    .Y(n_10215));
 AOI21xp5_ASAP7_75t_SL g165848 (.A1(n_16797),
    .A2(n_10196),
    .B(n_2609),
    .Y(n_10218));
 AOI22xp5_ASAP7_75t_SL g165857 (.A1(n_3320),
    .A2(n_66026),
    .B1(\u8_mem[2] [20]),
    .B2(n_16900),
    .Y(n_10227));
 AOI22xp5_ASAP7_75t_SL g165860 (.A1(n_3420),
    .A2(n_33024),
    .B1(\u6_mem[0] [20]),
    .B2(n_3425),
    .Y(n_10230));
 AOI22xp5_ASAP7_75t_SL g165861 (.A1(n_10247),
    .A2(n_32163),
    .B1(\u5_mem[1] [20]),
    .B2(n_13500),
    .Y(n_10231));
 AOI22xp5_ASAP7_75t_SL g165864 (.A1(n_33024),
    .A2(n_14386),
    .B1(\u6_mem[1] [20]),
    .B2(n_31741),
    .Y(n_10234));
 AOI22xp5_ASAP7_75t_SL g165868 (.A1(n_3285),
    .A2(n_33024),
    .B1(\u5_mem[2] [20]),
    .B2(n_43028),
    .Y(n_10238));
 AOI22xp5_ASAP7_75t_SL g165870 (.A1(n_3188),
    .A2(n_33024),
    .B1(\u7_mem[2] [20]),
    .B2(n_13333),
    .Y(n_10240));
 AOI22xp5_ASAP7_75t_SL g165871 (.A1(n_24633),
    .A2(n_66026),
    .B1(\u4_mem[2] [20]),
    .B2(n_13312),
    .Y(n_10241));
 AOI22xp5_ASAP7_75t_SL g165872 (.A1(n_33024),
    .A2(n_3454),
    .B1(\u8_mem[0] [20]),
    .B2(n_3453),
    .Y(n_10242));
 AOI21xp5_ASAP7_75t_SL g165874 (.A1(n_16797),
    .A2(n_66026),
    .B(n_2623),
    .Y(n_10244));
 AOI22xp5_ASAP7_75t_SL g165884 (.A1(n_3320),
    .A2(n_73996),
    .B1(\u8_mem[2] [21]),
    .B2(n_16900),
    .Y(n_10254));
 AOI22xp5_ASAP7_75t_SL g165887 (.A1(n_3420),
    .A2(n_32916),
    .B1(\u6_mem[0] [21]),
    .B2(n_3425),
    .Y(n_10257));
 AOI22xp5_ASAP7_75t_SL g165889 (.A1(n_32916),
    .A2(n_16009),
    .B1(\u3_mem[1] [21]),
    .B2(n_22505),
    .Y(n_10259));
 AOI22xp5_ASAP7_75t_SL g165890 (.A1(n_66016),
    .A2(n_32163),
    .B1(\u5_mem[1] [21]),
    .B2(n_13508),
    .Y(n_10260));
 AOI22xp5_ASAP7_75t_SL g165895 (.A1(n_3285),
    .A2(n_32916),
    .B1(\u5_mem[2] [21]),
    .B2(n_43020),
    .Y(n_10265));
 AOI22xp5_ASAP7_75t_SL g165897 (.A1(n_3188),
    .A2(n_32916),
    .B1(\u7_mem[2] [21]),
    .B2(n_13325),
    .Y(n_10267));
 AOI22xp5_ASAP7_75t_SL g165898 (.A1(n_24633),
    .A2(n_73996),
    .B1(\u4_mem[2] [21]),
    .B2(n_13312),
    .Y(n_10268));
 AOI22xp5_ASAP7_75t_SL g165899 (.A1(n_32916),
    .A2(n_3454),
    .B1(\u8_mem[0] [21]),
    .B2(n_3453),
    .Y(n_10269));
 AOI21xp5_ASAP7_75t_SL g165902 (.A1(n_16797),
    .A2(n_73996),
    .B(n_2620),
    .Y(n_10272));
 AOI22xp5_ASAP7_75t_SL g165918 (.A1(n_65941),
    .A2(n_14386),
    .B1(\u6_mem[1] [22]),
    .B2(n_31741),
    .Y(n_10288));
 AOI22xp5_ASAP7_75t_SL g165922 (.A1(n_3285),
    .A2(n_65941),
    .B1(\u5_mem[2] [22]),
    .B2(n_43028),
    .Y(n_10292));
 BUFx2_ASAP7_75t_R g165932 (.A(n_65937),
    .Y(n_10302));
 AOI22xp5_ASAP7_75t_SL g165936 (.A1(n_3320),
    .A2(n_65930),
    .B1(\u8_mem[2] [23]),
    .B2(n_16900),
    .Y(n_10306));
 AOI22xp5_ASAP7_75t_SL g165940 (.A1(n_3420),
    .A2(n_28381),
    .B1(\u6_mem[0] [23]),
    .B2(n_3415),
    .Y(n_10310));
 AOI22xp5_ASAP7_75t_SL g165945 (.A1(n_65930),
    .A2(n_32164),
    .B1(n_13500),
    .B2(\u5_mem[1] [23]),
    .Y(n_10315));
 AOI22xp5_ASAP7_75t_SL g165947 (.A1(n_65930),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [23]),
    .Y(n_10317));
 AOI22xp5_ASAP7_75t_SL g165951 (.A1(n_3285),
    .A2(n_65930),
    .B1(\u5_mem[2] [23]),
    .B2(n_43020),
    .Y(n_10321));
 AOI22xp5_ASAP7_75t_SL g165953 (.A1(n_3188),
    .A2(n_65930),
    .B1(\u7_mem[2] [23]),
    .B2(n_13333),
    .Y(n_10323));
 AOI22xp5_ASAP7_75t_SL g165954 (.A1(n_24633),
    .A2(n_28381),
    .B1(\u4_mem[2] [23]),
    .B2(n_13304),
    .Y(n_10324));
 AOI22xp5_ASAP7_75t_SL g165956 (.A1(n_28381),
    .A2(n_3454),
    .B1(\u8_mem[0] [23]),
    .B2(n_3460),
    .Y(n_10326));
 AOI21xp5_ASAP7_75t_SL g165957 (.A1(n_16797),
    .A2(n_65930),
    .B(n_2619),
    .Y(n_10327));
 BUFx2_ASAP7_75t_R g165959 (.A(n_65929),
    .Y(n_10329));
 AOI22xp5_ASAP7_75t_SL g165965 (.A1(n_3285),
    .A2(n_65902),
    .B1(\u5_mem[2] [31]),
    .B2(n_43020),
    .Y(n_10335));
 AOI22xp5_ASAP7_75t_SL g165966 (.A1(n_3320),
    .A2(n_65902),
    .B1(\u8_mem[2] [31]),
    .B2(n_16900),
    .Y(n_10336));
 AOI22xp5_ASAP7_75t_SL g165969 (.A1(n_3420),
    .A2(n_15920),
    .B1(\u6_mem[0] [31]),
    .B2(n_3425),
    .Y(n_10339));
 AOI22xp5_ASAP7_75t_SL g165974 (.A1(n_65902),
    .A2(n_32164),
    .B1(\u5_mem[1] [31]),
    .B2(n_13500),
    .Y(n_10344));
 AOI22xp5_ASAP7_75t_SL g165976 (.A1(n_15920),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [31]),
    .Y(n_10346));
 AOI22xp5_ASAP7_75t_SL g165980 (.A1(n_3188),
    .A2(n_65902),
    .B1(\u7_mem[2] [31]),
    .B2(n_13333),
    .Y(n_10350));
 AOI22xp5_ASAP7_75t_SL g165981 (.A1(n_24633),
    .A2(n_15920),
    .B1(\u4_mem[2] [31]),
    .B2(n_13304),
    .Y(n_10351));
 AOI22xp5_ASAP7_75t_SL g165982 (.A1(n_65900),
    .A2(n_3461),
    .B1(\u8_mem[0] [31]),
    .B2(n_3460),
    .Y(n_10352));
 AOI22xp5_ASAP7_75t_SL g165993 (.A1(n_3320),
    .A2(n_22640),
    .B1(\u8_mem[2] [28]),
    .B2(n_16900),
    .Y(n_10363));
 AOI22xp5_ASAP7_75t_SL g165996 (.A1(n_3420),
    .A2(n_65920),
    .B1(\u6_mem[0] [28]),
    .B2(n_3425),
    .Y(n_10366));
 AOI22xp5_ASAP7_75t_SL g165999 (.A1(n_22640),
    .A2(n_73997),
    .B1(\u8_mem[1] [28]),
    .B2(n_31460),
    .Y(n_10369));
 INVxp33_ASAP7_75t_R g166 (.A(wb_data_i[9]),
    .Y(n_65992));
 AOI22xp5_ASAP7_75t_SL g166000 (.A1(n_65920),
    .A2(n_32163),
    .B1(\u5_mem[1] [28]),
    .B2(n_13508),
    .Y(n_10370));
 AOI22xp5_ASAP7_75t_SL g166002 (.A1(n_22640),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [28]),
    .Y(n_10372));
 AOI22xp5_ASAP7_75t_SL g166006 (.A1(n_3285),
    .A2(n_65920),
    .B1(\u5_mem[2] [28]),
    .B2(n_43020),
    .Y(n_10376));
 AOI22xp5_ASAP7_75t_SL g166007 (.A1(n_3188),
    .A2(n_22640),
    .B1(\u7_mem[2] [28]),
    .B2(n_13333),
    .Y(n_10377));
 AOI22xp33_ASAP7_75t_SL g166008 (.A1(n_24633),
    .A2(n_65920),
    .B1(\u4_mem[2] [28]),
    .B2(n_13304),
    .Y(n_10378));
 AOI22xp5_ASAP7_75t_SL g166009 (.A1(n_22640),
    .A2(n_3461),
    .B1(\u8_mem[0] [28]),
    .B2(n_3453),
    .Y(n_10379));
 AOI22xp5_ASAP7_75t_SL g166042 (.A1(n_3320),
    .A2(n_65915),
    .B1(\u8_mem[2] [24]),
    .B2(n_16900),
    .Y(n_10413));
 AOI22xp5_ASAP7_75t_SL g166043 (.A1(n_3420),
    .A2(n_65915),
    .B1(\u6_mem[0] [24]),
    .B2(n_3415),
    .Y(n_10414));
 AOI22xp5_ASAP7_75t_SL g166049 (.A1(n_65917),
    .A2(n_32163),
    .B1(\u5_mem[1] [24]),
    .B2(n_13500),
    .Y(n_10420));
 AOI22xp5_ASAP7_75t_SL g166051 (.A1(n_65917),
    .A2(n_14386),
    .B1(n_31741),
    .B2(\u6_mem[1] [24]),
    .Y(n_10422));
 AOI22xp5_ASAP7_75t_SL g166055 (.A1(n_3285),
    .A2(n_65915),
    .B1(\u5_mem[2] [24]),
    .B2(n_43020),
    .Y(n_10426));
 AOI22xp5_ASAP7_75t_SL g166058 (.A1(n_3188),
    .A2(n_28424),
    .B1(\u7_mem[2] [24]),
    .B2(n_13325),
    .Y(n_10429));
 AOI22xp5_ASAP7_75t_SL g166059 (.A1(n_24633),
    .A2(n_65914),
    .B1(\u4_mem[2] [24]),
    .B2(n_13304),
    .Y(n_10430));
 AOI22xp5_ASAP7_75t_SL g166060 (.A1(n_28424),
    .A2(n_3461),
    .B1(\u8_mem[0] [24]),
    .B2(n_3460),
    .Y(n_10431));
 AOI22xp33_ASAP7_75t_SL g166068 (.A1(n_3320),
    .A2(n_65924),
    .B1(\u8_mem[2] [25]),
    .B2(n_16900),
    .Y(n_10439));
 AOI22xp5_ASAP7_75t_SL g166071 (.A1(n_3420),
    .A2(n_65925),
    .B1(\u6_mem[0] [25]),
    .B2(n_3415),
    .Y(n_10442));
 AOI22xp5_ASAP7_75t_SL g166075 (.A1(n_65927),
    .A2(n_32164),
    .B1(\u5_mem[1] [25]),
    .B2(n_13508),
    .Y(n_10446));
 AOI22xp5_ASAP7_75t_SL g166081 (.A1(n_3285),
    .A2(n_65924),
    .B1(\u5_mem[2] [25]),
    .B2(n_43028),
    .Y(n_10452));
 AOI22xp33_ASAP7_75t_SL g166084 (.A1(n_3188),
    .A2(n_28316),
    .B1(\u7_mem[2] [25]),
    .B2(n_13333),
    .Y(n_10455));
 AOI22xp5_ASAP7_75t_SL g166085 (.A1(n_24633),
    .A2(n_65925),
    .B1(\u4_mem[2] [25]),
    .B2(n_13304),
    .Y(n_10456));
 AOI22xp5_ASAP7_75t_SL g166086 (.A1(n_28316),
    .A2(n_3454),
    .B1(\u8_mem[0] [25]),
    .B2(n_3460),
    .Y(n_10457));
 AOI22xp5_ASAP7_75t_SL g166092 (.A1(n_3320),
    .A2(n_35437),
    .B1(\u8_mem[2] [26]),
    .B2(n_16900),
    .Y(n_10464));
 AOI22xp5_ASAP7_75t_SL g166096 (.A1(n_3420),
    .A2(n_66010),
    .B1(\u6_mem[0] [26]),
    .B2(n_3425),
    .Y(n_10467));
 AOI22xp5_ASAP7_75t_SL g166099 (.A1(n_35437),
    .A2(n_73997),
    .B1(\u8_mem[1] [26]),
    .B2(n_31464),
    .Y(n_10470));
 AOI22xp5_ASAP7_75t_SL g166100 (.A1(n_66011),
    .A2(n_32163),
    .B1(\u5_mem[1] [26]),
    .B2(n_13508),
    .Y(n_10471));
 AOI22xp5_ASAP7_75t_SL g166102 (.A1(n_66010),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [26]),
    .Y(n_10473));
 AOI22xp5_ASAP7_75t_SL g166106 (.A1(n_3285),
    .A2(n_66011),
    .B1(\u5_mem[2] [26]),
    .B2(n_43020),
    .Y(n_10477));
 AOI22xp5_ASAP7_75t_SL g166110 (.A1(n_3188),
    .A2(n_66011),
    .B1(\u7_mem[2] [26]),
    .B2(n_13325),
    .Y(n_10481));
 AOI22xp5_ASAP7_75t_SL g166111 (.A1(n_24633),
    .A2(n_35437),
    .B1(\u4_mem[2] [26]),
    .B2(n_13304),
    .Y(n_10482));
 AOI22xp5_ASAP7_75t_SL g166112 (.A1(n_66010),
    .A2(n_3454),
    .B1(\u8_mem[0] [26]),
    .B2(n_3460),
    .Y(n_10483));
 AOI22xp5_ASAP7_75t_SL g166118 (.A1(n_3320),
    .A2(n_62940),
    .B1(\u8_mem[2] [27]),
    .B2(n_16900),
    .Y(n_10490));
 AOI22xp5_ASAP7_75t_SL g166122 (.A1(n_3420),
    .A2(n_65910),
    .B1(\u6_mem[0] [27]),
    .B2(n_3425),
    .Y(n_10493));
 AOI22xp5_ASAP7_75t_SL g166125 (.A1(n_62940),
    .A2(n_73997),
    .B1(\u8_mem[1] [27]),
    .B2(n_73399),
    .Y(n_10496));
 AOI22xp5_ASAP7_75t_SL g166126 (.A1(n_65910),
    .A2(n_32163),
    .B1(\u5_mem[1] [27]),
    .B2(n_13500),
    .Y(n_10497));
 AOI22xp5_ASAP7_75t_SL g166128 (.A1(n_65908),
    .A2(n_14386),
    .B1(n_31741),
    .B2(\u6_mem[1] [27]),
    .Y(n_10499));
 AOI22xp5_ASAP7_75t_SL g166132 (.A1(n_3285),
    .A2(n_65908),
    .B1(\u5_mem[2] [27]),
    .B2(n_43028),
    .Y(n_10503));
 AOI22xp5_ASAP7_75t_SL g166135 (.A1(n_3188),
    .A2(n_62940),
    .B1(\u7_mem[2] [27]),
    .B2(n_13333),
    .Y(n_10506));
 AOI22xp5_ASAP7_75t_SL g166136 (.A1(n_24633),
    .A2(n_65908),
    .B1(\u4_mem[2] [27]),
    .B2(n_13304),
    .Y(n_10507));
 AOI22xp5_ASAP7_75t_SL g166138 (.A1(n_65908),
    .A2(n_3454),
    .B1(\u8_mem[0] [27]),
    .B2(n_3460),
    .Y(n_10509));
 INVx1_ASAP7_75t_SL g166190 (.A(n_28895),
    .Y(n_10565));
 NAND2x1p5_ASAP7_75t_L g166192 (.A(wb_addr_i[3]),
    .B(wb_addr_i[2]),
    .Y(n_10563));
 OR2x6_ASAP7_75t_SL g166238 (.A(n_8313),
    .B(n_8315),
    .Y(n_10613));
 AOI21xp33_ASAP7_75t_SL g166239 (.A1(n_2678),
    .A2(n_10614),
    .B(n_31821),
    .Y(n_10615));
 INVx4_ASAP7_75t_SL g166240 (.A(n_10613),
    .Y(n_10614));
 AOI21xp33_ASAP7_75t_SL g166242 (.A1(n_10614),
    .A2(n_2079),
    .B(n_11003),
    .Y(n_10617));
 AOI21xp5_ASAP7_75t_SL g166245 (.A1(n_2106),
    .A2(n_10614),
    .B(n_11010),
    .Y(n_10620));
 AOI22xp5_ASAP7_75t_L g166246 (.A1(n_14933),
    .A2(i6_dout[24]),
    .B1(n_10614),
    .B2(n_2024),
    .Y(n_10621));
 AOI21xp5_ASAP7_75t_SL g166247 (.A1(n_10614),
    .A2(n_2063),
    .B(n_10873),
    .Y(n_10622));
 AOI21xp33_ASAP7_75t_SL g166248 (.A1(n_10614),
    .A2(u13_ints_r[7]),
    .B(n_11013),
    .Y(n_10623));
 AOI21xp33_ASAP7_75t_SL g166249 (.A1(n_10614),
    .A2(u13_ints_r[12]),
    .B(n_11009),
    .Y(n_10624));
 AOI21xp33_ASAP7_75t_SL g166251 (.A1(n_10626),
    .A2(u13_ints_r[13]),
    .B(n_11007),
    .Y(n_10627));
 AOI21xp5_ASAP7_75t_SL g166252 (.A1(u13_ints_r[17]),
    .A2(n_10626),
    .B(n_10885),
    .Y(n_10628));
 AOI21xp5_ASAP7_75t_SL g166253 (.A1(n_10626),
    .A2(n_2065),
    .B(n_11004),
    .Y(n_10629));
 AOI21xp5_ASAP7_75t_SL g166255 (.A1(n_10626),
    .A2(n_2031),
    .B(n_11008),
    .Y(n_10631));
 AOI21xp5_ASAP7_75t_SL g166257 (.A1(n_10626),
    .A2(n_2036),
    .B(n_11017),
    .Y(n_10633));
 AOI21xp5_ASAP7_75t_SL g166259 (.A1(n_10626),
    .A2(n_2034),
    .B(n_26579),
    .Y(n_10635));
 AOI21xp5_ASAP7_75t_L g166260 (.A1(n_10626),
    .A2(n_2130),
    .B(n_11019),
    .Y(n_10636));
 AOI22xp5_ASAP7_75t_SL g166262 (.A1(n_3285),
    .A2(n_10640),
    .B1(\u5_mem[2] [30]),
    .B2(n_43020),
    .Y(n_10641));
 AOI22xp5_ASAP7_75t_SL g166263 (.A1(n_3320),
    .A2(n_10638),
    .B1(\u8_mem[2] [30]),
    .B2(n_16900),
    .Y(n_10642));
 AOI22xp5_ASAP7_75t_SL g166265 (.A1(n_3461),
    .A2(n_10638),
    .B1(\u8_mem[0] [30]),
    .B2(n_3453),
    .Y(n_10644));
 AOI22xp5_ASAP7_75t_SL g166270 (.A1(n_3420),
    .A2(n_10640),
    .B1(\u6_mem[0] [30]),
    .B2(n_3415),
    .Y(n_10649));
 AOI22xp5_ASAP7_75t_SL g166272 (.A1(n_32163),
    .A2(n_10640),
    .B1(\u5_mem[1] [30]),
    .B2(n_13500),
    .Y(n_10651));
 AOI22xp5_ASAP7_75t_SL g166275 (.A1(n_10638),
    .A2(n_14386),
    .B1(n_22396),
    .B2(\u6_mem[1] [30]),
    .Y(n_10654));
 AOI22xp5_ASAP7_75t_SL g166277 (.A1(n_3188),
    .A2(n_10638),
    .B1(\u7_mem[2] [30]),
    .B2(n_13325),
    .Y(n_10656));
 AOI22xp5_ASAP7_75t_SL g166278 (.A1(n_24633),
    .A2(n_10640),
    .B1(\u4_mem[2] [30]),
    .B2(n_13304),
    .Y(n_10657));
 HB1xp67_ASAP7_75t_R g166280 (.A(wb_din[30]),
    .Y(n_10659));
 HB1xp67_ASAP7_75t_SL g166281 (.A(wb_din[30]),
    .Y(n_10660));
 AOI22xp5_ASAP7_75t_SL g166285 (.A1(n_3461),
    .A2(n_22715),
    .B1(\u8_mem[0] [29]),
    .B2(n_3453),
    .Y(n_10665));
 AOI22xp5_ASAP7_75t_SL g166287 (.A1(n_3320),
    .A2(n_15952),
    .B1(\u8_mem[2] [29]),
    .B2(n_16900),
    .Y(n_10666));
 AOI22xp5_ASAP7_75t_SL g166290 (.A1(n_3420),
    .A2(n_22715),
    .B1(\u6_mem[0] [29]),
    .B2(n_3425),
    .Y(n_10669));
 AOI22xp5_ASAP7_75t_SL g166291 (.A1(n_32163),
    .A2(n_15952),
    .B1(\u5_mem[1] [29]),
    .B2(n_13508),
    .Y(n_10670));
 AOI22xp5_ASAP7_75t_SL g166297 (.A1(n_15952),
    .A2(n_14386),
    .B1(n_31741),
    .B2(\u6_mem[1] [29]),
    .Y(n_10676));
 AOI22xp5_ASAP7_75t_SL g166300 (.A1(n_3285),
    .A2(n_22715),
    .B1(\u5_mem[2] [29]),
    .B2(n_43020),
    .Y(n_10679));
 AOI22xp5_ASAP7_75t_SL g166301 (.A1(n_3188),
    .A2(n_15952),
    .B1(\u7_mem[2] [29]),
    .B2(n_13333),
    .Y(n_10680));
 AOI22xp5_ASAP7_75t_SL g166302 (.A1(n_24633),
    .A2(n_22715),
    .B1(\u4_mem[2] [29]),
    .B2(n_13304),
    .Y(n_10681));
 HB1xp67_ASAP7_75t_R g166304 (.A(wb_din[29]),
    .Y(n_10683));
 HB1xp67_ASAP7_75t_SL g166305 (.A(wb_din[29]),
    .Y(n_10684));
 NOR3x2_ASAP7_75t_SL g166481 (.B(wb_addr_i[3]),
    .C(wb_addr_i[2]),
    .Y(n_10867),
    .A(n_8296));
 OAI22xp5_ASAP7_75t_SL g166482 (.A1(n_1319),
    .A2(n_14909),
    .B1(n_263),
    .B2(n_10576),
    .Y(n_10869));
 OAI22xp33_ASAP7_75t_SL g166484 (.A1(n_1325),
    .A2(n_14909),
    .B1(n_166),
    .B2(n_10576),
    .Y(n_10870));
 OAI22xp5_ASAP7_75t_SL g166485 (.A1(n_76),
    .A2(n_14909),
    .B1(n_28669),
    .B2(n_57),
    .Y(n_10871));
 OAI22xp5_ASAP7_75t_SL g166487 (.A1(n_157),
    .A2(n_14909),
    .B1(n_10576),
    .B2(n_27003),
    .Y(n_10873));
 OAI22xp5_ASAP7_75t_SL g166491 (.A1(n_152),
    .A2(n_14909),
    .B1(n_97),
    .B2(n_6960),
    .Y(n_10877));
 OAI22xp33_ASAP7_75t_SL g166492 (.A1(n_95),
    .A2(n_14909),
    .B1(n_608),
    .B2(n_6960),
    .Y(n_10878));
 OAI22xp5_ASAP7_75t_SL g166494 (.A1(n_65),
    .A2(n_10889),
    .B1(n_6960),
    .B2(n_34532),
    .Y(n_10881));
 OAI22xp5_ASAP7_75t_SL g166495 (.A1(n_158),
    .A2(n_10889),
    .B1(n_28669),
    .B2(n_18900),
    .Y(n_10882));
 OAI22xp33_ASAP7_75t_SL g166497 (.A1(n_49),
    .A2(n_10889),
    .B1(n_6960),
    .B2(n_257),
    .Y(n_10884));
 OAI22xp5_ASAP7_75t_SL g166498 (.A1(n_1322),
    .A2(n_10889),
    .B1(n_10576),
    .B2(n_2640),
    .Y(n_10885));
 OAI22xp5_ASAP7_75t_SL g166500 (.A1(n_153),
    .A2(n_10889),
    .B1(n_41),
    .B2(n_6960),
    .Y(n_10887));
 OAI22xp33_ASAP7_75t_SL g166501 (.A1(n_99),
    .A2(n_10889),
    .B1(n_201),
    .B2(n_6960),
    .Y(n_10888));
 AOI22xp5_ASAP7_75t_SL g166503 (.A1(n_3320),
    .A2(n_10891),
    .B1(\u8_mem[2] [1]),
    .B2(n_16908),
    .Y(n_10892));
 AOI22xp5_ASAP7_75t_SL g166504 (.A1(n_3285),
    .A2(n_78044),
    .B1(\u5_mem[2] [1]),
    .B2(n_43020),
    .Y(n_10894));
 AOI22xp5_ASAP7_75t_SL g166505 (.A1(n_3188),
    .A2(n_78044),
    .B1(\u7_mem[2] [1]),
    .B2(n_13333),
    .Y(n_10895));
 AOI22xp5_ASAP7_75t_SL g166506 (.A1(n_24633),
    .A2(n_10891),
    .B1(\u4_mem[2] [1]),
    .B2(n_13312),
    .Y(n_10896));
 AOI22xp5_ASAP7_75t_SL g166512 (.A1(n_3420),
    .A2(n_10891),
    .B1(\u6_mem[0] [1]),
    .B2(n_3425),
    .Y(n_10902));
 AOI22xp5_ASAP7_75t_SL g166516 (.A1(n_10891),
    .A2(n_3454),
    .B1(\u8_mem[0] [1]),
    .B2(n_3453),
    .Y(n_10906));
 NAND3xp33_ASAP7_75t_L g166520 (.A(rf_we),
    .B(n_78044),
    .C(n_7196),
    .Y(n_10910));
 BUFx2_ASAP7_75t_L g166522 (.A(wb_din[1]),
    .Y(n_3815));
 NAND3xp33_ASAP7_75t_R g166526 (.A(n_75733),
    .B(rf_we),
    .C(n_7196),
    .Y(n_10916));
 AOI22xp5_ASAP7_75t_SL g166528 (.A1(n_24633),
    .A2(n_33203),
    .B1(\u4_mem[2] [0]),
    .B2(n_13304),
    .Y(n_10918));
 AOI22xp5_ASAP7_75t_SL g166529 (.A1(n_3188),
    .A2(n_33203),
    .B1(\u7_mem[2] [0]),
    .B2(n_13333),
    .Y(n_10919));
 AOI22xp5_ASAP7_75t_SL g166531 (.A1(n_3285),
    .A2(n_33203),
    .B1(\u5_mem[2] [0]),
    .B2(n_43020),
    .Y(n_10921));
 AOI22xp5_ASAP7_75t_SL g166532 (.A1(n_3320),
    .A2(n_75733),
    .B1(\u8_mem[2] [0]),
    .B2(n_16908),
    .Y(n_10922));
 AOI22xp5_ASAP7_75t_SL g166533 (.A1(n_75733),
    .A2(n_3454),
    .B1(\u8_mem[0] [0]),
    .B2(n_3453),
    .Y(n_10923));
 AOI22xp5_ASAP7_75t_SL g166538 (.A1(n_3420),
    .A2(n_10924),
    .B1(\u6_mem[0] [0]),
    .B2(n_3425),
    .Y(n_10929));
 NAND4xp25_ASAP7_75t_SL g166544 (.A(n_10935),
    .B(n_28955),
    .C(n_1059),
    .D(n_27257),
    .Y(n_10936));
 BUFx6f_ASAP7_75t_SL g166545 (.A(n_20426),
    .Y(n_10935));
 INVx5_ASAP7_75t_SL g166546 (.A(n_10935),
    .Y(n_10937));
 NAND2xp5_ASAP7_75t_L g166550 (.A(u11_din_tmp1[7]),
    .B(n_10935),
    .Y(n_10941));
 NAND2xp5_ASAP7_75t_SL g166551 (.A(u11_din_tmp1[6]),
    .B(n_10935),
    .Y(n_10942));
 NAND2xp5_ASAP7_75t_L g166552 (.A(u11_din_tmp1[11]),
    .B(n_10935),
    .Y(n_10943));
 NAND2xp5_ASAP7_75t_L g166553 (.A(u11_din_tmp1[15]),
    .B(n_10935),
    .Y(n_10944));
 AOI22xp5_ASAP7_75t_SL g166567 (.A1(n_21311),
    .A2(n_10891),
    .B1(oc4_cfg[1]),
    .B2(n_26541),
    .Y(n_10959));
 AOI22xp5_ASAP7_75t_SL g166568 (.A1(n_35041),
    .A2(n_21311),
    .B1(oc5_cfg[5]),
    .B2(n_26541),
    .Y(n_10960));
 AOI22xp5_ASAP7_75t_SL g166569 (.A1(n_66868),
    .A2(n_21311),
    .B1(oc4_cfg[5]),
    .B2(n_26541),
    .Y(n_10961));
 AOI22xp5_ASAP7_75t_SL g166570 (.A1(n_10026),
    .A2(n_21311),
    .B1(n_294),
    .B2(n_26541),
    .Y(n_10962));
 AOI22xp5_ASAP7_75t_SL g166571 (.A1(n_66842),
    .A2(n_21311),
    .B1(n_79193),
    .B2(n_26541),
    .Y(n_10963));
 AOI22xp5_ASAP7_75t_SL g166576 (.A1(n_66855),
    .A2(n_15272),
    .B1(n_50293),
    .B2(n_26541),
    .Y(n_10969));
 AOI22xp5_ASAP7_75t_SL g166577 (.A1(n_28330),
    .A2(n_15272),
    .B1(n_247),
    .B2(n_26541),
    .Y(n_10970));
 AOI22xp5_ASAP7_75t_SL g166578 (.A1(n_65969),
    .A2(n_15272),
    .B1(u13_occ1_r[7]),
    .B2(n_26541),
    .Y(n_10971));
 NAND2x1_ASAP7_75t_SL g166608 (.A(wb_addr_i[3]),
    .B(n_8238),
    .Y(n_11000));
 OAI22xp33_ASAP7_75t_SL g166609 (.A1(n_101),
    .A2(n_11011),
    .B1(n_264),
    .B2(n_28895),
    .Y(n_11003));
 OAI22xp5_ASAP7_75t_SL g166610 (.A1(n_11011),
    .A2(n_79192),
    .B1(n_10889),
    .B2(n_130),
    .Y(n_11004));
 OAI22xp5_ASAP7_75t_SL g166613 (.A1(n_11011),
    .A2(n_59),
    .B1(n_10576),
    .B2(n_1379),
    .Y(n_11007));
 OAI22xp33_ASAP7_75t_SL g166614 (.A1(n_35656),
    .A2(n_11011),
    .B1(n_10576),
    .B2(n_2645),
    .Y(n_11008));
 OAI22xp33_ASAP7_75t_SL g166615 (.A1(n_11011),
    .A2(n_293),
    .B1(n_28895),
    .B2(n_1501),
    .Y(n_11009));
 OAI22xp5_ASAP7_75t_SL g166616 (.A1(n_11011),
    .A2(n_103),
    .B1(n_28895),
    .B2(n_1503),
    .Y(n_11010));
 OAI22xp5_ASAP7_75t_SL g166617 (.A1(n_11011),
    .A2(n_70326),
    .B1(n_28895),
    .B2(n_8186),
    .Y(n_11012));
 OAI22xp5_ASAP7_75t_SL g166618 (.A1(n_11011),
    .A2(n_133),
    .B1(n_28895),
    .B2(n_1496),
    .Y(n_11013));
 OAI22xp5_ASAP7_75t_L g166620 (.A1(n_11011),
    .A2(n_81),
    .B1(n_10576),
    .B2(n_1494),
    .Y(n_11015));
 OAI22xp5_ASAP7_75t_SL g166622 (.A1(n_11011),
    .A2(n_229),
    .B1(n_10576),
    .B2(n_1376),
    .Y(n_11017));
 OAI22xp5_ASAP7_75t_SL g166624 (.A1(n_11011),
    .A2(n_1381),
    .B1(n_28895),
    .B2(n_25293),
    .Y(n_11019));
 INVx2_ASAP7_75t_SL g166696 (.A(u11_wp[2]),
    .Y(n_225));
 BUFx2_ASAP7_75t_SL g166713 (.A(n_26382),
    .Y(n_11124));
 AOI22xp5_ASAP7_75t_SL g166714 (.A1(n_11126),
    .A2(n_65952),
    .B1(\u5_mem[3] [17]),
    .B2(n_11125),
    .Y(n_11127));
 INVx5_ASAP7_75t_SL g166715 (.A(n_11125),
    .Y(n_11126));
 AOI22xp5_ASAP7_75t_SL g166717 (.A1(n_11128),
    .A2(n_65949),
    .B1(\u5_mem[3] [16]),
    .B2(n_11125),
    .Y(n_11129));
 AOI31xp33_ASAP7_75t_SL g166719 (.A1(n_11125),
    .A2(u5_wp[2]),
    .A3(n_35577),
    .B(n_35578),
    .Y(n_11130));
 AOI22xp33_ASAP7_75t_SL g166720 (.A1(n_11126),
    .A2(n_65902),
    .B1(\u5_mem[3] [31]),
    .B2(n_11125),
    .Y(n_11131));
 AOI22xp5_ASAP7_75t_SL g166721 (.A1(n_11128),
    .A2(n_10660),
    .B1(\u5_mem[3] [30]),
    .B2(n_11125),
    .Y(n_11132));
 AOI22xp5_ASAP7_75t_SL g166722 (.A1(n_11126),
    .A2(n_10684),
    .B1(\u5_mem[3] [29]),
    .B2(n_11125),
    .Y(n_11133));
 AOI22xp5_ASAP7_75t_SL g166723 (.A1(n_11128),
    .A2(n_65920),
    .B1(\u5_mem[3] [28]),
    .B2(n_11125),
    .Y(n_11134));
 AOI22xp5_ASAP7_75t_SL g166724 (.A1(n_11128),
    .A2(n_66010),
    .B1(\u5_mem[3] [26]),
    .B2(n_11135),
    .Y(n_11136));
 AOI22xp5_ASAP7_75t_SL g166725 (.A1(n_11126),
    .A2(n_65925),
    .B1(\u5_mem[3] [25]),
    .B2(n_11135),
    .Y(n_11137));
 AOI22xp5_ASAP7_75t_SL g166726 (.A1(n_11128),
    .A2(n_65915),
    .B1(\u5_mem[3] [24]),
    .B2(n_11135),
    .Y(n_11138));
 AOI22xp5_ASAP7_75t_SL g166727 (.A1(n_11128),
    .A2(n_10329),
    .B1(\u5_mem[3] [23]),
    .B2(n_11135),
    .Y(n_11139));
 AOI22xp5_ASAP7_75t_SL g166728 (.A1(n_11126),
    .A2(n_65941),
    .B1(\u5_mem[3] [22]),
    .B2(n_11135),
    .Y(n_11140));
 AOI22xp5_ASAP7_75t_SL g166729 (.A1(n_11126),
    .A2(n_66016),
    .B1(\u5_mem[3] [21]),
    .B2(n_11135),
    .Y(n_11141));
 AOI22xp5_ASAP7_75t_SL g166730 (.A1(n_11126),
    .A2(n_10247),
    .B1(\u5_mem[3] [20]),
    .B2(n_11135),
    .Y(n_11142));
 AOI22xp33_ASAP7_75t_SL g166731 (.A1(n_11128),
    .A2(n_65932),
    .B1(\u5_mem[3] [19]),
    .B2(n_11135),
    .Y(n_11143));
 AOI22xp5_ASAP7_75t_SL g166732 (.A1(n_11128),
    .A2(n_10194),
    .B1(\u5_mem[3] [18]),
    .B2(n_11135),
    .Y(n_11144));
 AOI22xp5_ASAP7_75t_SL g166769 (.A1(n_47390),
    .A2(n_66010),
    .B1(\u4_mem[3] [26]),
    .B2(n_35909),
    .Y(n_11183));
 AOI22xp5_ASAP7_75t_SL g166770 (.A1(n_47390),
    .A2(n_65925),
    .B1(\u4_mem[3] [25]),
    .B2(n_35909),
    .Y(n_11184));
 AOI22xp5_ASAP7_75t_SL g166771 (.A1(n_30253),
    .A2(n_65915),
    .B1(\u4_mem[3] [24]),
    .B2(n_35909),
    .Y(n_11185));
 AOI22xp5_ASAP7_75t_SL g166772 (.A1(n_30253),
    .A2(n_10329),
    .B1(\u4_mem[3] [23]),
    .B2(n_35909),
    .Y(n_11186));
 AOI22xp5_ASAP7_75t_SL g166773 (.A1(n_30253),
    .A2(n_10302),
    .B1(\u4_mem[3] [22]),
    .B2(n_35909),
    .Y(n_11187));
 AOI22xp33_ASAP7_75t_SL g166774 (.A1(n_47390),
    .A2(n_32916),
    .B1(\u4_mem[3] [21]),
    .B2(n_35909),
    .Y(n_11188));
 AOI22xp33_ASAP7_75t_SL g166776 (.A1(n_47390),
    .A2(n_65932),
    .B1(\u4_mem[3] [19]),
    .B2(n_35909),
    .Y(n_11190));
 AOI22xp33_ASAP7_75t_SL g166777 (.A1(n_30253),
    .A2(n_10194),
    .B1(\u4_mem[3] [18]),
    .B2(n_35909),
    .Y(n_11191));
 AOI22xp33_ASAP7_75t_SL g166783 (.A1(n_65952),
    .A2(n_64819),
    .B1(\u8_mem[3] [17]),
    .B2(n_72908),
    .Y(n_11197));
 AOI22xp33_ASAP7_75t_SL g166797 (.A1(n_64818),
    .A2(n_65932),
    .B1(\u8_mem[3] [19]),
    .B2(n_11204),
    .Y(n_11212));
 AOI22xp33_ASAP7_75t_SL g166841 (.A1(n_66856),
    .A2(n_14570),
    .B1(\u7_mem[3] [3]),
    .B2(n_33777),
    .Y(n_11259));
 AOI22xp5_ASAP7_75t_SL g166878 (.A1(n_3815),
    .A2(n_61228),
    .B1(\u6_mem[3] [1]),
    .B2(n_77233),
    .Y(n_11295));
 INVx1_ASAP7_75t_SL g166892 (.A(n_225),
    .Y(n_11312));
 INVxp33_ASAP7_75t_R g167 (.A(wb_data_i[12]),
    .Y(n_65995));
 AOI321xp33_ASAP7_75t_SL g167023 (.A1(n_1167),
    .A2(n_2788),
    .A3(i6_re),
    .B1(n_11477),
    .B2(n_2788),
    .C(n_2453),
    .Y(n_11478));
 AND2x6_ASAP7_75t_SL g167024 (.A(u11_rp[1]),
    .B(n_13027),
    .Y(n_11477));
 AOI321xp33_ASAP7_75t_SL g167058 (.A1(n_1171),
    .A2(n_375),
    .A3(i3_re),
    .B1(n_11512),
    .B2(n_375),
    .C(n_2452),
    .Y(n_11513));
 AND2x6_ASAP7_75t_SL g167059 (.A(u9_rp[1]),
    .B(n_13035),
    .Y(n_11512));
 AND2x6_ASAP7_75t_SL g167095 (.A(n_13761),
    .B(n_25439),
    .Y(n_11548));
 AOI22xp5_ASAP7_75t_SL g167096 (.A1(n_11548),
    .A2(\u10_mem[0] [11]),
    .B1(n_14825),
    .B2(\u10_mem[1] [11]),
    .Y(n_11550));
 AOI22xp5_ASAP7_75t_SL g167097 (.A1(n_11548),
    .A2(\u10_mem[0] [8]),
    .B1(n_14825),
    .B2(\u10_mem[1] [8]),
    .Y(n_11551));
 AOI22xp5_ASAP7_75t_SL g167098 (.A1(n_11548),
    .A2(\u10_mem[0] [10]),
    .B1(n_14825),
    .B2(\u10_mem[1] [10]),
    .Y(n_11552));
 AOI22xp5_ASAP7_75t_SL g167099 (.A1(n_11548),
    .A2(\u10_mem[0] [22]),
    .B1(n_14825),
    .B2(\u10_mem[1] [22]),
    .Y(n_11553));
 AOI22xp5_ASAP7_75t_SL g167100 (.A1(n_11548),
    .A2(\u10_mem[0] [28]),
    .B1(n_14825),
    .B2(\u10_mem[1] [28]),
    .Y(n_11554));
 AOI22xp5_ASAP7_75t_SL g167101 (.A1(n_11548),
    .A2(\u10_mem[0] [3]),
    .B1(n_14825),
    .B2(\u10_mem[1] [3]),
    .Y(n_11555));
 AOI22xp5_ASAP7_75t_SL g167102 (.A1(n_11548),
    .A2(\u10_mem[0] [31]),
    .B1(n_14825),
    .B2(\u10_mem[1] [31]),
    .Y(n_11556));
 AOI22xp5_ASAP7_75t_SL g167103 (.A1(n_11548),
    .A2(\u10_mem[0] [4]),
    .B1(n_14825),
    .B2(\u10_mem[1] [4]),
    .Y(n_11557));
 AOI22xp5_ASAP7_75t_SL g167104 (.A1(n_11548),
    .A2(\u10_mem[0] [27]),
    .B1(n_14825),
    .B2(\u10_mem[1] [27]),
    .Y(n_11558));
 AOI22xp5_ASAP7_75t_SL g167105 (.A1(n_11548),
    .A2(\u10_mem[0] [7]),
    .B1(n_14825),
    .B2(\u10_mem[1] [7]),
    .Y(n_11559));
 AOI22xp5_ASAP7_75t_SL g167106 (.A1(n_11548),
    .A2(\u10_mem[0] [30]),
    .B1(n_14825),
    .B2(\u10_mem[1] [30]),
    .Y(n_11560));
 AOI22xp5_ASAP7_75t_SL g167107 (.A1(n_11548),
    .A2(\u10_mem[0] [25]),
    .B1(n_14825),
    .B2(\u10_mem[1] [25]),
    .Y(n_11561));
 AOI22xp5_ASAP7_75t_SL g167108 (.A1(n_11548),
    .A2(\u10_mem[0] [24]),
    .B1(n_14825),
    .B2(\u10_mem[1] [24]),
    .Y(n_11562));
 AOI22xp5_ASAP7_75t_SL g167109 (.A1(n_11548),
    .A2(\u10_mem[0] [18]),
    .B1(n_14825),
    .B2(\u10_mem[1] [18]),
    .Y(n_11563));
 AOI22xp5_ASAP7_75t_SL g167110 (.A1(n_11548),
    .A2(\u10_mem[0] [2]),
    .B1(n_14825),
    .B2(\u10_mem[1] [2]),
    .Y(n_11564));
 AOI22xp5_ASAP7_75t_SL g167111 (.A1(n_11548),
    .A2(\u10_mem[0] [6]),
    .B1(n_14825),
    .B2(\u10_mem[1] [6]),
    .Y(n_11565));
 AOI22xp5_ASAP7_75t_SL g167112 (.A1(n_11548),
    .A2(\u10_mem[0] [12]),
    .B1(n_14825),
    .B2(\u10_mem[1] [12]),
    .Y(n_11566));
 AOI22xp5_ASAP7_75t_SL g167113 (.A1(n_11548),
    .A2(\u10_mem[0] [29]),
    .B1(n_14825),
    .B2(\u10_mem[1] [29]),
    .Y(n_11567));
 AOI22xp5_ASAP7_75t_SL g167114 (.A1(n_11548),
    .A2(\u10_mem[0] [17]),
    .B1(n_14825),
    .B2(\u10_mem[1] [17]),
    .Y(n_11568));
 AOI22xp5_ASAP7_75t_SL g167115 (.A1(n_11548),
    .A2(\u10_mem[0] [20]),
    .B1(n_14825),
    .B2(\u10_mem[1] [20]),
    .Y(n_11569));
 AOI22xp5_ASAP7_75t_SL g167116 (.A1(n_11548),
    .A2(\u10_mem[0] [1]),
    .B1(n_14825),
    .B2(\u10_mem[1] [1]),
    .Y(n_11570));
 AOI22xp5_ASAP7_75t_SL g167117 (.A1(n_11548),
    .A2(\u10_mem[0] [13]),
    .B1(n_14825),
    .B2(\u10_mem[1] [13]),
    .Y(n_11571));
 AOI22xp5_ASAP7_75t_SL g167118 (.A1(n_11548),
    .A2(\u10_mem[0] [26]),
    .B1(n_14825),
    .B2(\u10_mem[1] [26]),
    .Y(n_11572));
 AOI22xp5_ASAP7_75t_SL g167119 (.A1(n_11548),
    .A2(\u10_mem[0] [21]),
    .B1(n_14825),
    .B2(\u10_mem[1] [21]),
    .Y(n_11573));
 AOI22xp5_ASAP7_75t_SL g167120 (.A1(n_11548),
    .A2(\u10_mem[0] [19]),
    .B1(n_14825),
    .B2(\u10_mem[1] [19]),
    .Y(n_11574));
 AOI22xp5_ASAP7_75t_SL g167121 (.A1(n_11548),
    .A2(\u10_mem[0] [14]),
    .B1(n_14825),
    .B2(\u10_mem[1] [14]),
    .Y(n_11575));
 AOI22xp5_ASAP7_75t_SL g167122 (.A1(n_11548),
    .A2(\u10_mem[0] [0]),
    .B1(n_14825),
    .B2(\u10_mem[1] [0]),
    .Y(n_11576));
 AOI22xp5_ASAP7_75t_SL g167123 (.A1(n_11548),
    .A2(\u10_mem[0] [16]),
    .B1(n_14825),
    .B2(\u10_mem[1] [16]),
    .Y(n_11577));
 AOI22xp5_ASAP7_75t_SL g167124 (.A1(n_11548),
    .A2(\u10_mem[0] [15]),
    .B1(n_14825),
    .B2(\u10_mem[1] [15]),
    .Y(n_11578));
 AOI22xp5_ASAP7_75t_SL g167125 (.A1(n_11548),
    .A2(\u10_mem[0] [9]),
    .B1(n_14825),
    .B2(\u10_mem[1] [9]),
    .Y(n_11579));
 AOI22xp5_ASAP7_75t_SL g167126 (.A1(n_11548),
    .A2(\u10_mem[0] [5]),
    .B1(n_14825),
    .B2(\u10_mem[1] [5]),
    .Y(n_11580));
 AOI22xp5_ASAP7_75t_SL g167129 (.A1(n_11583),
    .A2(\u11_mem[0] [7]),
    .B1(n_11477),
    .B2(\u11_mem[2] [7]),
    .Y(n_11584));
 AND2x6_ASAP7_75t_SL g167130 (.A(n_13764),
    .B(n_13027),
    .Y(n_11583));
 AOI22xp5_ASAP7_75t_SL g167131 (.A1(n_11583),
    .A2(\u11_mem[0] [11]),
    .B1(n_11477),
    .B2(\u11_mem[2] [11]),
    .Y(n_11585));
 AOI22xp5_ASAP7_75t_SL g167132 (.A1(n_11583),
    .A2(\u11_mem[0] [31]),
    .B1(n_11477),
    .B2(\u11_mem[2] [31]),
    .Y(n_11586));
 AOI22xp5_ASAP7_75t_SL g167133 (.A1(n_11583),
    .A2(\u11_mem[0] [21]),
    .B1(n_11477),
    .B2(\u11_mem[2] [21]),
    .Y(n_11587));
 AOI22xp5_ASAP7_75t_SL g167134 (.A1(n_11583),
    .A2(\u11_mem[0] [15]),
    .B1(n_11477),
    .B2(\u11_mem[2] [15]),
    .Y(n_11588));
 AOI22xp5_ASAP7_75t_SL g167135 (.A1(n_11583),
    .A2(\u11_mem[0] [1]),
    .B1(n_11477),
    .B2(\u11_mem[2] [1]),
    .Y(n_11589));
 AOI22xp5_ASAP7_75t_SL g167136 (.A1(n_11583),
    .A2(\u11_mem[0] [2]),
    .B1(n_11477),
    .B2(\u11_mem[2] [2]),
    .Y(n_11590));
 AOI22xp5_ASAP7_75t_SL g167137 (.A1(n_11583),
    .A2(\u11_mem[0] [5]),
    .B1(n_11477),
    .B2(\u11_mem[2] [5]),
    .Y(n_11591));
 AOI22xp33_ASAP7_75t_SL g167138 (.A1(n_11583),
    .A2(\u11_mem[0] [13]),
    .B1(n_11477),
    .B2(\u11_mem[2] [13]),
    .Y(n_11592));
 AOI22xp5_ASAP7_75t_SL g167139 (.A1(n_11583),
    .A2(\u11_mem[0] [4]),
    .B1(n_11477),
    .B2(\u11_mem[2] [4]),
    .Y(n_11593));
 AOI22xp5_ASAP7_75t_SL g167140 (.A1(n_11583),
    .A2(\u11_mem[0] [8]),
    .B1(n_11477),
    .B2(\u11_mem[2] [8]),
    .Y(n_11594));
 AOI22xp5_ASAP7_75t_SL g167141 (.A1(n_11583),
    .A2(\u11_mem[0] [25]),
    .B1(n_11477),
    .B2(\u11_mem[2] [25]),
    .Y(n_11595));
 AOI22xp33_ASAP7_75t_SL g167142 (.A1(n_11583),
    .A2(\u11_mem[0] [26]),
    .B1(n_11477),
    .B2(\u11_mem[2] [26]),
    .Y(n_11596));
 AOI22xp5_ASAP7_75t_SL g167143 (.A1(n_11583),
    .A2(\u11_mem[0] [10]),
    .B1(n_11477),
    .B2(\u11_mem[2] [10]),
    .Y(n_11597));
 AOI22xp33_ASAP7_75t_SL g167144 (.A1(n_11583),
    .A2(\u11_mem[0] [28]),
    .B1(n_11477),
    .B2(\u11_mem[2] [28]),
    .Y(n_11598));
 AOI22xp5_ASAP7_75t_SL g167145 (.A1(n_11583),
    .A2(\u11_mem[0] [20]),
    .B1(n_11477),
    .B2(\u11_mem[2] [20]),
    .Y(n_11599));
 AOI22xp5_ASAP7_75t_SL g167146 (.A1(n_11583),
    .A2(\u11_mem[0] [23]),
    .B1(n_11477),
    .B2(\u11_mem[2] [23]),
    .Y(n_11600));
 AOI22xp5_ASAP7_75t_SL g167147 (.A1(n_11583),
    .A2(\u11_mem[0] [24]),
    .B1(n_11477),
    .B2(\u11_mem[2] [24]),
    .Y(n_11601));
 AOI22xp5_ASAP7_75t_SL g167148 (.A1(n_11583),
    .A2(\u11_mem[0] [17]),
    .B1(n_11477),
    .B2(\u11_mem[2] [17]),
    .Y(n_11602));
 AOI22xp5_ASAP7_75t_SL g167149 (.A1(n_11583),
    .A2(\u11_mem[0] [22]),
    .B1(n_11477),
    .B2(\u11_mem[2] [22]),
    .Y(n_11603));
 AOI22xp5_ASAP7_75t_SL g167150 (.A1(n_11583),
    .A2(\u11_mem[0] [19]),
    .B1(n_11477),
    .B2(\u11_mem[2] [19]),
    .Y(n_11604));
 AOI22xp5_ASAP7_75t_SL g167151 (.A1(n_11583),
    .A2(\u11_mem[0] [18]),
    .B1(n_11477),
    .B2(\u11_mem[2] [18]),
    .Y(n_11605));
 AOI22xp5_ASAP7_75t_SL g167152 (.A1(n_11583),
    .A2(\u11_mem[0] [12]),
    .B1(n_11477),
    .B2(\u11_mem[2] [12]),
    .Y(n_11606));
 AOI22xp5_ASAP7_75t_SL g167153 (.A1(n_11583),
    .A2(\u11_mem[0] [9]),
    .B1(n_11477),
    .B2(\u11_mem[2] [9]),
    .Y(n_11607));
 AOI22xp5_ASAP7_75t_SL g167154 (.A1(n_11583),
    .A2(\u11_mem[0] [6]),
    .B1(n_11477),
    .B2(\u11_mem[2] [6]),
    .Y(n_11608));
 AOI22xp5_ASAP7_75t_SL g167155 (.A1(n_11583),
    .A2(\u11_mem[0] [0]),
    .B1(n_11477),
    .B2(\u11_mem[2] [0]),
    .Y(n_11609));
 AOI22xp5_ASAP7_75t_SL g167156 (.A1(n_11583),
    .A2(\u11_mem[0] [29]),
    .B1(n_11477),
    .B2(\u11_mem[2] [29]),
    .Y(n_11610));
 AOI22xp5_ASAP7_75t_SL g167157 (.A1(n_11583),
    .A2(\u11_mem[0] [30]),
    .B1(n_11477),
    .B2(\u11_mem[2] [30]),
    .Y(n_11611));
 AOI22xp5_ASAP7_75t_SL g167158 (.A1(n_11583),
    .A2(\u11_mem[0] [3]),
    .B1(n_11477),
    .B2(\u11_mem[2] [3]),
    .Y(n_11612));
 AOI22xp33_ASAP7_75t_SL g167159 (.A1(n_11583),
    .A2(\u11_mem[0] [16]),
    .B1(n_11477),
    .B2(\u11_mem[2] [16]),
    .Y(n_11613));
 AOI22xp5_ASAP7_75t_SL g167160 (.A1(n_11583),
    .A2(\u11_mem[0] [27]),
    .B1(n_11477),
    .B2(\u11_mem[2] [27]),
    .Y(n_11614));
 AOI22xp5_ASAP7_75t_SL g167161 (.A1(n_11583),
    .A2(\u11_mem[0] [14]),
    .B1(n_11477),
    .B2(\u11_mem[2] [14]),
    .Y(n_11615));
 AOI22xp5_ASAP7_75t_SL g167164 (.A1(n_11618),
    .A2(\u9_mem[0] [17]),
    .B1(n_11512),
    .B2(\u9_mem[2] [17]),
    .Y(n_11619));
 AND2x6_ASAP7_75t_SL g167165 (.A(n_13035),
    .B(n_13758),
    .Y(n_11618));
 AOI22xp5_ASAP7_75t_SL g167166 (.A1(n_11618),
    .A2(\u9_mem[0] [15]),
    .B1(n_11512),
    .B2(\u9_mem[2] [15]),
    .Y(n_11620));
 AOI22xp5_ASAP7_75t_SL g167167 (.A1(n_11618),
    .A2(\u9_mem[0] [11]),
    .B1(n_11512),
    .B2(\u9_mem[2] [11]),
    .Y(n_11621));
 AOI22xp5_ASAP7_75t_SL g167168 (.A1(n_11618),
    .A2(\u9_mem[0] [1]),
    .B1(n_11512),
    .B2(\u9_mem[2] [1]),
    .Y(n_11622));
 AOI22xp5_ASAP7_75t_SL g167169 (.A1(n_11618),
    .A2(\u9_mem[0] [21]),
    .B1(n_11512),
    .B2(\u9_mem[2] [21]),
    .Y(n_11623));
 AOI22xp5_ASAP7_75t_SL g167170 (.A1(n_11618),
    .A2(\u9_mem[0] [29]),
    .B1(n_11512),
    .B2(\u9_mem[2] [29]),
    .Y(n_11624));
 AOI22xp5_ASAP7_75t_SL g167171 (.A1(n_11618),
    .A2(\u9_mem[0] [28]),
    .B1(n_11512),
    .B2(\u9_mem[2] [28]),
    .Y(n_11625));
 AOI22xp5_ASAP7_75t_SL g167172 (.A1(n_11618),
    .A2(\u9_mem[0] [27]),
    .B1(n_11512),
    .B2(\u9_mem[2] [27]),
    .Y(n_11626));
 AOI22xp5_ASAP7_75t_SL g167173 (.A1(n_11618),
    .A2(\u9_mem[0] [26]),
    .B1(n_11512),
    .B2(\u9_mem[2] [26]),
    .Y(n_11627));
 AOI22xp5_ASAP7_75t_SL g167174 (.A1(n_11618),
    .A2(\u9_mem[0] [25]),
    .B1(n_11512),
    .B2(\u9_mem[2] [25]),
    .Y(n_11628));
 AOI22xp33_ASAP7_75t_SL g167175 (.A1(n_11618),
    .A2(\u9_mem[0] [22]),
    .B1(n_11512),
    .B2(\u9_mem[2] [22]),
    .Y(n_11629));
 AOI22xp5_ASAP7_75t_SL g167176 (.A1(n_11618),
    .A2(\u9_mem[0] [20]),
    .B1(n_11512),
    .B2(\u9_mem[2] [20]),
    .Y(n_11630));
 AOI22xp5_ASAP7_75t_SL g167177 (.A1(n_11618),
    .A2(\u9_mem[0] [18]),
    .B1(n_11512),
    .B2(\u9_mem[2] [18]),
    .Y(n_11631));
 AOI22xp5_ASAP7_75t_SL g167178 (.A1(n_11618),
    .A2(\u9_mem[0] [16]),
    .B1(n_11512),
    .B2(\u9_mem[2] [16]),
    .Y(n_11632));
 AOI22xp5_ASAP7_75t_SL g167179 (.A1(n_11618),
    .A2(\u9_mem[0] [30]),
    .B1(n_11512),
    .B2(\u9_mem[2] [30]),
    .Y(n_11633));
 AOI22xp5_ASAP7_75t_SL g167180 (.A1(n_11618),
    .A2(\u9_mem[0] [10]),
    .B1(n_11512),
    .B2(\u9_mem[2] [10]),
    .Y(n_11634));
 AOI22xp5_ASAP7_75t_SL g167181 (.A1(n_11618),
    .A2(\u9_mem[0] [8]),
    .B1(n_11512),
    .B2(\u9_mem[2] [8]),
    .Y(n_11635));
 AOI22xp33_ASAP7_75t_SL g167182 (.A1(n_11618),
    .A2(\u9_mem[0] [7]),
    .B1(n_11512),
    .B2(\u9_mem[2] [7]),
    .Y(n_11636));
 AOI22xp5_ASAP7_75t_SL g167183 (.A1(n_11618),
    .A2(\u9_mem[0] [6]),
    .B1(n_11512),
    .B2(\u9_mem[2] [6]),
    .Y(n_11637));
 AOI22xp5_ASAP7_75t_SL g167184 (.A1(n_11618),
    .A2(\u9_mem[0] [2]),
    .B1(n_11512),
    .B2(\u9_mem[2] [2]),
    .Y(n_11638));
 AOI22xp5_ASAP7_75t_SL g167185 (.A1(n_11618),
    .A2(\u9_mem[0] [24]),
    .B1(n_11512),
    .B2(\u9_mem[2] [24]),
    .Y(n_11639));
 AOI22xp5_ASAP7_75t_SL g167186 (.A1(n_11618),
    .A2(\u9_mem[0] [31]),
    .B1(n_11512),
    .B2(\u9_mem[2] [31]),
    .Y(n_11640));
 AOI22xp5_ASAP7_75t_SL g167187 (.A1(n_11618),
    .A2(\u9_mem[0] [4]),
    .B1(n_11512),
    .B2(\u9_mem[2] [4]),
    .Y(n_11641));
 AOI22xp5_ASAP7_75t_SL g167188 (.A1(n_11618),
    .A2(\u9_mem[0] [5]),
    .B1(n_11512),
    .B2(\u9_mem[2] [5]),
    .Y(n_11642));
 AOI22xp5_ASAP7_75t_SL g167189 (.A1(n_11618),
    .A2(\u9_mem[0] [23]),
    .B1(n_11512),
    .B2(\u9_mem[2] [23]),
    .Y(n_11643));
 AOI22xp5_ASAP7_75t_SL g167190 (.A1(n_11618),
    .A2(\u9_mem[0] [9]),
    .B1(n_11512),
    .B2(\u9_mem[2] [9]),
    .Y(n_11644));
 AOI22xp5_ASAP7_75t_SL g167191 (.A1(n_11618),
    .A2(\u9_mem[0] [13]),
    .B1(n_11512),
    .B2(\u9_mem[2] [13]),
    .Y(n_11645));
 AOI22xp5_ASAP7_75t_SL g167192 (.A1(n_11618),
    .A2(\u9_mem[0] [12]),
    .B1(n_11512),
    .B2(\u9_mem[2] [12]),
    .Y(n_11646));
 AOI22xp33_ASAP7_75t_SL g167193 (.A1(n_11618),
    .A2(\u9_mem[0] [14]),
    .B1(n_11512),
    .B2(\u9_mem[2] [14]),
    .Y(n_11647));
 AOI22xp5_ASAP7_75t_SL g167194 (.A1(n_11618),
    .A2(\u9_mem[0] [0]),
    .B1(n_11512),
    .B2(\u9_mem[2] [0]),
    .Y(n_11648));
 AOI22xp33_ASAP7_75t_SL g167195 (.A1(n_11618),
    .A2(\u9_mem[0] [19]),
    .B1(n_11512),
    .B2(\u9_mem[2] [19]),
    .Y(n_11649));
 AOI22xp5_ASAP7_75t_SL g167196 (.A1(n_11618),
    .A2(\u9_mem[0] [3]),
    .B1(n_11512),
    .B2(\u9_mem[2] [3]),
    .Y(n_11650));
 INVx1_ASAP7_75t_L g167218 (.A(in_slt4[18]),
    .Y(n_11693));
 HB1xp67_ASAP7_75t_L g167355 (.A(n_77853),
    .Y(n_11874));
 AND2x4_ASAP7_75t_SL g167452_dup (.A(n_26497),
    .B(n_26498),
    .Y(n_26501));
 AOI22xp5_ASAP7_75t_SL g167520 (.A1(\u6_mem[2] [8]),
    .A2(n_77853),
    .B1(\u6_mem[3] [8]),
    .B2(n_41152),
    .Y(n_12053));
 AOI22xp33_ASAP7_75t_SL g167528 (.A1(n_2693),
    .A2(n_41152),
    .B1(u6_rp[3]),
    .B2(n_12061),
    .Y(n_12062));
 INVxp67_ASAP7_75t_SL g167529 (.A(n_41152),
    .Y(n_12061));
 AOI22xp5_ASAP7_75t_SL g167533 (.A1(\u6_mem[2] [11]),
    .A2(n_77853),
    .B1(\u6_mem[3] [11]),
    .B2(n_41152),
    .Y(n_12066));
 NAND2xp5_ASAP7_75t_SL g167534 (.A(n_41152),
    .B(u6_rp[0]),
    .Y(n_12067));
 AOI22xp5_ASAP7_75t_L g167537 (.A1(n_77853),
    .A2(\u6_mem[2] [3]),
    .B1(n_41152),
    .B2(\u6_mem[3] [3]),
    .Y(n_12070));
 OAI21xp5_ASAP7_75t_SL g167562 (.A1(n_12097),
    .A2(oc3_cfg[2]),
    .B(n_34234),
    .Y(n_12098));
 INVx1_ASAP7_75t_SL g167564 (.A(n_12098),
    .Y(n_12100));
 HB1xp67_ASAP7_75t_R g167577 (.A(n_12116),
    .Y(n_12117));
 NAND2xp5_ASAP7_75t_SL g167578 (.A(in_valid_s[1]),
    .B(u14_u7_en_out_l_44),
    .Y(n_12116));
 NOR2xp33_ASAP7_75t_SL g167580 (.A(n_12116),
    .B(u14_u7_en_out_l2),
    .Y(n_12119));
 AND2x2_ASAP7_75t_SL g167603 (.A(u3_wp[0]),
    .B(o3_we),
    .Y(n_12142));
 NAND2x1p5_ASAP7_75t_SL g167604 (.A(u3_wp[0]),
    .B(o3_we),
    .Y(n_12143));
 AND2x4_ASAP7_75t_SL g167677 (.A(rf_we),
    .B(n_22851),
    .Y(n_12219));
 INVx1_ASAP7_75t_SL g167682 (.A(n_77797),
    .Y(n_12225));
 AOI31xp33_ASAP7_75t_SL g167684 (.A1(n_18896),
    .A2(n_77797),
    .A3(n_2694),
    .B(oc3_int_set[2]),
    .Y(n_12226));
 OAI22xp33_ASAP7_75t_SL g167685 (.A1(n_12225),
    .A2(u6_rp[0]),
    .B1(n_678),
    .B2(n_77797),
    .Y(n_12227));
 INVx1_ASAP7_75t_SL g167730 (.A(u4_wp[0]),
    .Y(n_12275));
 AOI22xp5_ASAP7_75t_SL g167858 (.A1(n_12403),
    .A2(n_10924),
    .B1(\u7_mem[0] [0]),
    .B2(n_3365),
    .Y(n_12404));
 BUFx12f_ASAP7_75t_SL g167859 (.A(n_43534),
    .Y(n_12403));
 AOI22xp5_ASAP7_75t_SL g167860 (.A1(n_12403),
    .A2(n_78044),
    .B1(\u7_mem[0] [1]),
    .B2(n_3365),
    .Y(n_12405));
 AOI22xp5_ASAP7_75t_SL g167861 (.A1(n_12403),
    .A2(n_28424),
    .B1(\u7_mem[0] [24]),
    .B2(n_3365),
    .Y(n_12406));
 AOI22xp5_ASAP7_75t_SL g167862 (.A1(n_12403),
    .A2(n_65902),
    .B1(\u7_mem[0] [31]),
    .B2(n_3386),
    .Y(n_12407));
 AOI22xp5_ASAP7_75t_SL g167863 (.A1(n_12403),
    .A2(n_28381),
    .B1(\u7_mem[0] [23]),
    .B2(n_3365),
    .Y(n_12408));
 AOI22xp5_ASAP7_75t_SL g167864 (.A1(n_73996),
    .A2(n_12403),
    .B1(\u7_mem[0] [21]),
    .B2(n_3365),
    .Y(n_12409));
 AOI22xp5_ASAP7_75t_SL g167865 (.A1(n_10196),
    .A2(n_12403),
    .B1(\u7_mem[0] [19]),
    .B2(n_3365),
    .Y(n_12410));
 AOI22xp5_ASAP7_75t_SL g167866 (.A1(n_10194),
    .A2(n_12403),
    .B1(\u7_mem[0] [18]),
    .B2(n_3365),
    .Y(n_12411));
 AOI22xp5_ASAP7_75t_SL g167867 (.A1(n_65952),
    .A2(n_12403),
    .B1(\u7_mem[0] [17]),
    .B2(n_3386),
    .Y(n_12412));
 AOI22xp5_ASAP7_75t_SL g167868 (.A1(n_28276),
    .A2(n_12403),
    .B1(\u7_mem[0] [16]),
    .B2(n_3386),
    .Y(n_12413));
 AOI22xp5_ASAP7_75t_SL g167869 (.A1(n_35041),
    .A2(n_12403),
    .B1(\u7_mem[0] [13]),
    .B2(n_3386),
    .Y(n_12414));
 AOI22xp5_ASAP7_75t_SL g167870 (.A1(n_12403),
    .A2(n_66869),
    .B1(\u7_mem[0] [5]),
    .B2(n_3386),
    .Y(n_12415));
 AOI22xp5_ASAP7_75t_SL g167872 (.A1(n_65980),
    .A2(n_12403),
    .B1(\u7_mem[0] [8]),
    .B2(n_3386),
    .Y(n_12417));
 AOI22xp5_ASAP7_75t_SL g167873 (.A1(n_28913),
    .A2(n_12403),
    .B1(\u7_mem[0] [15]),
    .B2(n_3386),
    .Y(n_12418));
 AOI22xp5_ASAP7_75t_SL g167874 (.A1(n_12403),
    .A2(n_28251),
    .B1(\u7_mem[0] [14]),
    .B2(n_3386),
    .Y(n_12419));
 AOI22xp5_ASAP7_75t_SL g167875 (.A1(n_12403),
    .A2(n_15952),
    .B1(\u7_mem[0] [29]),
    .B2(n_3365),
    .Y(n_12420));
 AOI22xp5_ASAP7_75t_SL g167876 (.A1(n_12403),
    .A2(n_10638),
    .B1(\u7_mem[0] [30]),
    .B2(n_3386),
    .Y(n_12421));
 AOI22xp5_ASAP7_75t_SL g167877 (.A1(n_65910),
    .A2(n_12403),
    .B1(\u7_mem[0] [27]),
    .B2(n_3365),
    .Y(n_12422));
 AOI22xp5_ASAP7_75t_SL g167878 (.A1(n_12403),
    .A2(n_66010),
    .B1(\u7_mem[0] [26]),
    .B2(n_3386),
    .Y(n_12423));
 AOI22xp5_ASAP7_75t_SL g167879 (.A1(n_12403),
    .A2(n_28316),
    .B1(\u7_mem[0] [25]),
    .B2(n_3386),
    .Y(n_12424));
 AOI22xp5_ASAP7_75t_SL g167880 (.A1(n_12403),
    .A2(n_65920),
    .B1(\u7_mem[0] [28]),
    .B2(n_3365),
    .Y(n_12425));
 AOI22xp5_ASAP7_75t_SL g167882 (.A1(n_12403),
    .A2(n_10247),
    .B1(\u7_mem[0] [20]),
    .B2(n_3365),
    .Y(n_12427));
 AOI22xp5_ASAP7_75t_SL g167883 (.A1(n_10026),
    .A2(n_12403),
    .B1(\u7_mem[0] [12]),
    .B2(n_3386),
    .Y(n_12428));
 AOI22xp5_ASAP7_75t_SL g167884 (.A1(n_12403),
    .A2(n_66843),
    .B1(\u7_mem[0] [11]),
    .B2(n_3386),
    .Y(n_12429));
 AOI22xp5_ASAP7_75t_SL g167886 (.A1(n_9942),
    .A2(n_12403),
    .B1(\u7_mem[0] [9]),
    .B2(n_3386),
    .Y(n_12431));
 AOI22xp5_ASAP7_75t_SL g167887 (.A1(n_12403),
    .A2(n_15867),
    .B1(\u7_mem[0] [3]),
    .B2(n_3365),
    .Y(n_12432));
 AOI22xp5_ASAP7_75t_SL g167888 (.A1(n_12403),
    .A2(n_66000),
    .B1(\u7_mem[0] [2]),
    .B2(n_3365),
    .Y(n_12433));
 AOI22xp5_ASAP7_75t_SL g167889 (.A1(n_17578),
    .A2(n_12403),
    .B1(\u7_mem[0] [7]),
    .B2(n_3365),
    .Y(n_12434));
 AOI22xp5_ASAP7_75t_SL g167890 (.A1(n_12403),
    .A2(n_32644),
    .B1(\u7_mem[0] [6]),
    .B2(n_3365),
    .Y(n_12435));
 AOI22xp33_ASAP7_75t_SL g167892 (.A1(wb_din[30]),
    .A2(n_67247),
    .B1(oc3_cfg[6]),
    .B2(n_67248),
    .Y(n_12438));
 AOI22xp5_ASAP7_75t_SL g167895 (.A1(n_62940),
    .A2(n_67247),
    .B1(n_78041),
    .B2(n_29621),
    .Y(n_12440));
 AOI22xp33_ASAP7_75t_SL g167897 (.A1(n_35437),
    .A2(n_67247),
    .B1(n_4027),
    .B2(n_29621),
    .Y(n_12441));
 AOI22xp5_ASAP7_75t_SL g167898 (.A1(n_65924),
    .A2(n_67247),
    .B1(oc3_cfg[1]),
    .B2(n_29621),
    .Y(n_12442));
 AOI22xp5_ASAP7_75t_SL g167900 (.A1(n_15920),
    .A2(n_67247),
    .B1(u13_occ0_r[31]),
    .B2(n_67248),
    .Y(n_12444));
 AOI22xp33_ASAP7_75t_SL g167901 (.A1(n_10198),
    .A2(n_67247),
    .B1(n_644),
    .B2(n_67248),
    .Y(n_12445));
 AOI22xp5_ASAP7_75t_SL g167903 (.A1(n_10143),
    .A2(n_67247),
    .B1(oc2_cfg[1]),
    .B2(n_67248),
    .Y(n_12447));
 AOI22xp5_ASAP7_75t_SL g167904 (.A1(n_65955),
    .A2(n_67247),
    .B1(n_18902),
    .B2(n_67248),
    .Y(n_12448));
 AOI22xp5_ASAP7_75t_SL g167906 (.A1(n_10026),
    .A2(n_67247),
    .B1(n_139),
    .B2(n_29621),
    .Y(n_12450));
 AOI22xp5_ASAP7_75t_SL g167908 (.A1(n_65969),
    .A2(n_67247),
    .B1(u13_occ0_r[7]),
    .B2(n_29621),
    .Y(n_12452));
 AOI22xp5_ASAP7_75t_SL g167909 (.A1(n_66032),
    .A2(n_67247),
    .B1(n_360),
    .B2(n_29621),
    .Y(n_12453));
 AOI22xp5_ASAP7_75t_SL g167910 (.A1(n_67247),
    .A2(n_32650),
    .B1(n_356),
    .B2(n_29621),
    .Y(n_12454));
 AOI22xp33_ASAP7_75t_SL g167911 (.A1(n_75733),
    .A2(n_67247),
    .B1(n_552),
    .B2(n_67248),
    .Y(n_12455));
 AOI22xp5_ASAP7_75t_SL g167912 (.A1(n_10891),
    .A2(n_67247),
    .B1(oc0_cfg[1]),
    .B2(n_29621),
    .Y(n_12456));
 AOI22xp33_ASAP7_75t_SL g167913 (.A1(wb_din[29]),
    .A2(n_67247),
    .B1(oc3_cfg[5]),
    .B2(n_67248),
    .Y(n_12457));
 AOI22xp5_ASAP7_75t_SL g167914 (.A1(n_65914),
    .A2(n_67247),
    .B1(n_198),
    .B2(n_67248),
    .Y(n_12458));
 AOI22xp5_ASAP7_75t_SL g167915 (.A1(n_28381),
    .A2(n_67247),
    .B1(u13_occ0_r[23]),
    .B2(n_67248),
    .Y(n_12459));
 AOI22xp33_ASAP7_75t_SL g167917 (.A1(n_66015),
    .A2(n_67247),
    .B1(oc2_cfg[5]),
    .B2(n_67248),
    .Y(n_12461));
 AOI22xp5_ASAP7_75t_SL g167919 (.A1(n_28276),
    .A2(n_67247),
    .B1(n_35577),
    .B2(n_29621),
    .Y(n_12463));
 AOI22xp5_ASAP7_75t_SL g167922 (.A1(n_79972),
    .A2(n_67247),
    .B1(n_357),
    .B2(n_29621),
    .Y(n_12466));
 AOI22xp5_ASAP7_75t_SL g167924 (.A1(n_15867),
    .A2(n_67247),
    .B1(n_573),
    .B2(n_29621),
    .Y(n_12468));
 AOI22xp5_ASAP7_75t_SL g167925 (.A1(n_28330),
    .A2(n_67247),
    .B1(n_4028),
    .B2(n_67248),
    .Y(n_12469));
 AOI22xp5_ASAP7_75t_SL g167926 (.A1(n_65990),
    .A2(n_67247),
    .B1(u13_occ0_r[15]),
    .B2(n_67248),
    .Y(n_12470));
 INVxp33_ASAP7_75t_R g168 (.A(wb_data_i[26]),
    .Y(n_66007));
 INVx4_ASAP7_75t_SL g168295 (.A(n_12868),
    .Y(n_12869));
 INVx4_ASAP7_75t_SL g168298 (.A(n_12868),
    .Y(n_12871));
 AOI22xp33_ASAP7_75t_SL g168313 (.A1(\u9_mem[2] [4]),
    .A2(n_5258),
    .B1(n_48642),
    .B2(n_12871),
    .Y(n_12887));
 INVx1_ASAP7_75t_SL g168335 (.A(n_625),
    .Y(n_12908));
 OR2x2_ASAP7_75t_SL g168393_dup (.A(n_26255),
    .B(n_22267),
    .Y(n_22183));
 INVx4_ASAP7_75t_SL g168438 (.A(u11_rp[0]),
    .Y(n_13027));
 INVx4_ASAP7_75t_SL g168446 (.A(u9_rp[0]),
    .Y(n_13035));
 AOI22xp5_ASAP7_75t_SL g168463 (.A1(n_65908),
    .A2(n_21549),
    .B1(\u3_mem[3] [27]),
    .B2(n_21550),
    .Y(n_13063));
 AOI22xp5_ASAP7_75t_SL g168465 (.A1(n_66010),
    .A2(n_21549),
    .B1(\u3_mem[3] [26]),
    .B2(n_21550),
    .Y(n_13064));
 AOI22xp5_ASAP7_75t_SL g168466 (.A1(n_65927),
    .A2(n_21549),
    .B1(\u3_mem[3] [25]),
    .B2(n_21550),
    .Y(n_13065));
 AOI22xp5_ASAP7_75t_SL g168467 (.A1(n_65915),
    .A2(n_21549),
    .B1(\u3_mem[3] [24]),
    .B2(n_21550),
    .Y(n_13066));
 AOI22xp5_ASAP7_75t_SL g168468 (.A1(n_65920),
    .A2(n_21549),
    .B1(\u3_mem[3] [28]),
    .B2(n_21550),
    .Y(n_13067));
 AOI22xp5_ASAP7_75t_SL g168469 (.A1(n_65902),
    .A2(n_21549),
    .B1(\u3_mem[3] [31]),
    .B2(n_21550),
    .Y(n_13068));
 AOI22xp5_ASAP7_75t_SL g168470 (.A1(n_65930),
    .A2(n_21549),
    .B1(\u3_mem[3] [23]),
    .B2(n_21550),
    .Y(n_13069));
 AOI22xp5_ASAP7_75t_SL g168471 (.A1(n_10660),
    .A2(n_21549),
    .B1(\u3_mem[3] [30]),
    .B2(n_21550),
    .Y(n_13070));
 AOI22xp5_ASAP7_75t_SL g168472 (.A1(n_10684),
    .A2(n_21549),
    .B1(\u3_mem[3] [29]),
    .B2(n_21550),
    .Y(n_13071));
 AOI22xp5_ASAP7_75t_SL g168473 (.A1(n_10302),
    .A2(n_21549),
    .B1(\u3_mem[3] [22]),
    .B2(n_21550),
    .Y(n_13072));
 AOI22xp33_ASAP7_75t_SL g168476 (.A1(n_66026),
    .A2(n_21549),
    .B1(\u3_mem[3] [20]),
    .B2(n_21550),
    .Y(n_13075));
 AOI22xp5_ASAP7_75t_SL g168477 (.A1(n_65932),
    .A2(n_21549),
    .B1(\u3_mem[3] [19]),
    .B2(n_21550),
    .Y(n_13076));
 AOI22xp33_ASAP7_75t_SL g168478 (.A1(n_10194),
    .A2(n_21549),
    .B1(\u3_mem[3] [18]),
    .B2(n_21550),
    .Y(n_13077));
 AOI22xp33_ASAP7_75t_SL g168480 (.A1(n_65949),
    .A2(n_21549),
    .B1(\u3_mem[3] [16]),
    .B2(n_21550),
    .Y(n_13079));
 AOI22xp33_ASAP7_75t_SL g168481 (.A1(n_28913),
    .A2(n_21527),
    .B1(\u3_mem[3] [15]),
    .B2(n_21550),
    .Y(n_13080));
 AOI22xp33_ASAP7_75t_SL g168482 (.A1(n_66032),
    .A2(n_21527),
    .B1(\u3_mem[3] [14]),
    .B2(n_21550),
    .Y(n_13081));
 AOI22xp33_ASAP7_75t_SL g168483 (.A1(n_35041),
    .A2(n_21527),
    .B1(\u3_mem[3] [13]),
    .B2(n_21550),
    .Y(n_13082));
 AOI22xp33_ASAP7_75t_SL g168484 (.A1(n_65997),
    .A2(n_21527),
    .B1(\u3_mem[3] [12]),
    .B2(n_21550),
    .Y(n_13083));
 AOI22xp33_ASAP7_75t_SL g168485 (.A1(n_66843),
    .A2(n_21527),
    .B1(\u3_mem[3] [11]),
    .B2(n_21550),
    .Y(n_13084));
 AOI22xp33_ASAP7_75t_SL g168486 (.A1(n_65975),
    .A2(n_21527),
    .B1(\u3_mem[3] [10]),
    .B2(n_21550),
    .Y(n_13085));
 AOI22xp5_ASAP7_75t_SL g168487 (.A1(n_79971),
    .A2(n_21527),
    .B1(\u3_mem[3] [9]),
    .B2(n_21550),
    .Y(n_13086));
 AOI22xp5_ASAP7_75t_SL g168488 (.A1(n_65980),
    .A2(n_21527),
    .B1(\u3_mem[3] [8]),
    .B2(n_21550),
    .Y(n_13087));
 AOI22xp33_ASAP7_75t_SL g168489 (.A1(n_65969),
    .A2(n_21527),
    .B1(\u3_mem[3] [7]),
    .B2(n_21550),
    .Y(n_13088));
 AOI22xp5_ASAP7_75t_SL g168490 (.A1(n_32644),
    .A2(n_21527),
    .B1(\u3_mem[3] [6]),
    .B2(n_21550),
    .Y(n_13089));
 AOI22xp5_ASAP7_75t_SL g168491 (.A1(n_66868),
    .A2(n_21527),
    .B1(\u3_mem[3] [5]),
    .B2(n_21550),
    .Y(n_13090));
 AOI22xp5_ASAP7_75t_SL g168493 (.A1(n_66856),
    .A2(n_21527),
    .B1(\u3_mem[3] [3]),
    .B2(n_21550),
    .Y(n_13092));
 AOI22xp5_ASAP7_75t_SL g168494 (.A1(n_66000),
    .A2(n_21527),
    .B1(\u3_mem[3] [2]),
    .B2(n_21550),
    .Y(n_13093));
 AOI22xp5_ASAP7_75t_SL g168495 (.A1(n_75733),
    .A2(n_21527),
    .B1(\u3_mem[3] [0]),
    .B2(n_21550),
    .Y(n_13094));
 AOI22xp5_ASAP7_75t_SL g168496 (.A1(n_3815),
    .A2(n_21527),
    .B1(\u3_mem[3] [1]),
    .B2(n_21550),
    .Y(n_13095));
 AND3x4_ASAP7_75t_SL g168541 (.A(u3_wp[0]),
    .B(o3_we),
    .C(n_48427),
    .Y(n_13176));
 NAND2xp5_ASAP7_75t_SL g168586 (.A(n_13236),
    .B(u11_din_tmp1[13]),
    .Y(n_13237));
 NAND2xp5_ASAP7_75t_SL g168594 (.A(u11_din_tmp1[8]),
    .B(n_13236),
    .Y(n_13244));
 NAND2xp5_ASAP7_75t_SL g168596 (.A(u11_din_tmp1[4]),
    .B(n_13236),
    .Y(n_13246));
 NAND2xp5_ASAP7_75t_SL g168597 (.A(u11_din_tmp1[5]),
    .B(n_13236),
    .Y(n_13247));
 NAND2xp5_ASAP7_75t_SL g168599 (.A(u11_din_tmp1[10]),
    .B(n_13236),
    .Y(n_13249));
 OAI21xp5_ASAP7_75t_SL g168615 (.A1(n_477),
    .A2(n_79193),
    .B(n_21343),
    .Y(n_13266));
 INVx1_ASAP7_75t_SL g168616 (.A(n_13266),
    .Y(n_13269));
 NOR5xp2_ASAP7_75t_SL g168648 (.A(n_31535),
    .B(n_1920),
    .C(n_1919),
    .D(n_1),
    .E(u2_res_cnt[3]),
    .Y(n_13347));
 INVx4_ASAP7_75t_SL g168710 (.A(n_21261),
    .Y(n_13420));
 NAND2x1_ASAP7_75t_SL g168800 (.A(n_13546),
    .B(n_805),
    .Y(n_13547));
 AOI22xp5_ASAP7_75t_SL g168801 (.A1(n_58959),
    .A2(\u4_mem[0] [15]),
    .B1(\u4_mem[1] [15]),
    .B2(n_50709),
    .Y(n_13546));
 AOI22xp5_ASAP7_75t_SL g168808 (.A1(\u3_mem[2] [6]),
    .A2(n_50342),
    .B1(\u3_mem[0] [6]),
    .B2(n_50341),
    .Y(n_13557));
 AOI21xp33_ASAP7_75t_SL g168834 (.A1(n_13594),
    .A2(n_13595),
    .B(n_17399),
    .Y(n_13597));
 NOR3xp33_ASAP7_75t_R g168835 (.A(n_8186),
    .B(u14_u6_full_empty_r),
    .C(n_4075),
    .Y(n_13595));
 INVx1_ASAP7_75t_L g168946 (.A(n_79203),
    .Y(n_13734));
 OAI211xp5_ASAP7_75t_SL g168948 (.A1(n_41434),
    .A2(n_13734),
    .B(n_13736),
    .C(n_13737),
    .Y(n_13738));
 AOI22xp33_ASAP7_75t_R g168950 (.A1(\u8_mem[2] [26]),
    .A2(n_51488),
    .B1(\u8_mem[3] [26]),
    .B2(n_14001),
    .Y(n_13736));
 AOI222xp33_ASAP7_75t_SL g168951 (.A1(n_36528),
    .A2(n_71352),
    .B1(\u8_mem[0] [26]),
    .B2(n_27133),
    .C1(\u8_mem[1] [26]),
    .C2(n_27134),
    .Y(n_13737));
 AOI22xp5_ASAP7_75t_SL g168955 (.A1(n_58959),
    .A2(\u4_mem[0] [14]),
    .B1(\u4_mem[2] [14]),
    .B2(n_35632),
    .Y(n_13742));
 XOR2xp5_ASAP7_75t_SL g168960 (.A(n_506),
    .B(n_46235),
    .Y(n_13749));
 NAND2xp5_ASAP7_75t_SL g168964 (.A(n_32381),
    .B(i3_re),
    .Y(n_13751));
 AOI22xp5_ASAP7_75t_SL g168968 (.A1(n_53101),
    .A2(\u5_mem[0] [17]),
    .B1(\u5_mem[2] [17]),
    .B2(n_65643),
    .Y(n_13755));
 INVx3_ASAP7_75t_SL g168971 (.A(u9_rp[1]),
    .Y(n_13758));
 INVx3_ASAP7_75t_SL g168974 (.A(u10_rp[1]),
    .Y(n_13761));
 INVx2_ASAP7_75t_SL g168976 (.A(u11_rp[1]),
    .Y(n_13764));
 INVx1_ASAP7_75t_SL g168980 (.A(u11_wp[2]),
    .Y(n_543));
 AOI21x1_ASAP7_75t_SL g168986 (.A1(n_36071),
    .A2(n_31726),
    .B(n_36073),
    .Y(n_13777));
 AND2x2_ASAP7_75t_SL g168994 (.A(n_1338),
    .B(n_1346),
    .Y(n_13787));
 NOR2xp33_ASAP7_75t_SL g168999 (.A(n_1186),
    .B(n_27061),
    .Y(n_13794));
 INVxp33_ASAP7_75t_R g169 (.A(wb_data_i[21]),
    .Y(n_66014));
 NOR2xp33_ASAP7_75t_SL g169001 (.A(n_10889),
    .B(n_27061),
    .Y(n_13796));
 INVx2_ASAP7_75t_SL g169019 (.A(n_35457),
    .Y(n_4548));
 NAND2x1_ASAP7_75t_SL g169025 (.A(n_13820),
    .B(n_13821),
    .Y(n_13822));
 AOI22xp5_ASAP7_75t_SL g169026 (.A1(n_58959),
    .A2(\u4_mem[0] [11]),
    .B1(\u4_mem[2] [11]),
    .B2(n_35632),
    .Y(n_13820));
 AOI22xp5_ASAP7_75t_SL g169027 (.A1(\u4_mem[1] [11]),
    .A2(n_50709),
    .B1(\u4_mem[3] [11]),
    .B2(n_30078),
    .Y(n_13821));
 NAND2xp5_ASAP7_75t_SL g169028 (.A(n_24350),
    .B(n_13822),
    .Y(n_13824));
 INVx1_ASAP7_75t_SL g169029 (.A(n_13822),
    .Y(n_13825));
 OAI22xp5_ASAP7_75t_SL g169031 (.A1(n_13758),
    .A2(u9_wp[2]),
    .B1(u9_rp[1]),
    .B2(n_259),
    .Y(n_13827));
 NAND2xp5_ASAP7_75t_L g169034 (.A(u9_rp[0]),
    .B(n_24737),
    .Y(n_13829));
 OAI22xp5_ASAP7_75t_SL g169049 (.A1(n_13761),
    .A2(u10_wp[2]),
    .B1(u10_rp[1]),
    .B2(n_234),
    .Y(n_13855));
 NAND2xp33_ASAP7_75t_L g169052 (.A(u10_rp[0]),
    .B(n_25438),
    .Y(n_13857));
 INVxp33_ASAP7_75t_SL g169092 (.A(n_4645),
    .Y(n_13899));
 NAND2xp5_ASAP7_75t_L g169135 (.A(out_slt3[6]),
    .B(n_5024),
    .Y(n_13955));
 NOR3xp33_ASAP7_75t_SL g169148 (.A(n_3468),
    .B(n_70322),
    .C(n_459),
    .Y(n_13968));
 AOI22xp5_ASAP7_75t_SL g169156 (.A1(n_77853),
    .A2(\u6_mem[2] [0]),
    .B1(n_41152),
    .B2(\u6_mem[3] [0]),
    .Y(n_13974));
 AOI22xp5_ASAP7_75t_SL g169163 (.A1(\u8_mem[3] [12]),
    .A2(n_78273),
    .B1(\u8_mem[1] [12]),
    .B2(n_78274),
    .Y(n_13982));
 AOI22xp5_ASAP7_75t_L g169164 (.A1(n_78274),
    .A2(\u8_mem[1] [9]),
    .B1(n_78273),
    .B2(\u8_mem[3] [9]),
    .Y(n_13983));
 AOI22xp5_ASAP7_75t_SL g169169 (.A1(\u8_mem[1] [19]),
    .A2(n_78274),
    .B1(\u8_mem[3] [19]),
    .B2(n_78273),
    .Y(n_13988));
 AOI22xp33_ASAP7_75t_L g169170 (.A1(n_78274),
    .A2(\u8_mem[1] [16]),
    .B1(n_78273),
    .B2(\u8_mem[3] [16]),
    .Y(n_13989));
 NAND2xp5_ASAP7_75t_SL g169171 (.A(n_78273),
    .B(u8_rp[0]),
    .Y(n_13990));
 AOI22xp33_ASAP7_75t_SL g169176 (.A1(n_78274),
    .A2(\u8_mem[1] [13]),
    .B1(n_78273),
    .B2(\u8_mem[3] [13]),
    .Y(n_13995));
 AOI22xp5_ASAP7_75t_SL g169180 (.A1(\u8_mem[1] [7]),
    .A2(n_78274),
    .B1(\u8_mem[3] [7]),
    .B2(n_78273),
    .Y(n_13999));
 AND2x4_ASAP7_75t_SL g169182 (.A(n_636),
    .B(n_78273),
    .Y(n_14001));
 AOI22xp5_ASAP7_75t_L g169184 (.A1(n_78274),
    .A2(\u8_mem[1] [5]),
    .B1(n_78273),
    .B2(\u8_mem[3] [5]),
    .Y(n_14003));
 NAND2x1_ASAP7_75t_SL g169186 (.A(n_14004),
    .B(n_21231),
    .Y(n_14006));
 AOI22xp5_ASAP7_75t_SL g169187 (.A1(n_50341),
    .A2(\u3_mem[0] [0]),
    .B1(\u3_mem[1] [0]),
    .B2(n_43317),
    .Y(n_14004));
 AO22x1_ASAP7_75t_SL g169195 (.A1(n_26427),
    .A2(n_11124),
    .B1(n_379),
    .B2(n_14012),
    .Y(n_14013));
 NAND2xp5_ASAP7_75t_SL g169200 (.A(n_13742),
    .B(n_1175),
    .Y(n_14017));
 OAI22xp33_ASAP7_75t_SL g169206 (.A1(n_65997),
    .A2(n_33772),
    .B1(n_14570),
    .B2(\u7_mem[3] [12]),
    .Y(n_14030));
 AOI21xp33_ASAP7_75t_SL g169219 (.A1(n_1177),
    .A2(n_58960),
    .B(n_8113),
    .Y(n_14054));
 AOI22xp5_ASAP7_75t_SL g169254 (.A1(n_78044),
    .A2(n_16797),
    .B1(ic0_cfg[1]),
    .B2(n_14098),
    .Y(n_14099));
 NAND2xp5_ASAP7_75t_SL g169257 (.A(rf_we),
    .B(n_8247),
    .Y(n_14098));
 NAND2xp5_ASAP7_75t_SL g169265 (.A(n_1041),
    .B(n_35633),
    .Y(n_14108));
 NOR4xp25_ASAP7_75t_SL g169382 (.A(n_778),
    .B(n_1084),
    .C(n_1086),
    .D(n_14226),
    .Y(n_14227));
 INVx1_ASAP7_75t_L g169431 (.A(in_slt4[11]),
    .Y(n_14280));
 INVx2_ASAP7_75t_R g169439 (.A(in_slt4[15]),
    .Y(n_14288));
 INVx1_ASAP7_75t_L g169443 (.A(in_slt4[6]),
    .Y(n_14292));
 INVx1_ASAP7_75t_R g169452 (.A(in_slt3[7]),
    .Y(n_14301));
 INVx2_ASAP7_75t_R g169460 (.A(in_slt6[13]),
    .Y(n_14309));
 INVx1_ASAP7_75t_R g169464 (.A(in_slt6[6]),
    .Y(n_14313));
 INVxp67_ASAP7_75t_SL g169471 (.A(n_295),
    .Y(n_14319));
 AND2x2_ASAP7_75t_R g169475 (.A(u15_rdd2),
    .B(n_28884),
    .Y(n_14324));
 NOR2xp33_ASAP7_75t_SL g169477 (.A(n_14325),
    .B(crac_rd_done),
    .Y(n_14326));
 INVxp33_ASAP7_75t_R g169478 (.A(u15_rdd3),
    .Y(n_14325));
 NOR2xp33_ASAP7_75t_R g169480 (.A(u14_u0_en_out_l2),
    .B(n_14431),
    .Y(n_14328));
 HB1xp67_ASAP7_75t_SL g169481 (.A(out_slt0[12]),
    .Y(n_1042));
 INVxp33_ASAP7_75t_R g169483 (.A(n_14431),
    .Y(n_14333));
 AND2x2_ASAP7_75t_R g169494 (.A(n_31581),
    .B(n_3937),
    .Y(n_14343));
 NOR2xp33_ASAP7_75t_R g169496 (.A(u14_u4_en_out_l2),
    .B(n_26182),
    .Y(n_14345));
 INVxp33_ASAP7_75t_R g169500 (.A(n_26182),
    .Y(n_14350));
 INVx2_ASAP7_75t_SL g169536 (.A(n_69796),
    .Y(n_14385));
 AOI22xp5_ASAP7_75t_SL g169540 (.A1(n_75733),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [0]),
    .Y(n_14390));
 AOI22xp5_ASAP7_75t_SL g169541 (.A1(n_32644),
    .A2(n_78410),
    .B1(n_22396),
    .B2(\u6_mem[1] [6]),
    .Y(n_14391));
 AOI22xp5_ASAP7_75t_SL g169542 (.A1(n_17578),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [7]),
    .Y(n_14392));
 AOI22xp5_ASAP7_75t_SL g169543 (.A1(n_66000),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [2]),
    .Y(n_14393));
 AOI22xp5_ASAP7_75t_SL g169544 (.A1(n_15867),
    .A2(n_78410),
    .B1(n_22396),
    .B2(\u6_mem[1] [3]),
    .Y(n_14394));
 AOI22xp5_ASAP7_75t_SL g169545 (.A1(n_65980),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [8]),
    .Y(n_14395));
 AOI22xp5_ASAP7_75t_SL g169546 (.A1(n_9942),
    .A2(n_78410),
    .B1(n_22396),
    .B2(\u6_mem[1] [9]),
    .Y(n_14396));
 AOI22xp5_ASAP7_75t_SL g169548 (.A1(n_10058),
    .A2(n_78410),
    .B1(\u6_mem[1] [5]),
    .B2(n_22396),
    .Y(n_14398));
 AOI22xp5_ASAP7_75t_SL g169549 (.A1(n_65955),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [13]),
    .Y(n_14399));
 AOI22xp5_ASAP7_75t_SL g169550 (.A1(n_78410),
    .A2(n_10143),
    .B1(n_31741),
    .B2(\u6_mem[1] [17]),
    .Y(n_14400));
 AOI22xp5_ASAP7_75t_SL g169551 (.A1(n_10171),
    .A2(n_78410),
    .B1(\u6_mem[1] [18]),
    .B2(n_22396),
    .Y(n_14401));
 AOI22xp33_ASAP7_75t_SL g169552 (.A1(n_10198),
    .A2(n_78410),
    .B1(n_22396),
    .B2(\u6_mem[1] [19]),
    .Y(n_14402));
 AOI22xp5_ASAP7_75t_SL g169553 (.A1(n_32916),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [21]),
    .Y(n_14403));
 AOI22xp33_ASAP7_75t_SL g169555 (.A1(n_3815),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [1]),
    .Y(n_14405));
 OAI31xp33_ASAP7_75t_SL g169567 (.A1(oc0_cfg[4]),
    .A2(o3_status[1]),
    .A3(o3_status[0]),
    .B(n_14431),
    .Y(n_14432));
 INVx1_ASAP7_75t_SL g169569 (.A(o3_empty),
    .Y(n_14431));
 INVx1_ASAP7_75t_SL g169660 (.A(n_488),
    .Y(n_14546));
 NOR2xp33_ASAP7_75t_SL g169752 (.A(n_14976),
    .B(n_402),
    .Y(n_14680));
 HB1xp67_ASAP7_75t_L g169816 (.A(n_64814),
    .Y(n_14765));
 NAND3xp33_ASAP7_75t_SL g169838 (.A(n_14791),
    .B(n_14788),
    .C(n_14789),
    .Y(n_14792));
 AND3x1_ASAP7_75t_L g169866 (.A(n_13761),
    .B(u10_rp[0]),
    .C(i4_re),
    .Y(n_14820));
 AND2x6_ASAP7_75t_SL g169867 (.A(u10_rp[1]),
    .B(n_25439),
    .Y(n_14821));
 AND2x6_ASAP7_75t_SL g169869 (.A(u10_rp[0]),
    .B(n_13761),
    .Y(n_14825));
 AOI22xp33_ASAP7_75t_SL g169903 (.A1(n_64793),
    .A2(\u5_mem[0] [27]),
    .B1(\u5_mem[1] [27]),
    .B2(n_6071),
    .Y(n_14859));
 OAI211xp5_ASAP7_75t_SL g169906 (.A1(n_4405),
    .A2(n_2524),
    .B(n_59759),
    .C(n_2247),
    .Y(n_14864));
 OAI22xp33_ASAP7_75t_SL g169945 (.A1(n_4024),
    .A2(n_6960),
    .B1(n_14902),
    .B2(n_10889),
    .Y(n_14904));
 INVx1_ASAP7_75t_SL g169946 (.A(oc1_cfg[2]),
    .Y(n_4024));
 INVxp67_ASAP7_75t_SL g169948 (.A(crac_din[10]),
    .Y(n_14902));
 OAI21xp5_ASAP7_75t_SL g169950 (.A1(n_6960),
    .A2(n_14906),
    .B(n_14907),
    .Y(n_14908));
 INVx2_ASAP7_75t_SL g169951 (.A(n_8308),
    .Y(n_6960));
 NAND2xp5_ASAP7_75t_SL g169953 (.A(n_10867),
    .B(crac_din[14]),
    .Y(n_14907));
 INVx3_ASAP7_75t_SL g169954 (.A(n_10867),
    .Y(n_14909));
 INVx1_ASAP7_75t_L g169955 (.A(oc1_cfg[6]),
    .Y(n_14906));
 OAI22xp33_ASAP7_75t_SL g169957 (.A1(n_262),
    .A2(n_6960),
    .B1(n_14912),
    .B2(n_14909),
    .Y(n_14913));
 INVxp67_ASAP7_75t_SL g169958 (.A(crac_din[9]),
    .Y(n_14912));
 NAND2xp5_ASAP7_75t_SL g169959 (.A(n_1932),
    .B(n_7772),
    .Y(n_14914));
 INVx1_ASAP7_75t_SL g169961 (.A(n_1932),
    .Y(n_14918));
 NAND2xp33_ASAP7_75t_L g169962 (.A(n_14924),
    .B(n_64852),
    .Y(n_14925));
 OAI211xp5_ASAP7_75t_SL g169963 (.A1(n_4568),
    .A2(n_14918),
    .B(n_37051),
    .C(n_14924),
    .Y(n_14926));
 AND3x4_ASAP7_75t_SL g169965 (.A(n_8334),
    .B(n_7195),
    .C(n_8256),
    .Y(n_14933));
 NAND2xp5_ASAP7_75t_SL g169967 (.A(n_42621),
    .B(n_14933),
    .Y(n_14935));
 OAI21xp33_ASAP7_75t_SL g169975 (.A1(n_14944),
    .A2(n_706),
    .B(n_43468),
    .Y(n_14945));
 AND2x2_ASAP7_75t_R g169976 (.A(u2_to_cnt[2]),
    .B(n_705),
    .Y(n_14944));
 OAI22xp33_ASAP7_75t_SL g169996 (.A1(u10_rp[2]),
    .A2(n_132),
    .B1(n_28774),
    .B2(u10_wp[3]),
    .Y(n_14976));
 INVx2_ASAP7_75t_SL g17 (.A(n_65978),
    .Y(n_9880));
 INVxp33_ASAP7_75t_R g170 (.A(wb_data_i[14]),
    .Y(n_66030));
 NAND3xp33_ASAP7_75t_SL g170000 (.A(n_14982),
    .B(n_14983),
    .C(n_46111),
    .Y(n_14985));
 AOI22xp5_ASAP7_75t_R g170001 (.A1(i6_dout[10]),
    .A2(n_14933),
    .B1(i3_dout[10]),
    .B2(n_8235),
    .Y(n_14982));
 AOI221xp5_ASAP7_75t_SL g170002 (.A1(n_7083),
    .A2(u13_intm_r[10]),
    .B1(i4_dout[10]),
    .B2(n_8174),
    .C(n_14904),
    .Y(n_14983));
 AND2x2_ASAP7_75t_SL g170016 (.A(n_15005),
    .B(n_49309),
    .Y(n_15007));
 NOR2xp33_ASAP7_75t_SL g170017 (.A(n_21341),
    .B(n_70322),
    .Y(n_15005));
 NOR2xp33_ASAP7_75t_SL g170032 (.A(dma_ack_i[1]),
    .B(n_14906),
    .Y(n_15020));
 OAI21xp33_ASAP7_75t_SL g170033 (.A1(n_2980),
    .A2(n_2522),
    .B(n_43083),
    .Y(n_15023));
 INVx1_ASAP7_75t_SL g170035 (.A(n_19069),
    .Y(n_15024));
 INVx1_ASAP7_75t_SL g170036 (.A(n_14432),
    .Y(n_15025));
 NOR2xp33_ASAP7_75t_SL g170038 (.A(dma_ack_i[0]),
    .B(n_257),
    .Y(n_15026));
 NOR3xp33_ASAP7_75t_SL g170041 (.A(n_117),
    .B(n_15031),
    .C(dma_ack_i[8]),
    .Y(n_15032));
 INVx1_ASAP7_75t_SL g170042 (.A(ic2_cfg[0]),
    .Y(n_117));
 INVx1_ASAP7_75t_R g170043 (.A(ic2_cfg[6]),
    .Y(n_15031));
 OAI21xp33_ASAP7_75t_SL g170044 (.A1(n_2371),
    .A2(n_2544),
    .B(ic2_cfg[0]),
    .Y(n_15034));
 INVxp33_ASAP7_75t_R g170049 (.A(dma_ack_i[4]),
    .Y(n_15037));
 OAI21xp33_ASAP7_75t_L g170050 (.A1(n_26183),
    .A2(n_2520),
    .B(n_41608),
    .Y(n_15040));
 OAI21xp33_ASAP7_75t_SL g170063 (.A1(n_70198),
    .A2(n_70199),
    .B(n_47740),
    .Y(n_15054));
 HB1xp67_ASAP7_75t_R g170065 (.A(n_24764),
    .Y(n_15056));
 INVx1_ASAP7_75t_SL g170076 (.A(n_28441),
    .Y(n_15079));
 AO21x1_ASAP7_75t_SL g170077 (.A1(n_13742),
    .A2(n_1175),
    .B(n_4548),
    .Y(n_15080));
 NAND2xp5_ASAP7_75t_SL g170083 (.A(n_1968),
    .B(n_573),
    .Y(n_15084));
 AOI22xp5_ASAP7_75t_SL g170084 (.A1(\u3_mem[2] [27]),
    .A2(n_77398),
    .B1(\u3_mem[3] [27]),
    .B2(n_22062),
    .Y(n_15085));
 AOI22xp33_ASAP7_75t_L g170086 (.A1(\u3_mem[0] [27]),
    .A2(n_24512),
    .B1(\u3_mem[1] [27]),
    .B2(n_24513),
    .Y(n_15087));
 NAND2xp5_ASAP7_75t_SL g170087 (.A(n_643),
    .B(n_42031),
    .Y(n_15090));
 NAND4xp25_ASAP7_75t_SL g170089 (.A(n_15090),
    .B(n_31870),
    .C(n_15092),
    .D(n_15093),
    .Y(n_15094));
 AOI22xp5_ASAP7_75t_SL g170091 (.A1(n_64793),
    .A2(\u5_mem[0] [31]),
    .B1(\u5_mem[1] [31]),
    .B2(n_6071),
    .Y(n_15092));
 AOI22xp33_ASAP7_75t_L g170092 (.A1(\u5_mem[2] [31]),
    .A2(n_1459),
    .B1(\u5_mem[3] [31]),
    .B2(n_56865),
    .Y(n_15093));
 INVx2_ASAP7_75t_L g170097 (.A(n_50290),
    .Y(n_15100));
 INVxp67_ASAP7_75t_L g170098 (.A(n_1840),
    .Y(n_15101));
 AOI22xp33_ASAP7_75t_SL g170131 (.A1(n_29006),
    .A2(n_15136),
    .B1(n_20594),
    .B2(\u11_mem[3] [2]),
    .Y(n_15137));
 NAND2xp5_ASAP7_75t_SL g170132 (.A(n_15135),
    .B(n_15134),
    .Y(n_15136));
 NAND2xp5_ASAP7_75t_L g170133 (.A(u11_din_tmp1[2]),
    .B(n_13236),
    .Y(n_15134));
 AOI22xp33_ASAP7_75t_SL g170134 (.A1(in_slt6[4]),
    .A2(n_1361),
    .B1(in_slt6[2]),
    .B2(n_1362),
    .Y(n_15135));
 AOI22xp33_ASAP7_75t_SL g170135 (.A1(n_29006),
    .A2(n_27878),
    .B1(n_20594),
    .B2(\u11_mem[3] [3]),
    .Y(n_15141));
 NAND2xp33_ASAP7_75t_L g170137 (.A(u11_din_tmp1[3]),
    .B(n_13236),
    .Y(n_15138));
 AOI22xp33_ASAP7_75t_SL g170138 (.A1(in_slt6[5]),
    .A2(n_1361),
    .B1(in_slt6[3]),
    .B2(n_1362),
    .Y(n_15139));
 AOI22xp5_ASAP7_75t_SL g170156 (.A1(n_22505),
    .A2(\u3_mem[1] [5]),
    .B1(n_66869),
    .B2(n_16009),
    .Y(n_15166));
 AOI21xp5_ASAP7_75t_SL g170215 (.A1(n_26541),
    .A2(u13_occ1_r[15]),
    .B(n_28814),
    .Y(n_15271));
 OR2x2_ASAP7_75t_L g170220 (.A(wb_addr_i[4]),
    .B(wb_addr_i[2]),
    .Y(n_15269));
 NOR2x1p5_ASAP7_75t_SL g170221 (.A(n_15269),
    .B(n_21335),
    .Y(n_15272));
 AOI22xp5_ASAP7_75t_SL g170222 (.A1(oc5_cfg[6]),
    .A2(n_26541),
    .B1(n_66032),
    .B2(n_15272),
    .Y(n_15274));
 AOI22xp5_ASAP7_75t_SL g170248 (.A1(n_556),
    .A2(n_26541),
    .B1(n_28240),
    .B2(n_15272),
    .Y(n_15300));
 AOI22xp5_ASAP7_75t_SL g170302 (.A1(n_22505),
    .A2(\u3_mem[1] [31]),
    .B1(n_15920),
    .B2(n_15143),
    .Y(n_15426));
 AOI22xp5_ASAP7_75t_SL g170345 (.A1(n_22577),
    .A2(\u3_mem[1] [8]),
    .B1(n_65980),
    .B2(n_16009),
    .Y(n_15469));
 AOI22xp5_ASAP7_75t_SL g170349 (.A1(n_22577),
    .A2(\u3_mem[1] [13]),
    .B1(n_65955),
    .B2(n_16009),
    .Y(n_15473));
 AOI22xp33_ASAP7_75t_SL g170351 (.A1(n_22577),
    .A2(\u3_mem[1] [24]),
    .B1(n_28424),
    .B2(n_15143),
    .Y(n_15475));
 AOI22xp33_ASAP7_75t_SL g170356 (.A1(n_22577),
    .A2(\u3_mem[1] [16]),
    .B1(n_28276),
    .B2(n_15143),
    .Y(n_15481));
 AOI22xp33_ASAP7_75t_SL g170358 (.A1(n_22577),
    .A2(\u3_mem[1] [7]),
    .B1(n_17578),
    .B2(n_16009),
    .Y(n_15483));
 AOI22xp33_ASAP7_75t_SL g170362 (.A1(n_22577),
    .A2(\u3_mem[1] [14]),
    .B1(n_28251),
    .B2(n_16009),
    .Y(n_15487));
 NAND2x1_ASAP7_75t_SL g170366 (.A(n_14003),
    .B(n_51490),
    .Y(n_15491));
 AOI22xp33_ASAP7_75t_SL g170378 (.A1(n_22505),
    .A2(\u3_mem[1] [9]),
    .B1(n_79971),
    .B2(n_16009),
    .Y(n_15506));
 AOI22xp33_ASAP7_75t_SL g170387 (.A1(n_22505),
    .A2(\u3_mem[1] [12]),
    .B1(n_10026),
    .B2(n_16009),
    .Y(n_15515));
 AOI22xp33_ASAP7_75t_SL g170393 (.A1(n_22505),
    .A2(\u3_mem[1] [17]),
    .B1(n_10143),
    .B2(n_15143),
    .Y(n_15521));
 AOI22xp33_ASAP7_75t_SL g170405 (.A1(n_22505),
    .A2(\u3_mem[1] [18]),
    .B1(n_10171),
    .B2(n_15143),
    .Y(n_15534));
 AOI22xp5_ASAP7_75t_SL g170621 (.A1(n_22505),
    .A2(\u3_mem[1] [27]),
    .B1(n_62940),
    .B2(n_15143),
    .Y(n_15771));
 AOI22xp5_ASAP7_75t_SL g170623 (.A1(n_22577),
    .A2(\u3_mem[1] [28]),
    .B1(n_22640),
    .B2(n_15143),
    .Y(n_15773));
 AOI22xp5_ASAP7_75t_SL g170625 (.A1(n_22577),
    .A2(\u3_mem[1] [23]),
    .B1(n_28381),
    .B2(n_15143),
    .Y(n_15775));
 AOI22xp33_ASAP7_75t_SL g170689 (.A1(n_22577),
    .A2(\u3_mem[1] [26]),
    .B1(n_35437),
    .B2(n_15143),
    .Y(n_15854));
 INVx3_ASAP7_75t_SL g170703 (.A(n_9851),
    .Y(n_15867));
 AOI22xp5_ASAP7_75t_SL g170740 (.A1(n_28316),
    .A2(n_73997),
    .B1(\u8_mem[1] [25]),
    .B2(n_75735),
    .Y(n_15915));
 AOI22xp5_ASAP7_75t_SL g170748 (.A1(n_15920),
    .A2(n_73997),
    .B1(\u8_mem[1] [31]),
    .B2(n_75735),
    .Y(n_15923));
 INVx3_ASAP7_75t_SL g170749 (.A(n_10330),
    .Y(n_15920));
 AOI22xp5_ASAP7_75t_SL g170754 (.A1(n_33024),
    .A2(n_73997),
    .B1(\u8_mem[1] [20]),
    .B2(n_31464),
    .Y(n_15931));
 AND2x4_ASAP7_75t_SL g170821 (.A(n_48675),
    .B(n_12142),
    .Y(n_16009));
 AOI22xp5_ASAP7_75t_SL g170840 (.A1(n_22505),
    .A2(\u3_mem[1] [25]),
    .B1(n_28316),
    .B2(n_15143),
    .Y(n_16031));
 INVxp33_ASAP7_75t_R g171 (.A(wb_data_i[31]),
    .Y(n_65898));
 AOI22xp33_ASAP7_75t_SL g171075 (.A1(n_22505),
    .A2(\u3_mem[1] [11]),
    .B1(n_66842),
    .B2(n_16009),
    .Y(n_16304));
 AOI22xp5_ASAP7_75t_SL g171085 (.A1(\u8_mem[1] [16]),
    .A2(n_31460),
    .B1(n_28276),
    .B2(n_73997),
    .Y(n_16314));
 AOI22xp33_ASAP7_75t_SL g171168 (.A1(n_22577),
    .A2(\u3_mem[1] [2]),
    .B1(n_66000),
    .B2(n_16009),
    .Y(n_16416));
 AOI22xp33_ASAP7_75t_SL g171179 (.A1(n_22505),
    .A2(\u3_mem[1] [19]),
    .B1(n_10198),
    .B2(n_15143),
    .Y(n_16427));
 AOI22xp5_ASAP7_75t_SL g171189 (.A1(n_28953),
    .A2(n_31777),
    .B1(n_20593),
    .B2(\u11_mem[1] [9]),
    .Y(n_16439));
 OAI22xp5_ASAP7_75t_SL g171192 (.A1(n_36288),
    .A2(n_1705),
    .B1(n_21631),
    .B2(n_1679),
    .Y(n_16436));
 NAND2xp5_ASAP7_75t_SL g171209 (.A(n_51499),
    .B(n_23296),
    .Y(n_16458));
 AOI22xp33_ASAP7_75t_SL g171322 (.A1(n_22505),
    .A2(\u3_mem[1] [15]),
    .B1(n_28913),
    .B2(n_15143),
    .Y(n_16593));
 AOI22xp5_ASAP7_75t_SL g171378 (.A1(n_46477),
    .A2(\u10_mem[0] [19]),
    .B1(n_46478),
    .B2(n_50551),
    .Y(n_16664));
 AND2x2_ASAP7_75t_SL g171388 (.A(n_16671),
    .B(n_1244),
    .Y(n_16672));
 AOI22xp33_ASAP7_75t_SL g171389 (.A1(\u3_mem[0] [4]),
    .A2(n_50341),
    .B1(n_50388),
    .B2(\u3_mem[2] [4]),
    .Y(n_16671));
 AOI22xp5_ASAP7_75t_SL g171394 (.A1(n_65941),
    .A2(n_73997),
    .B1(\u8_mem[1] [22]),
    .B2(n_31460),
    .Y(n_16680));
 AOI22xp5_ASAP7_75t_SL g171397 (.A1(n_28381),
    .A2(n_73997),
    .B1(\u8_mem[1] [23]),
    .B2(n_31460),
    .Y(n_16684));
 NAND4xp25_ASAP7_75t_SL g171435 (.A(n_28901),
    .B(n_16720),
    .C(n_16721),
    .D(n_16722),
    .Y(n_16723));
 AOI21xp5_ASAP7_75t_SL g171436 (.A1(n_2095),
    .A2(n_10614),
    .B(n_10888),
    .Y(n_16720));
 AOI22xp5_ASAP7_75t_R g171437 (.A1(i4_dout[8]),
    .A2(n_8174),
    .B1(n_7083),
    .B2(n_301),
    .Y(n_16721));
 NAND3xp33_ASAP7_75t_SL g171438 (.A(n_16724),
    .B(n_2418),
    .C(n_7207),
    .Y(n_16725));
 AOI21xp33_ASAP7_75t_SL g171439 (.A1(n_10614),
    .A2(u13_ints_r[0]),
    .B(n_11012),
    .Y(n_16724));
 NAND4xp25_ASAP7_75t_SL g171440 (.A(n_16726),
    .B(n_10635),
    .C(n_16727),
    .D(n_7204),
    .Y(n_16728));
 AOI22xp5_ASAP7_75t_R g171441 (.A1(i4_dout[6]),
    .A2(n_8174),
    .B1(n_7083),
    .B2(u13_intm_r[6]),
    .Y(n_16727));
 NAND4xp25_ASAP7_75t_SL g171442 (.A(n_16730),
    .B(n_31732),
    .C(n_16731),
    .D(n_16732),
    .Y(n_16733));
 AOI21xp5_ASAP7_75t_SL g171445 (.A1(n_37200),
    .A2(n_41637),
    .B(n_16738),
    .Y(n_16739));
 OAI22xp5_ASAP7_75t_SL g171446 (.A1(n_64994),
    .A2(n_16736),
    .B1(n_16737),
    .B2(n_64993),
    .Y(n_16738));
 INVxp33_ASAP7_75t_R g171447 (.A(\u5_mem[0] [26]),
    .Y(n_16736));
 INVxp33_ASAP7_75t_R g171448 (.A(\u5_mem[1] [26]),
    .Y(n_16737));
 NAND2xp5_ASAP7_75t_SL g171451 (.A(n_78810),
    .B(n_34203),
    .Y(n_16749));
 AOI22xp33_ASAP7_75t_L g171452 (.A1(\u6_mem[1] [24]),
    .A2(n_48415),
    .B1(\u6_mem[3] [24]),
    .B2(n_17704),
    .Y(n_16750));
 NAND2xp5_ASAP7_75t_L g171453 (.A(n_12097),
    .B(n_34190),
    .Y(n_16751));
 AND2x2_ASAP7_75t_SL g171468 (.A(n_56859),
    .B(n_13755),
    .Y(n_16781));
 AOI22xp5_ASAP7_75t_SL g171473 (.A1(crac_out[20]),
    .A2(n_56881),
    .B1(n_66026),
    .B2(n_12219),
    .Y(n_16788));
 AND2x4_ASAP7_75t_SL g171483 (.A(n_6615),
    .B(rf_we),
    .Y(n_16797));
 INVxp33_ASAP7_75t_L g171484 (.A(n_15031),
    .Y(n_16798));
 AOI22xp5_ASAP7_75t_SL g171489 (.A1(n_16805),
    .A2(n_56879),
    .B1(n_10143),
    .B2(n_17579),
    .Y(n_16807));
 INVxp33_ASAP7_75t_R g171490 (.A(n_1322),
    .Y(n_16805));
 AOI22xp5_ASAP7_75t_SL g171492 (.A1(crac_out[31]),
    .A2(n_56879),
    .B1(n_65902),
    .B2(n_12219),
    .Y(n_16816));
 AOI22xp5_ASAP7_75t_SL g171495 (.A1(crac_out[16]),
    .A2(n_56879),
    .B1(n_65949),
    .B2(n_17579),
    .Y(n_16819));
 AOI22xp5_ASAP7_75t_SL g171504 (.A1(crac_out[19]),
    .A2(n_56879),
    .B1(n_10198),
    .B2(n_17579),
    .Y(n_16828));
 AOI21xp5_ASAP7_75t_SL g171521 (.A1(n_72062),
    .A2(n_72063),
    .B(n_16857),
    .Y(n_16858));
 NAND2xp5_ASAP7_75t_SL g171526 (.A(n_14763),
    .B(n_78135),
    .Y(n_16853));
 OAI21xp33_ASAP7_75t_SL g171528 (.A1(n_477),
    .A2(n_57084),
    .B(n_78936),
    .Y(n_16857));
 NOR2xp33_ASAP7_75t_SL g171550 (.A(n_51041),
    .B(n_19495),
    .Y(n_16880));
 NOR2xp33_ASAP7_75t_SL g171562 (.A(n_40417),
    .B(n_4261),
    .Y(n_16895));
 NAND3xp33_ASAP7_75t_SL g171722 (.A(n_31750),
    .B(n_19578),
    .C(n_2286),
    .Y(n_17079));
 O2A1O1Ixp5_ASAP7_75t_SL g171748 (.A1(n_17108),
    .A2(n_24580),
    .B(n_5077),
    .C(n_4457),
    .Y(n_17110));
 OAI21xp33_ASAP7_75t_SL g171749 (.A1(n_15100),
    .A2(n_27224),
    .B(n_2500),
    .Y(n_17108));
 O2A1O1Ixp5_ASAP7_75t_SL g171872 (.A1(n_24553),
    .A2(n_17252),
    .B(n_5077),
    .C(n_27227),
    .Y(n_17254));
 OAI21xp33_ASAP7_75t_SL g171873 (.A1(n_15100),
    .A2(n_2498),
    .B(n_27223),
    .Y(n_17252));
 INVx2_ASAP7_75t_SL g171917_dup (.A(n_38363),
    .Y(n_38374));
 AOI22xp5_ASAP7_75t_SL g172 (.A1(n_66026),
    .A2(n_15143),
    .B1(n_22577),
    .B2(\u3_mem[1] [20]),
    .Y(n_15145));
 AOI221xp5_ASAP7_75t_SL g172003 (.A1(u13_intm_r[9]),
    .A2(n_7082),
    .B1(n_8174),
    .B2(i4_dout[9]),
    .C(n_14913),
    .Y(n_17388));
 AOI21xp5_ASAP7_75t_SL g172010 (.A1(n_17400),
    .A2(n_17399),
    .B(ic0_int_set[2]),
    .Y(n_17401));
 NOR2xp33_ASAP7_75t_SL g172012 (.A(n_2226),
    .B(n_306),
    .Y(n_17400));
 NOR2xp33_ASAP7_75t_SL g172013 (.A(n_306),
    .B(n_7582),
    .Y(n_17402));
 INVxp33_ASAP7_75t_R g172014 (.A(n_2226),
    .Y(n_17403));
 NAND2xp5_ASAP7_75t_SL g172047 (.A(n_43468),
    .B(n_17440),
    .Y(n_17441));
 XOR2xp5_ASAP7_75t_SL g172048 (.A(n_1648),
    .B(n_1647),
    .Y(n_17440));
 OAI211xp5_ASAP7_75t_SL g172095 (.A1(n_46227),
    .A2(n_17489),
    .B(n_17490),
    .C(n_20759),
    .Y(n_17492));
 NAND2xp5_ASAP7_75t_SL g172097 (.A(n_18709),
    .B(n_425),
    .Y(n_17490));
 AOI22xp5_ASAP7_75t_SL g172114 (.A1(crac_out[1]),
    .A2(n_28367),
    .B1(n_12219),
    .B2(n_78044),
    .Y(n_17513));
 AOI22xp5_ASAP7_75t_SL g172124 (.A1(crac_out[8]),
    .A2(n_28367),
    .B1(n_65980),
    .B2(n_17579),
    .Y(n_17530));
 AOI22xp5_ASAP7_75t_SL g172126 (.A1(crac_out[2]),
    .A2(n_28367),
    .B1(n_66000),
    .B2(n_17579),
    .Y(n_17532));
 AOI22xp5_ASAP7_75t_SL g172128 (.A1(crac_out[14]),
    .A2(n_28367),
    .B1(n_66032),
    .B2(n_17579),
    .Y(n_17534));
 AOI22xp5_ASAP7_75t_SL g172136 (.A1(crac_out[15]),
    .A2(n_28367),
    .B1(n_28913),
    .B2(n_17579),
    .Y(n_17542));
 AOI22xp5_ASAP7_75t_SL g172155 (.A1(crac_out[3]),
    .A2(n_28367),
    .B1(n_15867),
    .B2(n_17579),
    .Y(n_17563));
 AOI22xp5_ASAP7_75t_SL g172157 (.A1(crac_out[9]),
    .A2(n_28367),
    .B1(n_17579),
    .B2(n_9942),
    .Y(n_17565));
 AOI22xp5_ASAP7_75t_SL g172159 (.A1(crac_out[5]),
    .A2(n_28367),
    .B1(n_17579),
    .B2(n_10058),
    .Y(n_17567));
 NOR2xp33_ASAP7_75t_SL g172163 (.A(n_37935),
    .B(n_41376),
    .Y(n_17569));
 OAI21xp5_ASAP7_75t_SL g172165 (.A1(n_32164),
    .A2(n_17573),
    .B(n_35577),
    .Y(n_17575));
 AND2x4_ASAP7_75t_SL g172166_dup (.A(n_32162),
    .B(n_675),
    .Y(n_32164));
 NOR2xp33_ASAP7_75t_R g172167 (.A(n_32162),
    .B(n_675),
    .Y(n_17573));
 AOI22xp5_ASAP7_75t_SL g172169 (.A1(crac_out[11]),
    .A2(n_28367),
    .B1(n_12219),
    .B2(n_10000),
    .Y(n_17577));
 INVx3_ASAP7_75t_SL g172172 (.A(n_9793),
    .Y(n_17578));
 AND2x4_ASAP7_75t_SL g172173 (.A(n_22851),
    .B(rf_we),
    .Y(n_17579));
 AOI22xp5_ASAP7_75t_SL g172175 (.A1(crac_out[13]),
    .A2(n_28367),
    .B1(n_35041),
    .B2(n_17579),
    .Y(n_17583));
 INVx1_ASAP7_75t_SL g172177 (.A(n_427),
    .Y(n_17584));
 OAI221xp5_ASAP7_75t_SL g172183 (.A1(n_14301),
    .A2(n_24883),
    .B1(n_1714),
    .B2(n_48057),
    .C(n_48645),
    .Y(n_17591));
 OA22x2_ASAP7_75t_SL g172187 (.A1(n_34492),
    .A2(n_48057),
    .B1(n_1820),
    .B2(n_24883),
    .Y(n_17594));
 OAI221xp5_ASAP7_75t_SL g172188 (.A1(n_24883),
    .A2(n_48052),
    .B1(n_48057),
    .B2(n_21673),
    .C(n_48646),
    .Y(n_17595));
 OAI221xp5_ASAP7_75t_SL g172189 (.A1(n_24883),
    .A2(n_34492),
    .B1(n_48057),
    .B2(n_34500),
    .C(n_48647),
    .Y(n_17596));
 OAI221xp5_ASAP7_75t_SL g172190 (.A1(n_24883),
    .A2(n_48056),
    .B1(n_48057),
    .B2(n_34488),
    .C(n_48638),
    .Y(n_17597));
 OAI221xp5_ASAP7_75t_SL g172192 (.A1(n_34500),
    .A2(n_24883),
    .B1(n_34504),
    .B2(n_48057),
    .C(n_48644),
    .Y(n_17599));
 INVx1_ASAP7_75t_SL g172193 (.A(n_336),
    .Y(n_17600));
 BUFx3_ASAP7_75t_SL g172200 (.A(n_17600),
    .Y(n_17606));
 NOR2xp67_ASAP7_75t_SL g172201 (.A(n_26827),
    .B(n_17606),
    .Y(n_17608));
 OAI22xp5_ASAP7_75t_SL g172202 (.A1(n_21878),
    .A2(n_330),
    .B1(n_14280),
    .B2(n_17606),
    .Y(n_17609));
 OAI221xp5_ASAP7_75t_SL g172206 (.A1(n_17606),
    .A2(n_21878),
    .B1(n_14288),
    .B2(n_330),
    .C(n_1201),
    .Y(n_17613));
 OAI221xp5_ASAP7_75t_SL g172207 (.A1(n_17606),
    .A2(n_21669),
    .B1(n_26807),
    .B2(n_330),
    .C(n_1214),
    .Y(n_17614));
 OAI221xp5_ASAP7_75t_SL g172208 (.A1(n_17606),
    .A2(n_14288),
    .B1(n_330),
    .B2(n_26811),
    .C(n_1208),
    .Y(n_17615));
 INVxp33_ASAP7_75t_L g172209 (.A(n_24594),
    .Y(n_17616));
 AND2x2_ASAP7_75t_SL g172210 (.A(n_51493),
    .B(n_13999),
    .Y(n_17617));
 NAND2xp33_ASAP7_75t_SL g172211 (.A(n_51493),
    .B(n_13999),
    .Y(n_17618));
 NAND2xp5_ASAP7_75t_SL g172216 (.A(n_36008),
    .B(n_35632),
    .Y(n_17623));
 OAI21xp33_ASAP7_75t_SL g172217 (.A1(n_59339),
    .A2(n_56),
    .B(n_17625),
    .Y(n_17626));
 AOI21xp5_ASAP7_75t_SL g172218 (.A1(\u5_mem[3] [28]),
    .A2(n_56865),
    .B(n_1770),
    .Y(n_17625));
 XNOR2xp5_ASAP7_75t_SL g172262 (.A(n_29366),
    .B(n_43077),
    .Y(n_17672));
 BUFx2_ASAP7_75t_SL g172264 (.A(n_29934),
    .Y(n_17686));
 INVx2_ASAP7_75t_SL g172266 (.A(n_29934),
    .Y(n_17687));
 NOR2xp33_ASAP7_75t_SL g172267 (.A(n_29934),
    .B(n_8306),
    .Y(n_17688));
 NOR3xp33_ASAP7_75t_L g172269 (.A(n_13761),
    .B(n_29934),
    .C(i4_re),
    .Y(n_17690));
 AND2x4_ASAP7_75t_SL g172283 (.A(n_37337),
    .B(n_41152),
    .Y(n_17704));
 NAND4xp25_ASAP7_75t_SL g172284 (.A(n_28371),
    .B(n_2098),
    .C(n_17705),
    .D(n_1403),
    .Y(n_17706));
 AOI22xp5_ASAP7_75t_L g172285 (.A1(n_48415),
    .A2(\u6_mem[1] [27]),
    .B1(\u6_mem[3] [27]),
    .B2(n_17704),
    .Y(n_17705));
 INVxp67_ASAP7_75t_SL g172292 (.A(n_18684),
    .Y(n_17711));
 AOI22xp5_ASAP7_75t_SL g172326 (.A1(n_35041),
    .A2(n_64819),
    .B1(\u8_mem[3] [13]),
    .B2(n_70622),
    .Y(n_17778));
 AOI22xp5_ASAP7_75t_SL g172330 (.A1(n_28240),
    .A2(n_64818),
    .B1(n_70622),
    .B2(\u8_mem[3] [8]),
    .Y(n_17785));
 AOI22xp5_ASAP7_75t_SL g172332 (.A1(n_65949),
    .A2(n_64818),
    .B1(\u8_mem[3] [16]),
    .B2(n_70622),
    .Y(n_17787));
 AOI22xp33_ASAP7_75t_SL g172336 (.A1(n_65972),
    .A2(n_64818),
    .B1(\u8_mem[3] [10]),
    .B2(n_70622),
    .Y(n_17801));
 AOI22xp5_ASAP7_75t_SL g172340 (.A1(n_32644),
    .A2(n_64819),
    .B1(n_70622),
    .B2(\u8_mem[3] [6]),
    .Y(n_17809));
 AOI22xp5_ASAP7_75t_SL g172431 (.A1(n_46587),
    .A2(\u9_mem[0] [18]),
    .B1(n_31720),
    .B2(n_49625),
    .Y(n_17927));
 NOR2x2_ASAP7_75t_SL g172433 (.A(n_17924),
    .B(n_13420),
    .Y(n_17925));
 BUFx2_ASAP7_75t_L g172434 (.A(n_522),
    .Y(n_17924));
 AOI22xp5_ASAP7_75t_SL g172438 (.A1(n_9942),
    .A2(n_64818),
    .B1(\u8_mem[3] [9]),
    .B2(n_70622),
    .Y(n_17938));
 AOI22xp5_ASAP7_75t_SL g172475 (.A1(n_66868),
    .A2(n_64819),
    .B1(\u8_mem[3] [5]),
    .B2(n_70622),
    .Y(n_17979));
 AOI22xp5_ASAP7_75t_SL g172501 (.A1(n_17578),
    .A2(n_64818),
    .B1(\u8_mem[3] [7]),
    .B2(n_70622),
    .Y(n_18018));
 AOI22xp5_ASAP7_75t_SL g172533 (.A1(n_15867),
    .A2(n_64819),
    .B1(\u8_mem[3] [3]),
    .B2(n_70622),
    .Y(n_18058));
 AOI22xp5_ASAP7_75t_SL g172535 (.A1(n_66843),
    .A2(n_64819),
    .B1(\u8_mem[3] [11]),
    .B2(n_70622),
    .Y(n_18060));
 AOI22xp5_ASAP7_75t_SL g172541 (.A1(n_46478),
    .A2(n_18707),
    .B1(\u10_mem[0] [9]),
    .B2(n_46477),
    .Y(n_18068));
 OA22x2_ASAP7_75t_SL g172542 (.A1(n_14280),
    .A2(n_330),
    .B1(n_26815),
    .B2(n_17606),
    .Y(n_18066));
 AOI22xp5_ASAP7_75t_SL g172560 (.A1(n_29006),
    .A2(n_31779),
    .B1(n_20594),
    .B2(\u11_mem[3] [14]),
    .Y(n_18092));
 OAI22xp5_ASAP7_75t_SL g172563 (.A1(n_1681),
    .A2(n_1705),
    .B1(n_1704),
    .B2(n_1679),
    .Y(n_18089));
 AOI22xp5_ASAP7_75t_SL g172635 (.A1(n_28251),
    .A2(n_64818),
    .B1(\u8_mem[3] [14]),
    .B2(n_70622),
    .Y(n_18195));
 AOI22xp5_ASAP7_75t_SL g172710 (.A1(n_66000),
    .A2(n_64819),
    .B1(\u8_mem[3] [2]),
    .B2(n_70622),
    .Y(n_18289));
 AOI22xp5_ASAP7_75t_SL g172840 (.A1(n_28913),
    .A2(n_64819),
    .B1(n_70622),
    .B2(\u8_mem[3] [15]),
    .Y(n_18448));
 AOI22xp5_ASAP7_75t_SL g172860 (.A1(n_28953),
    .A2(n_31781),
    .B1(n_20593),
    .B2(\u11_mem[1] [12]),
    .Y(n_18483));
 OAI22xp5_ASAP7_75t_SL g172863 (.A1(n_1704),
    .A2(n_1705),
    .B1(n_21646),
    .B2(n_1679),
    .Y(n_18480));
 AOI22xp33_ASAP7_75t_SL g172868 (.A1(n_10026),
    .A2(n_64818),
    .B1(\u8_mem[3] [12]),
    .B2(n_70622),
    .Y(n_18491));
 OA22x2_ASAP7_75t_SL g172898 (.A1(n_26819),
    .A2(n_330),
    .B1(n_26823),
    .B2(n_17606),
    .Y(n_18524));
 AOI22xp5_ASAP7_75t_SL g172949 (.A1(n_46478),
    .A2(n_61243),
    .B1(\u10_mem[0] [11]),
    .B2(n_46477),
    .Y(n_18591));
 AND2x4_ASAP7_75t_SL g173 (.A(n_48675),
    .B(n_12142),
    .Y(n_15143));
 NAND2xp5_ASAP7_75t_SL g173001 (.A(n_18652),
    .B(n_18654),
    .Y(n_18655));
 INVxp67_ASAP7_75t_R g173002 (.A(n_4390),
    .Y(n_18652));
 XOR2xp5_ASAP7_75t_SL g173003 (.A(n_28852),
    .B(n_18653),
    .Y(n_18654));
 INVx1_ASAP7_75t_R g173004 (.A(n_366),
    .Y(n_18653));
 NAND3xp33_ASAP7_75t_SL g173006 (.A(n_2124),
    .B(n_31834),
    .C(n_18658),
    .Y(n_18660));
 INVxp67_ASAP7_75t_SL g173007 (.A(n_2164),
    .Y(n_18658));
 NAND3xp33_ASAP7_75t_SL g173013 (.A(n_38705),
    .B(n_18667),
    .C(n_18666),
    .Y(n_18668));
 INVxp67_ASAP7_75t_SL g173014 (.A(n_37340),
    .Y(n_18666));
 AOI22xp33_ASAP7_75t_L g173015 (.A1(n_2458),
    .A2(n_24742),
    .B1(n_1113),
    .B2(n_24741),
    .Y(n_18667));
 INVx1_ASAP7_75t_SL g173024 (.A(n_29688),
    .Y(n_18679));
 NAND2xp5_ASAP7_75t_SL g173027 (.A(n_18683),
    .B(n_742),
    .Y(n_18684));
 AOI22xp5_ASAP7_75t_SL g173028 (.A1(n_58959),
    .A2(\u4_mem[0] [1]),
    .B1(\u4_mem[2] [1]),
    .B2(n_35632),
    .Y(n_18683));
 NAND2x1_ASAP7_75t_SL g173047 (.A(n_56846),
    .B(n_1153),
    .Y(n_18704));
 NAND2x1_ASAP7_75t_SL g173050 (.A(n_18066),
    .B(n_18706),
    .Y(n_18707));
 NAND2xp5_ASAP7_75t_L g173051 (.A(n_24336),
    .B(u10_din_tmp1[9]),
    .Y(n_18706));
 NAND2x1_ASAP7_75t_SL g173053 (.A(n_7417),
    .B(n_1241),
    .Y(n_18709));
 NAND4xp25_ASAP7_75t_SL g173054 (.A(n_2174),
    .B(n_18710),
    .C(n_1745),
    .D(n_1779),
    .Y(n_18711));
 NAND2xp5_ASAP7_75t_SL g173055 (.A(n_18709),
    .B(n_47551),
    .Y(n_18710));
 NOR2xp33_ASAP7_75t_SL g173086 (.A(n_20673),
    .B(n_77796),
    .Y(n_18742));
 NAND2xp5_ASAP7_75t_SL g173089 (.A(n_77796),
    .B(u6_rp[0]),
    .Y(n_18745));
 AOI221xp5_ASAP7_75t_SL g173186 (.A1(n_24513),
    .A2(\u3_mem[1] [20]),
    .B1(n_24512),
    .B2(\u3_mem[0] [20]),
    .C(n_1784),
    .Y(n_18841));
 OR2x2_ASAP7_75t_SL g173202 (.A(dma_ack_i[3]),
    .B(n_2517),
    .Y(n_18857));
 AO21x1_ASAP7_75t_SL g173212 (.A1(n_15025),
    .A2(n_15024),
    .B(n_34534),
    .Y(n_18871));
 INVx1_ASAP7_75t_SL g173213 (.A(n_18872),
    .Y(n_18873));
 OAI21xp5_ASAP7_75t_SL g173214 (.A1(n_2371),
    .A2(n_2544),
    .B(n_15032),
    .Y(n_18872));
 AO21x1_ASAP7_75t_SL g173216 (.A1(n_30060),
    .A2(n_30059),
    .B(n_30061),
    .Y(n_18875));
 NOR2xp33_ASAP7_75t_SL g173226 (.A(n_1661),
    .B(u12_we2),
    .Y(n_18885));
 NAND3xp33_ASAP7_75t_L g173227 (.A(wb_stb_i),
    .B(wb_we_i),
    .C(wb_cyc_i),
    .Y(n_18886));
 OR3x1_ASAP7_75t_R g173228 (.A(wb_addr_i[30]),
    .B(wb_addr_i[31]),
    .C(wb_addr_i[29]),
    .Y(n_18887));
 OR2x2_ASAP7_75t_SL g173229 (.A(n_18885),
    .B(n_18888),
    .Y(n_18889));
 OR2x2_ASAP7_75t_L g173230 (.A(n_18886),
    .B(n_18887),
    .Y(n_18888));
 AO22x2_ASAP7_75t_SL g173237 (.A1(n_69795),
    .A2(n_18895),
    .B1(n_24742),
    .B2(n_18894),
    .Y(n_18896));
 INVxp33_ASAP7_75t_R g173250 (.A(in_valid_s1[2]),
    .Y(n_18928));
 HB1xp67_ASAP7_75t_SL g173253 (.A(in_valid_s[2]),
    .Y(n_18931));
 HB1xp67_ASAP7_75t_SL g173254 (.A(in_valid_s[2]),
    .Y(n_18933));
 O2A1O1Ixp33_ASAP7_75t_L g173312 (.A1(o6_status[0]),
    .A2(oc2_cfg[4]),
    .B(o6_status[1]),
    .C(oc2_cfg[5]),
    .Y(n_19006));
 AOI22xp5_ASAP7_75t_SL g173313 (.A1(n_66026),
    .A2(n_67247),
    .B1(n_19004),
    .B2(n_29621),
    .Y(n_19005));
 HB1xp67_ASAP7_75t_R g173314 (.A(oc2_cfg[4]),
    .Y(n_19004));
 OAI31xp33_ASAP7_75t_SL g173315 (.A1(oc2_cfg[4]),
    .A2(o6_status[1]),
    .A3(o6_status[0]),
    .B(n_2950),
    .Y(n_19007));
 AOI22xp33_ASAP7_75t_L g173316 (.A1(oc2_cfg[4]),
    .A2(n_8212),
    .B1(u13_intm_r[20]),
    .B2(n_7082),
    .Y(n_19008));
 HB1xp67_ASAP7_75t_SL g173339 (.A(u10_wp[1]),
    .Y(n_19045));
 NAND2xp5_ASAP7_75t_SL g173340 (.A(n_47768),
    .B(n_19045),
    .Y(n_19046));
 O2A1O1Ixp33_ASAP7_75t_SL g173357 (.A1(oc0_cfg[4]),
    .A2(o3_status[0]),
    .B(o3_status[1]),
    .C(oc0_cfg[5]),
    .Y(n_19069));
 AOI22xp5_ASAP7_75t_SL g173358 (.A1(n_66868),
    .A2(n_67247),
    .B1(n_19067),
    .B2(n_67248),
    .Y(n_19068));
 HB1xp67_ASAP7_75t_R g173359 (.A(oc0_cfg[5]),
    .Y(n_19067));
 NAND2x1_ASAP7_75t_SL g173416 (.A(out_slt0[12]),
    .B(n_19132),
    .Y(n_19133));
 AOI22xp5_ASAP7_75t_SL g173512 (.A1(n_10684),
    .A2(n_64861),
    .B1(\u6_mem[3] [29]),
    .B2(n_72084),
    .Y(n_19234));
 AOI22xp5_ASAP7_75t_SL g173513 (.A1(n_10660),
    .A2(n_64861),
    .B1(\u6_mem[3] [30]),
    .B2(n_72084),
    .Y(n_19235));
 AOI22xp5_ASAP7_75t_SL g173515 (.A1(n_65900),
    .A2(n_64861),
    .B1(\u6_mem[3] [31]),
    .B2(n_72084),
    .Y(n_19237));
 AOI22xp5_ASAP7_75t_SL g173519 (.A1(n_35437),
    .A2(n_64861),
    .B1(\u6_mem[3] [26]),
    .B2(n_72084),
    .Y(n_19241));
 AND3x1_ASAP7_75t_R g173649 (.A(n_40978),
    .B(n_64816),
    .C(n_15867),
    .Y(n_19378));
 AND3x4_ASAP7_75t_SL g173655 (.A(n_78931),
    .B(o9_we),
    .C(n_64816),
    .Y(n_19383));
 AO22x1_ASAP7_75t_SL g173763 (.A1(\u7_mem[1] [19]),
    .A2(n_49617),
    .B1(\u7_mem[3] [19]),
    .B2(n_49618),
    .Y(n_19495));
 AOI22xp33_ASAP7_75t_SL g173764 (.A1(n_49617),
    .A2(\u7_mem[1] [17]),
    .B1(n_49618),
    .B2(\u7_mem[3] [17]),
    .Y(n_19496));
 AOI22xp33_ASAP7_75t_SL g173765 (.A1(n_49617),
    .A2(\u7_mem[1] [16]),
    .B1(n_49618),
    .B2(\u7_mem[3] [16]),
    .Y(n_19497));
 AOI22xp5_ASAP7_75t_SL g173769 (.A1(n_49617),
    .A2(\u7_mem[1] [3]),
    .B1(\u7_mem[3] [3]),
    .B2(n_49618),
    .Y(n_19501));
 AOI22xp5_ASAP7_75t_SL g173770 (.A1(n_49617),
    .A2(\u7_mem[1] [2]),
    .B1(\u7_mem[3] [2]),
    .B2(n_49618),
    .Y(n_19502));
 AOI22xp5_ASAP7_75t_SL g173771 (.A1(\u7_mem[1] [18]),
    .A2(n_49617),
    .B1(\u7_mem[3] [18]),
    .B2(n_49618),
    .Y(n_19503));
 AOI22xp33_ASAP7_75t_SL g173772 (.A1(\u7_mem[1] [9]),
    .A2(n_49617),
    .B1(\u7_mem[3] [9]),
    .B2(n_49618),
    .Y(n_19504));
 AOI22xp5_ASAP7_75t_SL g173773 (.A1(\u7_mem[1] [10]),
    .A2(n_49617),
    .B1(\u7_mem[3] [10]),
    .B2(n_49618),
    .Y(n_19505));
 AOI22xp5_ASAP7_75t_SL g173774 (.A1(\u7_mem[1] [8]),
    .A2(n_49617),
    .B1(\u7_mem[3] [8]),
    .B2(n_49618),
    .Y(n_19506));
 AOI22xp33_ASAP7_75t_SL g173777 (.A1(n_2691),
    .A2(n_49618),
    .B1(u7_rp[3]),
    .B2(n_19509),
    .Y(n_19510));
 INVxp67_ASAP7_75t_SL g173778 (.A(n_49618),
    .Y(n_19509));
 NAND2x1_ASAP7_75t_SL g173837 (.A(n_19577),
    .B(n_19576),
    .Y(n_19578));
 NOR3xp33_ASAP7_75t_SL g173838 (.A(n_258),
    .B(u2_to_cnt[1]),
    .C(u2_to_cnt[4]),
    .Y(n_19576));
 NOR3xp33_ASAP7_75t_SL g173839 (.A(n_5),
    .B(u2_to_cnt[2]),
    .C(u2_to_cnt[3]),
    .Y(n_19577));
 INVx1_ASAP7_75t_L g173872 (.A(u5_wp[0]),
    .Y(n_19615));
 INVx1_ASAP7_75t_SL g173874 (.A(n_169),
    .Y(n_19617));
 AOI22xp33_ASAP7_75t_L g173875 (.A1(n_13405),
    .A2(n_19619),
    .B1(n_19620),
    .B2(u5_rp[0]),
    .Y(n_19621));
 AOI22xp5_ASAP7_75t_SL g173876 (.A1(n_19616),
    .A2(n_19615),
    .B1(n_7869),
    .B2(n_19617),
    .Y(n_19619));
 INVx1_ASAP7_75t_SL g173878 (.A(n_19619),
    .Y(n_19620));
 AOI31xp33_ASAP7_75t_SL g173879 (.A1(n_14013),
    .A2(n_19622),
    .A3(n_2695),
    .B(oc2_int_set[2]),
    .Y(n_19623));
 HB1xp67_ASAP7_75t_SL g173880 (.A(n_19619),
    .Y(n_19622));
 NAND2xp33_ASAP7_75t_SL g173925 (.A(n_27129),
    .B(n_78810),
    .Y(n_19672));
 AOI22xp33_ASAP7_75t_SL g173927 (.A1(n_77853),
    .A2(\u6_mem[2] [1]),
    .B1(n_41152),
    .B2(\u6_mem[3] [1]),
    .Y(n_19669));
 NAND2xp5_ASAP7_75t_L g173940 (.A(n_28239),
    .B(n_50290),
    .Y(n_19687));
 AOI22xp33_ASAP7_75t_L g174 (.A1(n_8235),
    .A2(i3_dout[8]),
    .B1(n_14933),
    .B2(i6_dout[8]),
    .Y(n_16722));
 AND3x2_ASAP7_75t_SL g174069_dup202286 (.A(n_41910),
    .B(n_48432),
    .C(o3_we),
    .Y(n_52892));
 NAND4xp25_ASAP7_75t_SL g174499 (.A(n_14680),
    .B(n_21696),
    .C(n_24336),
    .D(n_25440),
    .Y(n_20245));
 NAND3xp33_ASAP7_75t_SL g174501 (.A(n_21696),
    .B(n_25440),
    .C(n_14976),
    .Y(n_20246));
 INVxp67_ASAP7_75t_SL g174502 (.A(n_25440),
    .Y(n_20247));
 XNOR2xp5_ASAP7_75t_SL g174550 (.A(n_24588),
    .B(n_20316),
    .Y(n_20317));
 NAND2xp5_ASAP7_75t_L g174551 (.A(n_40417),
    .B(u3_rp[0]),
    .Y(n_20316));
 NOR2xp33_ASAP7_75t_SL g174553 (.A(n_2454),
    .B(n_20317),
    .Y(n_20319));
 AND2x2_ASAP7_75t_SL g174613 (.A(n_7693),
    .B(n_7692),
    .Y(n_20426));
 NAND2xp5_ASAP7_75t_L g174906 (.A(n_695),
    .B(n_71974),
    .Y(n_20759));
 AOI22xp33_ASAP7_75t_SL g174908 (.A1(\u3_mem[0] [19]),
    .A2(n_50341),
    .B1(n_50342),
    .B2(\u3_mem[2] [19]),
    .Y(n_20756));
 NAND2xp5_ASAP7_75t_SL g174910 (.A(n_573),
    .B(n_71974),
    .Y(n_20760));
 NAND2xp5_ASAP7_75t_SL g174933 (.A(n_278),
    .B(n_171),
    .Y(n_20783));
 INVxp33_ASAP7_75t_R g174970 (.A(in_valid_s1[0]),
    .Y(n_20821));
 HB1xp67_ASAP7_75t_SL g174972 (.A(in_valid_s[0]),
    .Y(n_20824));
 AOI221x1_ASAP7_75t_SL g175 (.A1(n_79104),
    .A2(n_47682),
    .B1(n_12519),
    .B2(n_38373),
    .C(n_38367),
    .Y(n_47683));
 NAND2x1_ASAP7_75t_SL g175104 (.A(n_20972),
    .B(n_752),
    .Y(n_20973));
 AOI22xp5_ASAP7_75t_SL g175105 (.A1(n_58959),
    .A2(\u4_mem[0] [8]),
    .B1(\u4_mem[1] [8]),
    .B2(n_50709),
    .Y(n_20972));
 NAND2x1_ASAP7_75t_SL g175146 (.A(n_31892),
    .B(n_56851),
    .Y(n_21015));
 HB1xp67_ASAP7_75t_SL g175148 (.A(n_21024),
    .Y(n_2188));
 INVx1_ASAP7_75t_SL g175149 (.A(n_7671),
    .Y(n_21024));
 AO21x1_ASAP7_75t_L g175150 (.A1(n_56859),
    .A2(n_13755),
    .B(n_21026),
    .Y(n_21027));
 INVxp67_ASAP7_75t_SL g175151 (.A(n_2188),
    .Y(n_21026));
 BUFx6f_ASAP7_75t_SL g175200 (.A(n_6141),
    .Y(n_21076));
 INVx2_ASAP7_75t_SL g175201 (.A(n_21076),
    .Y(n_12097));
 AND2x4_ASAP7_75t_SL g175212 (.A(u10_rp[1]),
    .B(u10_rp[0]),
    .Y(n_21092));
 AOI22xp33_ASAP7_75t_SL g175213 (.A1(n_14821),
    .A2(\u10_mem[2] [2]),
    .B1(n_21093),
    .B2(\u10_mem[3] [2]),
    .Y(n_21094));
 BUFx12f_ASAP7_75t_SL g175214 (.A(n_21092),
    .Y(n_21093));
 AOI22xp33_ASAP7_75t_SL g175215 (.A1(n_14821),
    .A2(\u10_mem[2] [26]),
    .B1(n_21093),
    .B2(\u10_mem[3] [26]),
    .Y(n_21095));
 AOI22xp33_ASAP7_75t_SL g175216 (.A1(n_14821),
    .A2(\u10_mem[2] [3]),
    .B1(n_21093),
    .B2(\u10_mem[3] [3]),
    .Y(n_21096));
 AOI22xp33_ASAP7_75t_SL g175217 (.A1(n_14821),
    .A2(\u10_mem[2] [8]),
    .B1(n_21093),
    .B2(\u10_mem[3] [8]),
    .Y(n_21097));
 AOI22xp33_ASAP7_75t_SL g175218 (.A1(n_14821),
    .A2(\u10_mem[2] [12]),
    .B1(n_21093),
    .B2(\u10_mem[3] [12]),
    .Y(n_21098));
 AOI22xp33_ASAP7_75t_SL g175219 (.A1(n_14821),
    .A2(\u10_mem[2] [16]),
    .B1(n_21093),
    .B2(\u10_mem[3] [16]),
    .Y(n_21099));
 AOI22xp33_ASAP7_75t_SL g175220 (.A1(n_14821),
    .A2(\u10_mem[2] [22]),
    .B1(n_21093),
    .B2(\u10_mem[3] [22]),
    .Y(n_21100));
 AOI22xp33_ASAP7_75t_SL g175221 (.A1(n_14821),
    .A2(\u10_mem[2] [31]),
    .B1(n_21093),
    .B2(\u10_mem[3] [31]),
    .Y(n_21101));
 AOI22xp33_ASAP7_75t_SL g175222 (.A1(n_14821),
    .A2(\u10_mem[2] [10]),
    .B1(n_21093),
    .B2(\u10_mem[3] [10]),
    .Y(n_21102));
 AOI22xp33_ASAP7_75t_SL g175223 (.A1(n_14821),
    .A2(\u10_mem[2] [0]),
    .B1(n_21093),
    .B2(\u10_mem[3] [0]),
    .Y(n_21103));
 AOI22xp5_ASAP7_75t_SL g175224 (.A1(n_14821),
    .A2(\u10_mem[2] [19]),
    .B1(n_21093),
    .B2(\u10_mem[3] [19]),
    .Y(n_21104));
 AOI22xp5_ASAP7_75t_SL g175225 (.A1(n_14821),
    .A2(\u10_mem[2] [18]),
    .B1(n_21093),
    .B2(\u10_mem[3] [18]),
    .Y(n_21105));
 AOI22xp5_ASAP7_75t_SL g175226 (.A1(n_14821),
    .A2(\u10_mem[2] [28]),
    .B1(n_21093),
    .B2(\u10_mem[3] [28]),
    .Y(n_21106));
 AOI22xp5_ASAP7_75t_SL g175227 (.A1(n_14821),
    .A2(\u10_mem[2] [1]),
    .B1(n_21093),
    .B2(\u10_mem[3] [1]),
    .Y(n_21107));
 AOI22xp5_ASAP7_75t_SL g175228 (.A1(n_14821),
    .A2(\u10_mem[2] [4]),
    .B1(n_21093),
    .B2(\u10_mem[3] [4]),
    .Y(n_21108));
 AOI22xp5_ASAP7_75t_SL g175229 (.A1(n_14821),
    .A2(\u10_mem[2] [5]),
    .B1(n_21093),
    .B2(\u10_mem[3] [5]),
    .Y(n_21109));
 AOI22xp5_ASAP7_75t_SL g175230 (.A1(n_14821),
    .A2(\u10_mem[2] [6]),
    .B1(n_21093),
    .B2(\u10_mem[3] [6]),
    .Y(n_21110));
 AOI22xp5_ASAP7_75t_SL g175231 (.A1(n_14821),
    .A2(\u10_mem[2] [7]),
    .B1(n_21093),
    .B2(\u10_mem[3] [7]),
    .Y(n_21111));
 AOI22xp5_ASAP7_75t_SL g175232 (.A1(n_14821),
    .A2(\u10_mem[2] [9]),
    .B1(n_21093),
    .B2(\u10_mem[3] [9]),
    .Y(n_21112));
 AOI22xp5_ASAP7_75t_SL g175233 (.A1(n_14821),
    .A2(\u10_mem[2] [13]),
    .B1(n_21093),
    .B2(\u10_mem[3] [13]),
    .Y(n_21113));
 AOI22xp5_ASAP7_75t_SL g175234 (.A1(n_14821),
    .A2(\u10_mem[2] [15]),
    .B1(n_21093),
    .B2(\u10_mem[3] [15]),
    .Y(n_21114));
 AOI22xp5_ASAP7_75t_SL g175235 (.A1(n_14821),
    .A2(\u10_mem[2] [17]),
    .B1(n_21093),
    .B2(\u10_mem[3] [17]),
    .Y(n_21115));
 AOI22xp5_ASAP7_75t_SL g175236 (.A1(n_14821),
    .A2(\u10_mem[2] [20]),
    .B1(n_21093),
    .B2(\u10_mem[3] [20]),
    .Y(n_21116));
 AOI22xp5_ASAP7_75t_SL g175237 (.A1(n_14821),
    .A2(\u10_mem[2] [21]),
    .B1(n_21093),
    .B2(\u10_mem[3] [21]),
    .Y(n_21117));
 AOI22xp5_ASAP7_75t_SL g175238 (.A1(n_14821),
    .A2(\u10_mem[2] [27]),
    .B1(n_21093),
    .B2(\u10_mem[3] [27]),
    .Y(n_21118));
 AOI22xp5_ASAP7_75t_SL g175239 (.A1(n_14821),
    .A2(\u10_mem[2] [30]),
    .B1(n_21093),
    .B2(\u10_mem[3] [30]),
    .Y(n_21119));
 AOI22xp33_ASAP7_75t_SL g175240 (.A1(n_14821),
    .A2(\u10_mem[2] [29]),
    .B1(n_21093),
    .B2(\u10_mem[3] [29]),
    .Y(n_21120));
 AOI22xp5_ASAP7_75t_SL g175241 (.A1(n_14821),
    .A2(\u10_mem[2] [25]),
    .B1(n_21093),
    .B2(\u10_mem[3] [25]),
    .Y(n_21121));
 AOI22xp33_ASAP7_75t_SL g175242 (.A1(n_14821),
    .A2(\u10_mem[2] [11]),
    .B1(n_21093),
    .B2(\u10_mem[3] [11]),
    .Y(n_21122));
 AOI22xp5_ASAP7_75t_SL g175243 (.A1(n_14821),
    .A2(\u10_mem[2] [24]),
    .B1(n_21093),
    .B2(\u10_mem[3] [24]),
    .Y(n_21123));
 AOI22xp33_ASAP7_75t_SL g175244 (.A1(n_14821),
    .A2(\u10_mem[2] [14]),
    .B1(n_21093),
    .B2(\u10_mem[3] [14]),
    .Y(n_21124));
 NAND2xp5_ASAP7_75t_L g175263 (.A(n_49617),
    .B(\u7_mem[1] [4]),
    .Y(n_21141));
 O2A1O1Ixp33_ASAP7_75t_SL g175268 (.A1(i4_re),
    .A2(n_25439),
    .B(n_21147),
    .C(n_29934),
    .Y(n_21148));
 NAND2xp33_ASAP7_75t_SL g175269 (.A(n_25439),
    .B(i4_re),
    .Y(n_21147));
 OR2x2_ASAP7_75t_SL g175310 (.A(n_14763),
    .B(n_78135),
    .Y(n_21190));
 OAI22xp5_ASAP7_75t_SL g175346 (.A1(n_18931),
    .A2(u14_u8_en_out_l_44),
    .B1(in_slt0[9]),
    .B2(n_2640),
    .Y(n_21225));
 AND3x1_ASAP7_75t_SL g175347 (.A(n_7695),
    .B(in_valid_s[2]),
    .C(u14_u8_en_out_l_44),
    .Y(n_21226));
 NOR2xp33_ASAP7_75t_SL g175352 (.A(n_24594),
    .B(n_21507),
    .Y(n_21234));
 AND2x4_ASAP7_75t_SL g175375 (.A(n_710),
    .B(n_17399),
    .Y(n_21261));
 AOI22xp5_ASAP7_75t_SL g175414 (.A1(n_10924),
    .A2(n_21311),
    .B1(n_549),
    .B2(n_26541),
    .Y(n_21312));
 NOR2x1p5_ASAP7_75t_SL g175415 (.A(n_21332),
    .B(n_21335),
    .Y(n_21311));
 OAI221xp5_ASAP7_75t_SL g175420 (.A1(n_1679),
    .A2(n_21638),
    .B1(n_1705),
    .B2(n_21646),
    .C(n_13249),
    .Y(n_21317));
 OAI221xp5_ASAP7_75t_SL g175424 (.A1(n_1679),
    .A2(n_21709),
    .B1(n_1705),
    .B2(n_21638),
    .C(n_13244),
    .Y(n_21321));
 OAI221xp5_ASAP7_75t_SL g175428 (.A1(n_1679),
    .A2(n_1707),
    .B1(n_1705),
    .B2(n_14313),
    .C(n_13246),
    .Y(n_21325));
 INVx3_ASAP7_75t_SL g175436 (.A(wb_addr_i[2]),
    .Y(n_21331));
 NAND2x1p5_ASAP7_75t_SL g175437 (.A(wb_addr_i[3]),
    .B(rf_we),
    .Y(n_21335));
 AND3x1_ASAP7_75t_SL g175440 (.A(n_21342),
    .B(n_36068),
    .C(n_47740),
    .Y(n_21343));
 INVx1_ASAP7_75t_SL g175441 (.A(n_21341),
    .Y(n_21342));
 NAND2x1_ASAP7_75t_SL g175442 (.A(out_slt0[6]),
    .B(n_67329),
    .Y(n_21341));
 NAND2xp5_ASAP7_75t_SL g175581 (.A(n_43082),
    .B(u15_valid_r),
    .Y(n_21513));
 INVxp33_ASAP7_75t_R g175582 (.A(crac_out[31]),
    .Y(n_21514));
 NAND2xp33_ASAP7_75t_SL g175584 (.A(n_21513),
    .B(n_21516),
    .Y(n_21517));
 INVx1_ASAP7_75t_SL g175585 (.A(n_2063),
    .Y(n_21516));
 NAND2xp5_ASAP7_75t_R g175586 (.A(n_21516),
    .B(n_23),
    .Y(n_21518));
 INVxp67_ASAP7_75t_SL g175588 (.A(n_21520),
    .Y(n_21521));
 INVx2_ASAP7_75t_SL g175589 (.A(n_12143),
    .Y(n_21520));
 INVxp67_ASAP7_75t_R g175593 (.A(\u3_mem[3] [21]),
    .Y(n_8));
 AND2x4_ASAP7_75t_SL g175594 (.A(n_48428),
    .B(n_21520),
    .Y(n_21527));
 OAI221xp5_ASAP7_75t_SL g175597 (.A1(n_24883),
    .A2(n_1714),
    .B1(n_48057),
    .B2(n_1820),
    .C(n_48636),
    .Y(n_21530));
 OAI221xp5_ASAP7_75t_SL g175601 (.A1(n_24883),
    .A2(n_24886),
    .B1(n_48057),
    .B2(n_48053),
    .C(n_48635),
    .Y(n_21534));
 OAI22xp5_ASAP7_75t_SL g175604 (.A1(n_21538),
    .A2(n_21539),
    .B1(n_27257),
    .B2(n_21540),
    .Y(n_21541));
 INVx1_ASAP7_75t_SL g175605 (.A(n_27257),
    .Y(n_21538));
 NAND2xp5_ASAP7_75t_L g175607 (.A(u11_rp[0]),
    .B(n_28954),
    .Y(n_21539));
 INVxp67_ASAP7_75t_R g175608 (.A(n_21539),
    .Y(n_21540));
 INVxp67_ASAP7_75t_SL g175610 (.A(n_21520),
    .Y(n_21543));
 INVxp33_ASAP7_75t_R g175614 (.A(\u3_mem[3] [17]),
    .Y(n_21546));
 AND2x4_ASAP7_75t_SL g175615 (.A(n_48428),
    .B(n_21520),
    .Y(n_21549));
 OR2x6_ASAP7_75t_SL g175616 (.A(n_48427),
    .B(n_12143),
    .Y(n_21550));
 OAI21xp5_ASAP7_75t_SL g175618 (.A1(n_1707),
    .A2(n_10937),
    .B(n_744),
    .Y(n_21552));
 XNOR2xp5_ASAP7_75t_SL g175646 (.A(n_13829),
    .B(n_13827),
    .Y(n_21599));
 INVx1_ASAP7_75t_SL g175647 (.A(n_13827),
    .Y(n_21600));
 INVx1_ASAP7_75t_L g175677 (.A(in_slt6[9]),
    .Y(n_21631));
 INVx1_ASAP7_75t_L g175684 (.A(in_slt6[10]),
    .Y(n_21638));
 INVx1_ASAP7_75t_L g175692 (.A(in_slt6[12]),
    .Y(n_21646));
 INVx1_ASAP7_75t_R g175711 (.A(in_slt3[5]),
    .Y(n_21665));
 INVx1_ASAP7_75t_L g175715 (.A(in_slt4[14]),
    .Y(n_21669));
 INVx1_ASAP7_75t_R g175719 (.A(in_slt3[16]),
    .Y(n_21673));
 XNOR2xp5_ASAP7_75t_SL g175741 (.A(n_13857),
    .B(n_13855),
    .Y(n_21695));
 INVx1_ASAP7_75t_SL g175742 (.A(n_13855),
    .Y(n_21696));
 INVx1_ASAP7_75t_R g175743 (.A(in_slt6[17]),
    .Y(n_21697));
 INVx1_ASAP7_75t_R g175751 (.A(in_slt6[15]),
    .Y(n_21705));
 INVx1_ASAP7_75t_L g175755 (.A(in_slt6[8]),
    .Y(n_21709));
 AND3x1_ASAP7_75t_SL g175809 (.A(n_184),
    .B(n_24764),
    .C(u26_cnt[2]),
    .Y(n_21776));
 NOR4xp25_ASAP7_75t_L g175810 (.A(n_21777),
    .B(n_339),
    .C(n_15056),
    .D(u26_cnt[2]),
    .Y(n_21778));
 OR3x1_ASAP7_75t_SL g175811 (.A(n_31535),
    .B(n_21776),
    .C(ac97_rst_force),
    .Y(n_21777));
 NOR4xp25_ASAP7_75t_SL g175813 (.A(n_550),
    .B(n_31535),
    .C(n_21776),
    .D(ac97_rst_force),
    .Y(n_21780));
 INVxp67_ASAP7_75t_R g175814 (.A(n_339),
    .Y(n_550));
 INVxp67_ASAP7_75t_SL g175817 (.A(n_21780),
    .Y(n_21784));
 AOI21xp5_ASAP7_75t_SL g175819 (.A1(n_21793),
    .A2(n_29314),
    .B(n_21794),
    .Y(n_21795));
 XNOR2xp5_ASAP7_75t_SL g175821 (.A(u3_rp[3]),
    .B(n_616),
    .Y(n_21793));
 OAI22xp33_ASAP7_75t_SL g175822 (.A1(n_34541),
    .A2(n_2687),
    .B1(n_4261),
    .B2(n_908),
    .Y(n_21794));
 AOI21xp5_ASAP7_75t_SL g175892 (.A1(n_63999),
    .A2(n_550),
    .B(n_21780),
    .Y(n_21865));
 A2O1A1Ixp33_ASAP7_75t_SL g175895 (.A1(n_303),
    .A2(n_50090),
    .B(n_14947),
    .C(n_63999),
    .Y(n_21867));
 OAI21xp5_ASAP7_75t_SL g175898 (.A1(n_719),
    .A2(n_720),
    .B(n_63999),
    .Y(n_21871));
 OAI21xp5_ASAP7_75t_SL g175899 (.A1(n_47539),
    .A2(n_1292),
    .B(n_63999),
    .Y(n_21872));
 INVxp67_ASAP7_75t_L g175901 (.A(n_63999),
    .Y(n_21874));
 AOI22xp33_ASAP7_75t_SL g175904 (.A1(u8_rp[3]),
    .A2(n_13980),
    .B1(n_2689),
    .B2(n_78273),
    .Y(n_21876));
 INVx1_ASAP7_75t_L g175906 (.A(in_slt4[13]),
    .Y(n_21878));
 AOI22xp33_ASAP7_75t_SL g175956 (.A1(n_46478),
    .A2(n_65879),
    .B1(\u10_mem[0] [6]),
    .B2(n_46477),
    .Y(n_21938));
 AOI22xp33_ASAP7_75t_SL g175968 (.A1(n_31786),
    .A2(n_46478),
    .B1(\u10_mem[0] [8]),
    .B2(n_46477),
    .Y(n_21947));
 AOI21xp5_ASAP7_75t_SL g176 (.A1(n_43604),
    .A2(n_43605),
    .B(n_43606),
    .Y(n_43607));
 NAND2xp5_ASAP7_75t_L g176012 (.A(n_20973),
    .B(n_24350),
    .Y(n_21996));
 INVxp67_ASAP7_75t_SL g176040 (.A(n_10870),
    .Y(n_22025));
 AND2x4_ASAP7_75t_SL g176041_dup (.A(n_33774),
    .B(n_30452),
    .Y(n_25387));
 NAND4xp25_ASAP7_75t_SL g176064 (.A(n_2108),
    .B(n_1999),
    .C(n_22059),
    .D(n_1418),
    .Y(n_22060));
 AOI22xp33_ASAP7_75t_L g176065 (.A1(n_79305),
    .A2(\u6_mem[0] [22]),
    .B1(\u6_mem[2] [22]),
    .B2(n_79306),
    .Y(n_22059));
 AND2x2_ASAP7_75t_SL g176067 (.A(n_695),
    .B(n_71972),
    .Y(n_22062));
 OAI211xp5_ASAP7_75t_SL g176068 (.A1(n_2524),
    .A2(n_66198),
    .B(n_27341),
    .C(n_2238),
    .Y(n_22064));
 NOR2xp33_ASAP7_75t_SL g176147 (.A(n_2596),
    .B(n_5748),
    .Y(n_22163));
 OAI21xp33_ASAP7_75t_SL g176152 (.A1(u13_ints_r[12]),
    .A2(oc3_int_set[1]),
    .B(n_22174),
    .Y(n_22175));
 OR2x2_ASAP7_75t_SL g176153 (.A(n_26255),
    .B(n_22267),
    .Y(n_22174));
 OAI21xp33_ASAP7_75t_SL g176154 (.A1(u13_ints_r[22]),
    .A2(ic0_int_set[2]),
    .B(n_22174),
    .Y(n_22176));
 OAI21xp33_ASAP7_75t_SL g176155 (.A1(u13_ints_r[15]),
    .A2(oc4_int_set[1]),
    .B(n_22174),
    .Y(n_22177));
 OAI21xp33_ASAP7_75t_SL g176156 (.A1(u13_ints_r[13]),
    .A2(oc3_int_set[2]),
    .B(n_22174),
    .Y(n_22178));
 OAI21xp33_ASAP7_75t_SL g176157 (.A1(u13_ints_r[0]),
    .A2(n_42736),
    .B(n_22174),
    .Y(n_22179));
 OAI21xp33_ASAP7_75t_SL g176158 (.A1(n_2038),
    .A2(oc0_int_set[1]),
    .B(n_22174),
    .Y(n_22180));
 OAI21xp33_ASAP7_75t_SL g176159 (.A1(n_2036),
    .A2(oc0_int_set[2]),
    .B(n_22174),
    .Y(n_22181));
 OAI21xp33_ASAP7_75t_SL g176160 (.A1(n_2034),
    .A2(oc1_int_set[1]),
    .B(n_22174),
    .Y(n_22182));
 OAI21xp33_ASAP7_75t_SL g176161 (.A1(u13_ints_r[7]),
    .A2(oc1_int_set[2]),
    .B(n_22183),
    .Y(n_22184));
 OAI21xp33_ASAP7_75t_SL g176162 (.A1(n_2031),
    .A2(oc2_int_set[1]),
    .B(n_22183),
    .Y(n_22185));
 OAI21xp33_ASAP7_75t_SL g176163 (.A1(n_2029),
    .A2(oc2_int_set[2]),
    .B(n_22183),
    .Y(n_22186));
 OAI21xp33_ASAP7_75t_SL g176164 (.A1(u13_ints_r[16]),
    .A2(oc4_int_set[2]),
    .B(n_22183),
    .Y(n_22187));
 OAI21xp33_ASAP7_75t_SL g176165 (.A1(u13_ints_r[19]),
    .A2(oc5_int_set[2]),
    .B(n_22183),
    .Y(n_22188));
 OAI21xp33_ASAP7_75t_SL g176166 (.A1(n_2024),
    .A2(ic1_int_set[1]),
    .B(n_22183),
    .Y(n_22189));
 OAI21xp33_ASAP7_75t_SL g176167 (.A1(u13_ints_r[25]),
    .A2(ic1_int_set[2]),
    .B(n_22183),
    .Y(n_22190));
 NAND4xp25_ASAP7_75t_SL g176214 (.A(n_50291),
    .B(n_22247),
    .C(n_22248),
    .D(n_53372),
    .Y(n_22250));
 NAND2xp5_ASAP7_75t_SL g176215 (.A(n_34645),
    .B(n_50290),
    .Y(n_22247));
 AOI22xp33_ASAP7_75t_SL g176216 (.A1(\u7_mem[0] [30]),
    .A2(n_65055),
    .B1(n_65056),
    .B2(\u7_mem[1] [30]),
    .Y(n_22248));
 AOI221xp5_ASAP7_75t_SL g176218 (.A1(n_22256),
    .A2(n_5077),
    .B1(n_4225),
    .B2(out_slt8[15]),
    .C(n_4453),
    .Y(n_22257));
 NAND4xp25_ASAP7_75t_SL g176219 (.A(n_22252),
    .B(n_22253),
    .C(n_22254),
    .D(n_53371),
    .Y(n_22256));
 NAND2xp5_ASAP7_75t_SL g176220 (.A(n_41491),
    .B(n_666),
    .Y(n_22252));
 NAND2xp5_ASAP7_75t_SL g176221 (.A(n_49620),
    .B(n_50290),
    .Y(n_22253));
 AOI22xp33_ASAP7_75t_L g176222 (.A1(\u7_mem[0] [27]),
    .A2(n_65055),
    .B1(\u7_mem[1] [27]),
    .B2(n_65056),
    .Y(n_22254));
 NAND4xp75_ASAP7_75t_SL g176228 (.A(n_8220),
    .B(n_8311),
    .C(wb_addr_i[4]),
    .D(wb_addr_i[3]),
    .Y(n_22267));
 NAND3xp33_ASAP7_75t_SL g176229 (.A(n_21517),
    .B(n_22268),
    .C(n_21518),
    .Y(n_22269));
 OAI21xp33_ASAP7_75t_SL g176237 (.A1(ic1_int_set[0]),
    .A2(n_2678),
    .B(n_22276),
    .Y(n_22277));
 OAI21xp33_ASAP7_75t_SL g176238 (.A1(ic0_int_set[0]),
    .A2(u13_ints_r[20]),
    .B(n_22276),
    .Y(n_22278));
 OAI21xp33_ASAP7_75t_SL g176239 (.A1(ic2_int_set[0]),
    .A2(n_219),
    .B(n_22276),
    .Y(n_22279));
 OAI21xp33_ASAP7_75t_SL g176240 (.A1(n_2048),
    .A2(oc5_int_set[1]),
    .B(n_22276),
    .Y(n_22280));
 OAI21xp33_ASAP7_75t_SL g176241 (.A1(u13_ints_r[27]),
    .A2(ic2_int_set[1]),
    .B(n_22276),
    .Y(n_22281));
 OAI21xp33_ASAP7_75t_SL g176242 (.A1(u13_ints_r[21]),
    .A2(ic0_int_set[1]),
    .B(n_22276),
    .Y(n_22282));
 OAI21xp33_ASAP7_75t_SL g176243 (.A1(u13_ints_r[28]),
    .A2(ic2_int_set[2]),
    .B(n_22276),
    .Y(n_22283));
 AOI22xp5_ASAP7_75t_SL g176265 (.A1(n_22577),
    .A2(\u3_mem[1] [6]),
    .B1(n_32644),
    .B2(n_16009),
    .Y(n_22311));
 AOI22xp5_ASAP7_75t_SL g176269 (.A1(n_65949),
    .A2(n_64861),
    .B1(\u6_mem[3] [16]),
    .B2(n_77233),
    .Y(n_22315));
 AOI22xp5_ASAP7_75t_SL g176310 (.A1(n_22505),
    .A2(\u3_mem[1] [29]),
    .B1(n_22715),
    .B2(n_15143),
    .Y(n_22371));
 OR2x6_ASAP7_75t_SL g176333 (.A(n_47787),
    .B(n_18964),
    .Y(n_22396));
 AOI22xp5_ASAP7_75t_SL g176342 (.A1(\u9_mem[3] [23]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25673),
    .Y(n_22407));
 AOI22xp5_ASAP7_75t_SL g176348 (.A1(\u9_mem[3] [24]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25674),
    .Y(n_22413));
 AOI22xp5_ASAP7_75t_SL g176350 (.A1(\u9_mem[3] [28]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25682),
    .Y(n_22415));
 AOI22xp5_ASAP7_75t_SL g176359 (.A1(\u9_mem[3] [29]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25679),
    .Y(n_22424));
 AOI22xp5_ASAP7_75t_SL g176365 (.A1(\u9_mem[3] [31]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25681),
    .Y(n_22430));
 AOI22xp5_ASAP7_75t_SL g176367 (.A1(\u9_mem[3] [1]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_12482),
    .Y(n_22432));
 AOI22xp5_ASAP7_75t_SL g176413 (.A1(\u9_mem[3] [30]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_25680),
    .Y(n_22482));
 AOI22xp33_ASAP7_75t_SL g176436 (.A1(n_22505),
    .A2(\u3_mem[1] [30]),
    .B1(n_10640),
    .B2(n_15143),
    .Y(n_22506));
 INVx4_ASAP7_75t_SL g176437 (.A(n_13176),
    .Y(n_22505));
 AOI22xp5_ASAP7_75t_SL g176438 (.A1(n_75733),
    .A2(n_64819),
    .B1(\u8_mem[3] [0]),
    .B2(n_70622),
    .Y(n_22508));
 AOI22xp33_ASAP7_75t_L g176460 (.A1(n_19593),
    .A2(n_37200),
    .B1(n_7863),
    .B2(n_698),
    .Y(n_22530));
 AOI22xp5_ASAP7_75t_SL g176500 (.A1(n_22577),
    .A2(\u3_mem[1] [3]),
    .B1(n_15867),
    .B2(n_16009),
    .Y(n_22578));
 INVx4_ASAP7_75t_SL g176501 (.A(n_13176),
    .Y(n_22577));
 OAI221xp5_ASAP7_75t_SL g176529 (.A1(n_21665),
    .A2(n_50452),
    .B1(n_48057),
    .B2(n_14301),
    .C(n_48634),
    .Y(n_22632));
 AOI22xp5_ASAP7_75t_SL g176537 (.A1(n_22640),
    .A2(n_64861),
    .B1(\u6_mem[3] [28]),
    .B2(n_72084),
    .Y(n_22642));
 INVx3_ASAP7_75t_SL g176538 (.A(n_10356),
    .Y(n_22640));
 AOI22xp5_ASAP7_75t_SL g176607 (.A1(n_22715),
    .A2(n_73997),
    .B1(\u8_mem[1] [29]),
    .B2(n_75735),
    .Y(n_22718));
 INVx2_ASAP7_75t_SL g176608 (.A(n_10661),
    .Y(n_22715));
 INVxp33_ASAP7_75t_R g176647 (.A(u15_rdd1),
    .Y(n_22774));
 OAI21xp33_ASAP7_75t_R g176648 (.A1(u15_valid_r),
    .A2(u15_rdd1),
    .B(u15_crac_rd),
    .Y(n_22775));
 NOR2xp33_ASAP7_75t_SL g176660 (.A(n_22827),
    .B(n_22828),
    .Y(n_22829));
 NOR2xp33_ASAP7_75t_L g176661 (.A(n_5849),
    .B(n_4496),
    .Y(n_22827));
 OAI22xp33_ASAP7_75t_SL g176662 (.A1(n_43090),
    .A2(n_65325),
    .B1(n_28122),
    .B2(n_24641),
    .Y(n_22828));
 NOR3xp33_ASAP7_75t_SL g176667 (.A(n_47541),
    .B(n_22835),
    .C(n_24725),
    .Y(n_22837));
 INVxp33_ASAP7_75t_SL g176669 (.A(n_19013),
    .Y(n_22835));
 INVx1_ASAP7_75t_SL g176672 (.A(n_37355),
    .Y(n_22839));
 INVxp33_ASAP7_75t_SL g176676 (.A(n_73154),
    .Y(n_22841));
 NAND4xp25_ASAP7_75t_SL g176677 (.A(n_22844),
    .B(n_10629),
    .C(n_7152),
    .D(n_22845),
    .Y(n_22846));
 INVxp67_ASAP7_75t_SL g176678 (.A(n_26803),
    .Y(n_22844));
 NAND2xp5_ASAP7_75t_L g176679 (.A(i3_dout[11]),
    .B(n_8341),
    .Y(n_22845));
 AOI22xp5_ASAP7_75t_SL g176743 (.A1(crac_out[0]),
    .A2(n_28367),
    .B1(n_10924),
    .B2(n_12219),
    .Y(n_22919));
 INVx1_ASAP7_75t_SL g176748 (.A(n_70201),
    .Y(n_22922));
 NOR2xp33_ASAP7_75t_R g176749 (.A(dma_ack_i[5]),
    .B(n_119),
    .Y(n_22923));
 NOR2xp33_ASAP7_75t_R g176756 (.A(dma_ack_i[1]),
    .B(n_131),
    .Y(n_22932));
 INVxp33_ASAP7_75t_R g176761 (.A(n_2227),
    .Y(n_22938));
 AOI22xp5_ASAP7_75t_SL g176786 (.A1(\u9_mem[3] [25]),
    .A2(n_45330),
    .B1(n_24735),
    .B2(n_5173),
    .Y(n_22964));
 AOI22xp33_ASAP7_75t_L g176883 (.A1(\u6_mem[1] [26]),
    .A2(n_48415),
    .B1(\u6_mem[3] [26]),
    .B2(n_17704),
    .Y(n_23079));
 AOI21xp33_ASAP7_75t_SL g176896 (.A1(n_15024),
    .A2(n_15025),
    .B(n_34534),
    .Y(n_23099));
 NOR2xp33_ASAP7_75t_R g176897 (.A(dma_ack_i[0]),
    .B(n_46),
    .Y(n_23100));
 AOI22xp5_ASAP7_75t_SL g176906 (.A1(n_58959),
    .A2(\u4_mem[0] [9]),
    .B1(\u4_mem[2] [9]),
    .B2(n_35632),
    .Y(n_23110));
 NAND2xp5_ASAP7_75t_SL g176922 (.A(n_58960),
    .B(n_1177),
    .Y(n_23129));
 NAND4xp25_ASAP7_75t_SL g176923 (.A(n_7755),
    .B(n_23130),
    .C(n_1757),
    .D(n_1805),
    .Y(n_23131));
 NAND2xp5_ASAP7_75t_SL g176924 (.A(n_23129),
    .B(n_1932),
    .Y(n_23130));
 NAND3xp33_ASAP7_75t_SL g176941 (.A(n_23150),
    .B(n_31754),
    .C(n_31538),
    .Y(n_23154));
 AOI21xp33_ASAP7_75t_SL g176943 (.A1(n_698),
    .A2(n_28691),
    .B(n_19621),
    .Y(n_23150));
 INVxp33_ASAP7_75t_R g177 (.A(wb_data_i[15]),
    .Y(n_65989));
 NAND2xp5_ASAP7_75t_SL g177057 (.A(n_28954),
    .B(n_226),
    .Y(n_23285));
 INVx4_ASAP7_75t_SL g177058 (.A(n_29005),
    .Y(n_23286));
 AOI22xp5_ASAP7_75t_SL g177066 (.A1(n_78274),
    .A2(\u8_mem[1] [11]),
    .B1(\u8_mem[0] [11]),
    .B2(n_59474),
    .Y(n_23296));
 AOI22xp5_ASAP7_75t_SL g177081 (.A1(n_79104),
    .A2(n_23393),
    .B1(n_38371),
    .B2(n_7597),
    .Y(n_23394));
 INVx1_ASAP7_75t_L g177136 (.A(n_2753),
    .Y(n_549));
 INVxp33_ASAP7_75t_R g177137 (.A(n_503),
    .Y(n_23508));
 XNOR2xp5_ASAP7_75t_SL g177158 (.A(n_23526),
    .B(n_50814),
    .Y(n_23529));
 NAND2xp5_ASAP7_75t_L g177159 (.A(n_30078),
    .B(n_36008),
    .Y(n_23530));
 AND2x2_ASAP7_75t_SL g177160 (.A(n_30078),
    .B(n_36008),
    .Y(n_23531));
 OAI21xp33_ASAP7_75t_SL g177279 (.A1(n_23655),
    .A2(n_23656),
    .B(n_23660),
    .Y(n_23661));
 INVx2_ASAP7_75t_L g177280 (.A(n_36528),
    .Y(n_23655));
 INVx1_ASAP7_75t_L g177281 (.A(n_1723),
    .Y(n_23656));
 AOI21xp5_ASAP7_75t_SL g177282 (.A1(n_65293),
    .A2(n_79193),
    .B(n_23659),
    .Y(n_23660));
 AOI21xp33_ASAP7_75t_SL g177284 (.A1(n_51487),
    .A2(n_7544),
    .B(n_57084),
    .Y(n_23659));
 AND2x2_ASAP7_75t_SL g177292 (.A(n_801),
    .B(n_1054),
    .Y(n_23671));
 AOI22xp5_ASAP7_75t_SL g177544 (.A1(n_10194),
    .A2(n_64819),
    .B1(\u8_mem[3] [18]),
    .B2(n_11204),
    .Y(n_23971));
 AND2x2_ASAP7_75t_SL g177835 (.A(u7_wp[0]),
    .B(o8_we),
    .Y(n_24316));
 BUFx6f_ASAP7_75t_SL g177855 (.A(n_684),
    .Y(n_24336));
 NAND2xp5_ASAP7_75t_SL g177857 (.A(n_24336),
    .B(u10_din_tmp1[6]),
    .Y(n_24337));
 AOI22xp5_ASAP7_75t_SL g177859 (.A1(n_8212),
    .A2(n_78041),
    .B1(n_7082),
    .B2(u13_intm_r[27]),
    .Y(n_24341));
 INVx3_ASAP7_75t_SL g177868 (.A(n_8113),
    .Y(n_24350));
 OAI22xp5_ASAP7_75t_SL g177869 (.A1(n_104),
    .A2(n_1762),
    .B1(n_106),
    .B2(n_36011),
    .Y(n_24351));
 NOR5xp2_ASAP7_75t_SL g177886 (.A(n_34540),
    .B(n_24373),
    .C(n_48675),
    .D(n_2748),
    .E(u3_wp[2]),
    .Y(n_24374));
 NOR2xp33_ASAP7_75t_R g177888 (.A(n_40417),
    .B(n_24373),
    .Y(n_24375));
 OAI22xp5_ASAP7_75t_SL g178 (.A1(n_2691),
    .A2(n_42249),
    .B1(n_64103),
    .B2(n_19510),
    .Y(n_43606));
 OAI21xp33_ASAP7_75t_R g178023 (.A1(n_24509),
    .A2(n_1285),
    .B(n_24510),
    .Y(n_24511));
 NAND3xp33_ASAP7_75t_SL g178024 (.A(n_695),
    .B(n_50341),
    .C(\u3_mem[0] [21]),
    .Y(n_24510));
 AND2x4_ASAP7_75t_SL g178025 (.A(n_50341),
    .B(n_695),
    .Y(n_24512));
 INVx2_ASAP7_75t_SL g178026 (.A(n_1285),
    .Y(n_24513));
 AO22x1_ASAP7_75t_SL g178030 (.A1(n_65055),
    .A2(\u7_mem[0] [25]),
    .B1(n_65056),
    .B2(\u7_mem[1] [25]),
    .Y(n_24516));
 INVx1_ASAP7_75t_SL g178037 (.A(n_26183),
    .Y(n_24523));
 INVx1_ASAP7_75t_L g178038 (.A(n_2520),
    .Y(n_24524));
 OAI21xp33_ASAP7_75t_SL g178044 (.A1(n_2373),
    .A2(n_2546),
    .B(n_375),
    .Y(n_24532));
 OAI21xp33_ASAP7_75t_SL g178049 (.A1(n_19006),
    .A2(n_19007),
    .B(n_78094),
    .Y(n_24536));
 NAND2xp5_ASAP7_75t_SL g178060 (.A(n_37142),
    .B(n_31742),
    .Y(n_24553));
 NAND2xp5_ASAP7_75t_SL g178081 (.A(n_50619),
    .B(n_31743),
    .Y(n_24580));
 AND2x2_ASAP7_75t_SL g178098 (.A(n_24594),
    .B(out_slt3[2]),
    .Y(n_24595));
 INVx2_ASAP7_75t_SL g178099 (.A(n_34541),
    .Y(n_24594));
 O2A1O1Ixp33_ASAP7_75t_SL g178124 (.A1(oc3_cfg[4]),
    .A2(o7_status[0]),
    .B(o7_status[1]),
    .C(oc3_cfg[5]),
    .Y(n_24624));
 AOI22xp33_ASAP7_75t_SL g178125 (.A1(n_65919),
    .A2(n_67247),
    .B1(n_24622),
    .B2(n_29621),
    .Y(n_24623));
 HB1xp67_ASAP7_75t_R g178126 (.A(oc3_cfg[4]),
    .Y(n_24622));
 OAI31xp33_ASAP7_75t_SL g178127 (.A1(oc3_cfg[4]),
    .A2(o7_status[0]),
    .A3(o7_status[1]),
    .B(n_2990),
    .Y(n_24625));
 AOI22xp33_ASAP7_75t_SL g178128 (.A1(oc3_cfg[4]),
    .A2(n_8212),
    .B1(u13_intm_r[28]),
    .B2(n_7082),
    .Y(n_24626));
 AND2x2_ASAP7_75t_SL g178129 (.A(o4_we),
    .B(u4_wp[0]),
    .Y(n_24628));
 NOR2xp33_ASAP7_75t_SL g178130 (.A(n_6960),
    .B(n_27061),
    .Y(n_24627));
 INVx1_ASAP7_75t_L g178134 (.A(o4_we),
    .Y(n_24632));
 AND3x4_ASAP7_75t_SL g178135 (.A(n_27057),
    .B(n_48105),
    .C(o4_we),
    .Y(n_24633));
 AOI22xp33_ASAP7_75t_SL g178136 (.A1(n_488),
    .A2(n_24632),
    .B1(n_12275),
    .B2(o4_we),
    .Y(n_24635));
 NAND3xp33_ASAP7_75t_SL g178142 (.A(n_4548),
    .B(n_7766),
    .C(n_26379),
    .Y(n_24641));
 OR2x6_ASAP7_75t_SL g178143 (.A(n_35457),
    .B(n_71392),
    .Y(n_8113));
 AOI22xp5_ASAP7_75t_SL g178167 (.A1(n_24669),
    .A2(n_26541),
    .B1(n_32650),
    .B2(n_15272),
    .Y(n_24670));
 HB1xp67_ASAP7_75t_R g178168 (.A(oc4_cfg[6]),
    .Y(n_24669));
 INVx1_ASAP7_75t_L g178169 (.A(oc4_cfg[6]),
    .Y(n_24672));
 HB1xp67_ASAP7_75t_SL g178193 (.A(u9_wp[1]),
    .Y(n_24730));
 NAND2xp5_ASAP7_75t_SL g178194 (.A(n_13420),
    .B(n_24730),
    .Y(n_24732));
 NAND2x1_ASAP7_75t_SL g178196 (.A(n_21261),
    .B(u9_wp[1]),
    .Y(n_24736));
 INVx4_ASAP7_75t_SL g178197 (.A(u9_wp[1]),
    .Y(n_24737));
 OAI22xp5_ASAP7_75t_SL g178198 (.A1(u9_rp[0]),
    .A2(u9_wp[1]),
    .B1(n_24737),
    .B2(n_13035),
    .Y(n_24738));
 AND3x4_ASAP7_75t_SL g178199 (.A(n_340),
    .B(n_21261),
    .C(u9_wp[1]),
    .Y(n_24739));
 AOI22xp5_ASAP7_75t_SL g178210 (.A1(n_67247),
    .A2(n_65934),
    .B1(n_28689),
    .B2(n_29621),
    .Y(n_24753));
 NOR2xp33_ASAP7_75t_R g178214 (.A(ac97_rst_force),
    .B(u26_cnt[1]),
    .Y(n_24763));
 O2A1O1Ixp33_ASAP7_75t_SL g178215 (.A1(n_21780),
    .A2(n_63999),
    .B(n_24759),
    .C(n_24761),
    .Y(n_24762));
 HB1xp67_ASAP7_75t_SL g178216 (.A(u26_cnt[1]),
    .Y(n_24759));
 NOR3xp33_ASAP7_75t_SL g178217 (.A(n_21777),
    .B(n_339),
    .C(n_24759),
    .Y(n_24761));
 INVx1_ASAP7_75t_SL g178219 (.A(u26_cnt[1]),
    .Y(n_24764));
 AND2x2_ASAP7_75t_SL g178256 (.A(u10_wp[1]),
    .B(n_234),
    .Y(n_24801));
 BUFx3_ASAP7_75t_SL g178258 (.A(u3_wp[1]),
    .Y(n_24804));
 INVx2_ASAP7_75t_SL g178259 (.A(u3_wp[0]),
    .Y(n_24805));
 AOI22xp5_ASAP7_75t_SL g178260 (.A1(n_24806),
    .A2(n_22640),
    .B1(\u3_mem[2] [28]),
    .B2(n_15954),
    .Y(n_24807));
 AND3x4_ASAP7_75t_SL g178261 (.A(n_24805),
    .B(n_24804),
    .C(o3_we),
    .Y(n_24806));
 AOI22xp5_ASAP7_75t_SL g178262 (.A1(n_24806),
    .A2(n_28316),
    .B1(\u3_mem[2] [25]),
    .B2(n_15954),
    .Y(n_24808));
 AOI22xp5_ASAP7_75t_SL g178263 (.A1(n_24806),
    .A2(n_28424),
    .B1(\u3_mem[2] [24]),
    .B2(n_15954),
    .Y(n_24809));
 AOI22xp5_ASAP7_75t_SL g178264 (.A1(n_24806),
    .A2(n_28381),
    .B1(\u3_mem[2] [23]),
    .B2(n_15954),
    .Y(n_24810));
 AOI22xp5_ASAP7_75t_SL g178265 (.A1(n_24806),
    .A2(n_28913),
    .B1(\u3_mem[2] [15]),
    .B2(n_15954),
    .Y(n_24811));
 AOI22xp5_ASAP7_75t_SL g178266 (.A1(n_24806),
    .A2(n_33203),
    .B1(\u3_mem[2] [0]),
    .B2(n_13295),
    .Y(n_24812));
 AOI22xp5_ASAP7_75t_SL g178267 (.A1(n_24806),
    .A2(n_10198),
    .B1(\u3_mem[2] [19]),
    .B2(n_13295),
    .Y(n_24813));
 AOI22xp5_ASAP7_75t_SL g178268 (.A1(n_24806),
    .A2(n_66026),
    .B1(\u3_mem[2] [20]),
    .B2(n_13295),
    .Y(n_24814));
 AOI22xp33_ASAP7_75t_SL g178269 (.A1(n_24806),
    .A2(n_10143),
    .B1(\u3_mem[2] [17]),
    .B2(n_13295),
    .Y(n_24815));
 AOI22xp5_ASAP7_75t_SL g178270 (.A1(n_24806),
    .A2(n_66032),
    .B1(\u3_mem[2] [14]),
    .B2(n_13295),
    .Y(n_24816));
 AOI22xp5_ASAP7_75t_SL g178271 (.A1(n_24806),
    .A2(n_65969),
    .B1(\u3_mem[2] [7]),
    .B2(n_13295),
    .Y(n_24817));
 AOI22xp5_ASAP7_75t_SL g178272 (.A1(n_24806),
    .A2(n_66856),
    .B1(\u3_mem[2] [3]),
    .B2(n_13295),
    .Y(n_24818));
 AOI22xp5_ASAP7_75t_SL g178273 (.A1(n_24806),
    .A2(n_78044),
    .B1(\u3_mem[2] [1]),
    .B2(n_15954),
    .Y(n_24819));
 AOI22xp5_ASAP7_75t_SL g178274 (.A1(n_24806),
    .A2(n_65997),
    .B1(\u3_mem[2] [12]),
    .B2(n_15954),
    .Y(n_24820));
 AOI22xp5_ASAP7_75t_SL g178275 (.A1(n_24806),
    .A2(n_10000),
    .B1(\u3_mem[2] [11]),
    .B2(n_15954),
    .Y(n_24821));
 AOI22xp5_ASAP7_75t_SL g178276 (.A1(n_24806),
    .A2(n_28330),
    .B1(\u3_mem[2] [2]),
    .B2(n_13295),
    .Y(n_24822));
 AOI22xp5_ASAP7_75t_SL g178277 (.A1(n_24806),
    .A2(n_10058),
    .B1(\u3_mem[2] [5]),
    .B2(n_13295),
    .Y(n_24823));
 AOI22xp33_ASAP7_75t_SL g178278 (.A1(n_24806),
    .A2(n_65972),
    .B1(\u3_mem[2] [10]),
    .B2(n_15954),
    .Y(n_24824));
 AOI22xp5_ASAP7_75t_SL g178279 (.A1(n_24806),
    .A2(n_65949),
    .B1(\u3_mem[2] [16]),
    .B2(n_13295),
    .Y(n_24825));
 AOI22xp5_ASAP7_75t_SL g178280 (.A1(n_24806),
    .A2(n_10171),
    .B1(\u3_mem[2] [18]),
    .B2(n_13295),
    .Y(n_24826));
 AOI22xp5_ASAP7_75t_SL g178281 (.A1(n_24806),
    .A2(n_65902),
    .B1(\u3_mem[2] [31]),
    .B2(n_15954),
    .Y(n_24827));
 AOI22xp5_ASAP7_75t_SL g178282 (.A1(n_24806),
    .A2(n_10638),
    .B1(\u3_mem[2] [30]),
    .B2(n_13295),
    .Y(n_24828));
 AOI22xp5_ASAP7_75t_SL g178283 (.A1(n_24806),
    .A2(n_28240),
    .B1(\u3_mem[2] [8]),
    .B2(n_15954),
    .Y(n_24829));
 AOI22xp5_ASAP7_75t_SL g178284 (.A1(n_24806),
    .A2(n_65955),
    .B1(\u3_mem[2] [13]),
    .B2(n_13295),
    .Y(n_24830));
 AOI22xp5_ASAP7_75t_SL g178285 (.A1(n_24806),
    .A2(n_32644),
    .B1(\u3_mem[2] [6]),
    .B2(n_15954),
    .Y(n_24831));
 AOI22xp5_ASAP7_75t_SL g178286 (.A1(n_24806),
    .A2(n_9942),
    .B1(\u3_mem[2] [9]),
    .B2(n_13295),
    .Y(n_24832));
 AOI22xp5_ASAP7_75t_SL g178287 (.A1(n_24806),
    .A2(n_73996),
    .B1(\u3_mem[2] [21]),
    .B2(n_13295),
    .Y(n_24833));
 AOI22xp5_ASAP7_75t_SL g178289 (.A1(n_24806),
    .A2(n_62940),
    .B1(\u3_mem[2] [27]),
    .B2(n_15954),
    .Y(n_24835));
 AOI22xp5_ASAP7_75t_SL g178291 (.A1(n_24806),
    .A2(n_15952),
    .B1(\u3_mem[2] [29]),
    .B2(n_15954),
    .Y(n_24837));
 AOI22xp5_ASAP7_75t_SL g178292 (.A1(n_24806),
    .A2(n_66010),
    .B1(\u3_mem[2] [26]),
    .B2(n_15954),
    .Y(n_24838));
 BUFx2_ASAP7_75t_SL g178335 (.A(n_17584),
    .Y(n_24883));
 INVx1_ASAP7_75t_SL g178338 (.A(in_slt3[10]),
    .Y(n_24886));
 OAI221xp5_ASAP7_75t_SL g178340 (.A1(n_34488),
    .A2(n_24883),
    .B1(n_48057),
    .B2(n_24886),
    .C(n_48640),
    .Y(n_24888));
 AOI22xp5_ASAP7_75t_SL g178423 (.A1(n_35121),
    .A2(\u10_mem[3] [19]),
    .B1(n_61242),
    .B2(n_50551),
    .Y(n_24978));
 NAND2x1_ASAP7_75t_SL g178425 (.A(n_33604),
    .B(u10_wp[1]),
    .Y(n_24975));
 INVx2_ASAP7_75t_SL g178426 (.A(u10_wp[2]),
    .Y(n_534));
 INVx1_ASAP7_75t_SL g178721 (.A(ic1_cfg[6]),
    .Y(n_25293));
 NOR2xp33_ASAP7_75t_SL g178723 (.A(n_25293),
    .B(dma_ack_i[7]),
    .Y(n_25294));
 AOI22xp5_ASAP7_75t_SL g178750 (.A1(n_33024),
    .A2(n_64861),
    .B1(\u6_mem[3] [20]),
    .B2(n_67568),
    .Y(n_25330));
 AOI22xp5_ASAP7_75t_SL g178751 (.A1(n_65932),
    .A2(n_64861),
    .B1(\u6_mem[3] [19]),
    .B2(n_67568),
    .Y(n_25331));
 AOI22xp33_ASAP7_75t_SL g178752 (.A1(n_10194),
    .A2(n_64861),
    .B1(\u6_mem[3] [18]),
    .B2(n_67568),
    .Y(n_25332));
 AOI22xp5_ASAP7_75t_SL g178753 (.A1(n_65952),
    .A2(n_64861),
    .B1(\u6_mem[3] [17]),
    .B2(n_67568),
    .Y(n_25333));
 AOI22xp5_ASAP7_75t_SL g178796 (.A1(n_66011),
    .A2(n_25378),
    .B1(\u7_mem[3] [26]),
    .B2(n_33777),
    .Y(n_25379));
 AND2x4_ASAP7_75t_SL g178797 (.A(n_33774),
    .B(n_30452),
    .Y(n_25378));
 AOI22xp5_ASAP7_75t_SL g178800 (.A1(n_65908),
    .A2(n_25378),
    .B1(n_33777),
    .B2(\u7_mem[3] [27]),
    .Y(n_25380));
 AOI22xp5_ASAP7_75t_SL g178801 (.A1(n_33203),
    .A2(n_25378),
    .B1(n_33777),
    .B2(\u7_mem[3] [0]),
    .Y(n_25381));
 AOI22xp5_ASAP7_75t_SL g178802 (.A1(n_65932),
    .A2(n_25378),
    .B1(\u7_mem[3] [19]),
    .B2(n_33777),
    .Y(n_25382));
 AOI22xp5_ASAP7_75t_SL g178803 (.A1(n_32916),
    .A2(n_25378),
    .B1(\u7_mem[3] [21]),
    .B2(n_33777),
    .Y(n_25383));
 AOI22xp5_ASAP7_75t_SL g178804 (.A1(n_10659),
    .A2(n_25378),
    .B1(n_33777),
    .B2(\u7_mem[3] [30]),
    .Y(n_25384));
 AOI22xp5_ASAP7_75t_SL g178805 (.A1(n_10683),
    .A2(n_25378),
    .B1(n_33777),
    .B2(\u7_mem[3] [29]),
    .Y(n_25385));
 AOI22xp5_ASAP7_75t_SL g178806 (.A1(n_65920),
    .A2(n_25378),
    .B1(n_33777),
    .B2(\u7_mem[3] [28]),
    .Y(n_25386));
 AOI22xp5_ASAP7_75t_SL g178807 (.A1(n_33777),
    .A2(\u7_mem[3] [20]),
    .B1(n_33024),
    .B2(n_25387),
    .Y(n_25388));
 AOI22xp5_ASAP7_75t_SL g178808 (.A1(n_10329),
    .A2(n_25387),
    .B1(\u7_mem[3] [23]),
    .B2(n_33777),
    .Y(n_25389));
 AOI22xp5_ASAP7_75t_SL g178809 (.A1(n_3815),
    .A2(n_25387),
    .B1(n_33777),
    .B2(\u7_mem[3] [1]),
    .Y(n_25390));
 AOI22xp5_ASAP7_75t_SL g178810 (.A1(n_10302),
    .A2(n_25387),
    .B1(\u7_mem[3] [22]),
    .B2(n_33777),
    .Y(n_25391));
 AOI22xp5_ASAP7_75t_SL g178811 (.A1(n_66000),
    .A2(n_25387),
    .B1(\u7_mem[3] [2]),
    .B2(n_33777),
    .Y(n_25392));
 AOI22xp5_ASAP7_75t_SL g178812 (.A1(n_65900),
    .A2(n_25387),
    .B1(n_33777),
    .B2(\u7_mem[3] [31]),
    .Y(n_25393));
 AOI22xp5_ASAP7_75t_SL g178813 (.A1(n_65917),
    .A2(n_25387),
    .B1(\u7_mem[3] [24]),
    .B2(n_33777),
    .Y(n_25394));
 AOI22xp5_ASAP7_75t_SL g178814 (.A1(n_65927),
    .A2(n_25387),
    .B1(\u7_mem[3] [25]),
    .B2(n_33777),
    .Y(n_25395));
 AND2x2_ASAP7_75t_R g178817 (.A(u7_rp[0]),
    .B(n_2691),
    .Y(n_25398));
 OAI22xp5_ASAP7_75t_SL g178833 (.A1(u10_wp[1]),
    .A2(u10_rp[0]),
    .B1(n_25438),
    .B2(n_25439),
    .Y(n_25440));
 INVx4_ASAP7_75t_SL g178834 (.A(u10_rp[0]),
    .Y(n_25439));
 NAND2xp5_ASAP7_75t_SL g178918 (.A(n_25528),
    .B(n_25529),
    .Y(n_25530));
 AOI22xp33_ASAP7_75t_SL g178919 (.A1(u11_din_tmp1[1]),
    .A2(n_13236),
    .B1(in_slt6[3]),
    .B2(n_1523),
    .Y(n_25528));
 NAND2xp33_ASAP7_75t_R g178920 (.A(in_slt6[1]),
    .B(n_46192),
    .Y(n_25529));
 INVxp33_ASAP7_75t_L g179 (.A(n_52770),
    .Y(n_43605));
 NOR2x1_ASAP7_75t_L g179059 (.A(n_1820),
    .B(n_48637),
    .Y(n_25673));
 NOR2x1_ASAP7_75t_L g179061 (.A(n_48053),
    .B(n_48637),
    .Y(n_25674));
 NOR2xp67_ASAP7_75t_SL g179062 (.A(n_34488),
    .B(n_48637),
    .Y(n_25675));
 OAI21xp5_ASAP7_75t_SL g179063 (.A1(n_48637),
    .A2(n_48058),
    .B(n_50459),
    .Y(n_25677));
 OAI21xp5_ASAP7_75t_SL g179065 (.A1(n_21665),
    .A2(n_48637),
    .B(n_50457),
    .Y(n_25678));
 NOR2x1_ASAP7_75t_L g179066 (.A(n_34504),
    .B(n_48637),
    .Y(n_25679));
 NOR2xp67_ASAP7_75t_SL g179067 (.A(n_1678),
    .B(n_48637),
    .Y(n_25680));
 NOR2x1_ASAP7_75t_L g179068 (.A(n_1677),
    .B(n_48637),
    .Y(n_25681));
 NOR2xp67_ASAP7_75t_SL g179069 (.A(n_21673),
    .B(n_48637),
    .Y(n_25682));
 AND2x2_ASAP7_75t_SL g179262 (.A(n_51496),
    .B(n_13988),
    .Y(n_25928));
 BUFx3_ASAP7_75t_SL g179288 (.A(n_25953),
    .Y(n_25954));
 HB1xp67_ASAP7_75t_SL g179289 (.A(n_13968),
    .Y(n_25953));
 BUFx2_ASAP7_75t_SL g179291 (.A(n_25953),
    .Y(n_25956));
 AOI211xp5_ASAP7_75t_SL g179295 (.A1(n_79308),
    .A2(n_25956),
    .B(n_4423),
    .C(n_7735),
    .Y(n_25961));
 AOI21xp5_ASAP7_75t_SL g179298 (.A1(n_37342),
    .A2(n_25954),
    .B(n_14969),
    .Y(n_25964));
 AOI21xp5_ASAP7_75t_SL g179299 (.A1(n_14448),
    .A2(n_25954),
    .B(n_49181),
    .Y(n_25965));
 AOI211xp5_ASAP7_75t_SL g179301 (.A1(n_49180),
    .A2(n_25954),
    .B(n_36364),
    .C(n_49179),
    .Y(n_25967));
 NAND2x1p5_ASAP7_75t_SL g179383 (.A(u4_wp[0]),
    .B(o4_we),
    .Y(n_26050));
 AOI22xp33_ASAP7_75t_SL g179385 (.A1(n_30253),
    .A2(n_65908),
    .B1(n_35910),
    .B2(\u4_mem[3] [27]),
    .Y(n_26054));
 AOI22xp33_ASAP7_75t_SL g179388 (.A1(n_30253),
    .A2(n_65902),
    .B1(n_35910),
    .B2(\u4_mem[3] [31]),
    .Y(n_26055));
 AOI22xp33_ASAP7_75t_SL g179390 (.A1(n_30253),
    .A2(n_65920),
    .B1(\u4_mem[3] [28]),
    .B2(n_35910),
    .Y(n_26057));
 NAND2xp5_ASAP7_75t_SL g179414 (.A(n_56848),
    .B(n_52880),
    .Y(n_26098));
 OAI31xp33_ASAP7_75t_SL g179496 (.A1(oc4_cfg[4]),
    .A2(o8_status[0]),
    .A3(o8_status[1]),
    .B(n_26182),
    .Y(n_26183));
 INVx1_ASAP7_75t_SL g179498 (.A(o8_empty),
    .Y(n_26182));
 AND2x2_ASAP7_75t_SL g179532 (.A(n_33604),
    .B(n_31801),
    .Y(n_26250));
 NAND3x1_ASAP7_75t_SL g179534 (.A(u12_re1),
    .B(n_26254),
    .C(n_35636),
    .Y(n_26255));
 NOR3x1_ASAP7_75t_L g179537 (.A(n_38),
    .B(n_0),
    .C(wb_we_i),
    .Y(n_26254));
 NAND3xp33_ASAP7_75t_SL g179657 (.A(n_195),
    .B(n_36068),
    .C(n_519),
    .Y(n_26376));
 AND3x1_ASAP7_75t_SL g179660 (.A(n_36068),
    .B(n_519),
    .C(n_195),
    .Y(n_26379));
 INVx2_ASAP7_75t_SL g179663 (.A(u5_wp[1]),
    .Y(n_26382));
 AOI22xp33_ASAP7_75t_SL g179664 (.A1(n_26385),
    .A2(n_22715),
    .B1(\u5_mem[0] [29]),
    .B2(n_26386),
    .Y(n_26387));
 BUFx12f_ASAP7_75t_SL g179665 (.A(n_26384),
    .Y(n_26385));
 AND3x4_ASAP7_75t_SL g179666 (.A(n_26383),
    .B(o6_we),
    .C(n_26382),
    .Y(n_26384));
 INVx2_ASAP7_75t_SL g179667 (.A(u5_wp[0]),
    .Y(n_26383));
 INVx3_ASAP7_75t_SL g179668 (.A(n_26384),
    .Y(n_26386));
 AOI22xp5_ASAP7_75t_SL g179669 (.A1(n_26385),
    .A2(n_10640),
    .B1(\u5_mem[0] [30]),
    .B2(n_26386),
    .Y(n_26388));
 AOI22xp5_ASAP7_75t_SL g179670 (.A1(n_26385),
    .A2(n_15920),
    .B1(\u5_mem[0] [31]),
    .B2(n_26389),
    .Y(n_26390));
 INVx3_ASAP7_75t_SL g179671 (.A(n_26384),
    .Y(n_26389));
 AOI22xp5_ASAP7_75t_SL g179672 (.A1(n_26385),
    .A2(n_10198),
    .B1(\u5_mem[0] [19]),
    .B2(n_26386),
    .Y(n_26391));
 AOI22xp5_ASAP7_75t_SL g179673 (.A1(n_26385),
    .A2(n_10171),
    .B1(\u5_mem[0] [18]),
    .B2(n_26389),
    .Y(n_26392));
 AOI22xp5_ASAP7_75t_SL g179674 (.A1(n_26385),
    .A2(n_65952),
    .B1(\u5_mem[0] [17]),
    .B2(n_26386),
    .Y(n_26393));
 AOI22xp5_ASAP7_75t_SL g179675 (.A1(n_26385),
    .A2(n_28276),
    .B1(\u5_mem[0] [16]),
    .B2(n_26386),
    .Y(n_26394));
 AOI22xp5_ASAP7_75t_SL g179676 (.A1(n_26385),
    .A2(n_35041),
    .B1(\u5_mem[0] [13]),
    .B2(n_26386),
    .Y(n_26395));
 AOI22xp5_ASAP7_75t_SL g179677 (.A1(n_26385),
    .A2(n_66869),
    .B1(\u5_mem[0] [5]),
    .B2(n_26386),
    .Y(n_26396));
 AOI22xp5_ASAP7_75t_SL g179679 (.A1(n_26385),
    .A2(n_9942),
    .B1(\u5_mem[0] [9]),
    .B2(n_26386),
    .Y(n_26398));
 AOI22xp5_ASAP7_75t_SL g179680 (.A1(n_26385),
    .A2(n_65972),
    .B1(\u5_mem[0] [10]),
    .B2(n_26386),
    .Y(n_26399));
 AOI22xp5_ASAP7_75t_SL g179681 (.A1(n_65980),
    .A2(n_26385),
    .B1(\u5_mem[0] [8]),
    .B2(n_26386),
    .Y(n_26400));
 AOI22xp33_ASAP7_75t_SL g179682 (.A1(n_26385),
    .A2(n_66856),
    .B1(\u5_mem[0] [3]),
    .B2(n_26386),
    .Y(n_26401));
 AOI22xp5_ASAP7_75t_SL g179683 (.A1(n_26385),
    .A2(n_65969),
    .B1(\u5_mem[0] [7]),
    .B2(n_26389),
    .Y(n_26402));
 AOI22xp5_ASAP7_75t_SL g179684 (.A1(n_26385),
    .A2(n_32644),
    .B1(\u5_mem[0] [6]),
    .B2(n_26389),
    .Y(n_26403));
 AOI22xp5_ASAP7_75t_SL g179685 (.A1(n_26385),
    .A2(n_10000),
    .B1(\u5_mem[0] [11]),
    .B2(n_26386),
    .Y(n_26404));
 AOI22xp5_ASAP7_75t_SL g179686 (.A1(n_26385),
    .A2(n_65941),
    .B1(\u5_mem[0] [22]),
    .B2(n_26389),
    .Y(n_26405));
 AOI22xp5_ASAP7_75t_SL g179687 (.A1(n_26385),
    .A2(n_62940),
    .B1(\u5_mem[0] [27]),
    .B2(n_26386),
    .Y(n_26406));
 AOI22xp5_ASAP7_75t_SL g179688 (.A1(n_26385),
    .A2(n_65930),
    .B1(\u5_mem[0] [23]),
    .B2(n_26389),
    .Y(n_26407));
 AOI22xp5_ASAP7_75t_SL g179689 (.A1(n_26385),
    .A2(n_65925),
    .B1(\u5_mem[0] [25]),
    .B2(n_26389),
    .Y(n_26408));
 AOI22xp5_ASAP7_75t_SL g179690 (.A1(n_26385),
    .A2(n_10026),
    .B1(\u5_mem[0] [12]),
    .B2(n_26386),
    .Y(n_26409));
 AOI22xp33_ASAP7_75t_SL g179691 (.A1(n_26385),
    .A2(n_28330),
    .B1(\u5_mem[0] [2]),
    .B2(n_26386),
    .Y(n_26410));
 AOI22xp5_ASAP7_75t_SL g179692 (.A1(n_26385),
    .A2(n_32916),
    .B1(\u5_mem[0] [21]),
    .B2(n_26389),
    .Y(n_26411));
 AOI22xp5_ASAP7_75t_SL g179693 (.A1(n_26385),
    .A2(n_28424),
    .B1(\u5_mem[0] [24]),
    .B2(n_26389),
    .Y(n_26412));
 AOI22xp5_ASAP7_75t_SL g179694 (.A1(n_26385),
    .A2(n_65920),
    .B1(\u5_mem[0] [28]),
    .B2(n_26389),
    .Y(n_26413));
 AOI22xp5_ASAP7_75t_SL g179695 (.A1(n_26385),
    .A2(n_35437),
    .B1(\u5_mem[0] [26]),
    .B2(n_26389),
    .Y(n_26414));
 AOI22xp5_ASAP7_75t_SL g179696 (.A1(n_26385),
    .A2(n_33024),
    .B1(\u5_mem[0] [20]),
    .B2(n_26389),
    .Y(n_26415));
 AOI22xp5_ASAP7_75t_SL g179697 (.A1(n_26385),
    .A2(n_28913),
    .B1(\u5_mem[0] [15]),
    .B2(n_26389),
    .Y(n_26416));
 AOI22xp5_ASAP7_75t_SL g179698 (.A1(n_26385),
    .A2(n_66032),
    .B1(\u5_mem[0] [14]),
    .B2(n_26389),
    .Y(n_26417));
 AOI22xp33_ASAP7_75t_SL g179699 (.A1(n_26385),
    .A2(n_10891),
    .B1(\u5_mem[0] [1]),
    .B2(n_26386),
    .Y(n_26418));
 AOI22xp33_ASAP7_75t_SL g179700 (.A1(n_26385),
    .A2(n_10924),
    .B1(\u5_mem[0] [0]),
    .B2(n_26389),
    .Y(n_26419));
 AND2x4_ASAP7_75t_SL g179775 (.A(n_26497),
    .B(n_26498),
    .Y(n_26499));
 AND2x2_ASAP7_75t_SL g179776 (.A(u8_wp[0]),
    .B(o9_we),
    .Y(n_26497));
 INVx1_ASAP7_75t_SL g179777 (.A(n_64814),
    .Y(n_26498));
 INVx5_ASAP7_75t_SL g179813 (.A(n_26540),
    .Y(n_26541));
 AND2x2_ASAP7_75t_SL g179814 (.A(rf_we),
    .B(n_26539),
    .Y(n_26540));
 NOR2xp67_ASAP7_75t_L g179815 (.A(n_8177),
    .B(n_21332),
    .Y(n_26539));
 AOI22xp33_ASAP7_75t_SL g179827 (.A1(n_28520),
    .A2(n_26553),
    .B1(\u11_mem[2] [7]),
    .B2(n_61785),
    .Y(n_26556));
 OAI221xp5_ASAP7_75t_SL g179828 (.A1(n_1679),
    .A2(n_34484),
    .B1(n_1705),
    .B2(n_21631),
    .C(n_10941),
    .Y(n_26553));
 INVx1_ASAP7_75t_SL g179851 (.A(ic0_cfg[6]),
    .Y(n_26577));
 OAI22xp5_ASAP7_75t_SL g179852 (.A1(n_11011),
    .A2(n_24672),
    .B1(n_28895),
    .B2(n_26577),
    .Y(n_26579));
 NOR2xp33_ASAP7_75t_SL g179853 (.A(n_26577),
    .B(n_8306),
    .Y(n_26581));
 HB1xp67_ASAP7_75t_SL g179917 (.A(n_32299),
    .Y(n_26645));
 INVxp67_ASAP7_75t_R g179982 (.A(u16_u3_dma_req_r1),
    .Y(n_26711));
 NOR2xp33_ASAP7_75t_R g179983 (.A(dma_ack_i[3]),
    .B(n_25),
    .Y(n_26713));
 NAND2xp5_ASAP7_75t_SL g18 (.A(n_78810),
    .B(n_79326),
    .Y(n_79327));
 INVxp33_ASAP7_75t_R g180 (.A(wb_data_i[28]),
    .Y(n_65918));
 NAND2xp5_ASAP7_75t_SL g180001 (.A(n_23110),
    .B(n_36613),
    .Y(n_26733));
 BUFx3_ASAP7_75t_L g180062 (.A(n_35458),
    .Y(n_26801));
 NOR2xp33_ASAP7_75t_SL g180064 (.A(n_5741),
    .B(n_35458),
    .Y(n_26802));
 OAI22xp33_ASAP7_75t_SL g180065 (.A1(n_35458),
    .A2(n_6972),
    .B1(n_17600),
    .B2(n_28895),
    .Y(n_26803));
 NOR3xp33_ASAP7_75t_SL g180067 (.A(n_26801),
    .B(n_5741),
    .C(n_396),
    .Y(n_26806));
 INVx2_ASAP7_75t_L g180069 (.A(in_slt4[16]),
    .Y(n_26807));
 INVxp67_ASAP7_75t_R g180073 (.A(in_slt4[17]),
    .Y(n_26811));
 INVx1_ASAP7_75t_L g180077 (.A(in_slt4[9]),
    .Y(n_26815));
 INVx1_ASAP7_75t_L g180081 (.A(in_slt4[12]),
    .Y(n_26819));
 INVx1_ASAP7_75t_R g180085 (.A(in_slt4[10]),
    .Y(n_26823));
 INVx2_ASAP7_75t_R g180089 (.A(in_slt4[8]),
    .Y(n_26827));
 INVx1_ASAP7_75t_L g180093 (.A(in_slt4[5]),
    .Y(n_26831));
 INVx1_ASAP7_75t_L g180108 (.A(in_slt4[4]),
    .Y(n_26859));
 OR2x2_ASAP7_75t_SL g180146 (.A(n_1816),
    .B(n_1752),
    .Y(n_26904));
 OAI22xp33_ASAP7_75t_SL g180237 (.A1(u14_u6_en_out_l_44),
    .A2(in_valid_s[0]),
    .B1(n_27003),
    .B2(in_slt0[12]),
    .Y(n_27004));
 INVx1_ASAP7_75t_SL g180238 (.A(ic0_cfg[1]),
    .Y(n_27003));
 AND2x2_ASAP7_75t_SL g180246 (.A(n_31891),
    .B(n_56852),
    .Y(n_27013));
 AOI22xp5_ASAP7_75t_SL g180273 (.A1(n_43318),
    .A2(\u3_mem[0] [9]),
    .B1(\u3_mem[1] [9]),
    .B2(n_43317),
    .Y(n_27038));
 AND3x4_ASAP7_75t_SL g180289 (.A(n_27057),
    .B(n_48105),
    .C(o4_we),
    .Y(n_27058));
 INVx3_ASAP7_75t_SL g180290 (.A(u4_wp[0]),
    .Y(n_27057));
 NAND2x1p5_ASAP7_75t_SL g180291 (.A(n_27059),
    .B(n_27060),
    .Y(n_27061));
 NOR2x1_ASAP7_75t_L g180292 (.A(n_8236),
    .B(u12_we2),
    .Y(n_27059));
 INVx1_ASAP7_75t_SL g180293 (.A(n_1661),
    .Y(n_27060));
 NOR2xp33_ASAP7_75t_SL g180353 (.A(n_6138),
    .B(n_4117),
    .Y(n_27128));
 NAND2xp5_ASAP7_75t_SL g180354 (.A(n_19669),
    .B(n_78952),
    .Y(n_27129));
 AOI221xp5_ASAP7_75t_SL g180356 (.A1(n_27128),
    .A2(n_47631),
    .B1(n_27129),
    .B2(n_34235),
    .C(n_27131),
    .Y(n_27132));
 AND2x2_ASAP7_75t_L g180357 (.A(out_slt7[3]),
    .B(n_46182),
    .Y(n_27131));
 AND2x4_ASAP7_75t_SL g180358 (.A(n_636),
    .B(n_70885),
    .Y(n_27133));
 AND2x4_ASAP7_75t_SL g180359 (.A(n_636),
    .B(n_78274),
    .Y(n_27134));
 NAND4xp25_ASAP7_75t_SL g180360 (.A(n_41435),
    .B(n_2345),
    .C(n_1432),
    .D(n_27135),
    .Y(n_27136));
 AOI22xp33_ASAP7_75t_SL g180361 (.A1(\u8_mem[0] [30]),
    .A2(n_27133),
    .B1(n_27134),
    .B2(\u8_mem[1] [30]),
    .Y(n_27135));
 NAND2xp5_ASAP7_75t_SL g180428 (.A(n_28327),
    .B(n_78810),
    .Y(n_27219));
 A2O1A1Ixp33_ASAP7_75t_SL g180431 (.A1(n_27223),
    .A2(n_27224),
    .B(n_27225),
    .C(n_42258),
    .Y(n_27227));
 NAND2xp5_ASAP7_75t_SL g180432 (.A(n_35407),
    .B(n_50293),
    .Y(n_27223));
 INVx1_ASAP7_75t_L g180433 (.A(n_1842),
    .Y(n_27224));
 INVx4_ASAP7_75t_SL g180434 (.A(n_4788),
    .Y(n_27225));
 NAND3xp33_ASAP7_75t_SL g180441 (.A(n_27234),
    .B(n_27235),
    .C(n_27236),
    .Y(n_27237));
 NAND2xp33_ASAP7_75t_R g180442 (.A(n_40417),
    .B(n_24594),
    .Y(n_27234));
 A2O1A1Ixp33_ASAP7_75t_SL g180443 (.A1(n_40417),
    .A2(n_47551),
    .B(n_1229),
    .C(n_31844),
    .Y(n_27235));
 INVxp67_ASAP7_75t_SL g180444 (.A(n_16895),
    .Y(n_27236));
 AO22x2_ASAP7_75t_SL g180464 (.A1(n_13764),
    .A2(n_543),
    .B1(u11_rp[1]),
    .B2(u11_wp[2]),
    .Y(n_27257));
 AOI22xp5_ASAP7_75t_SL g180508 (.A1(\u4_mem[2] [2]),
    .A2(n_35632),
    .B1(\u4_mem[0] [2]),
    .B2(n_58959),
    .Y(n_27305));
 AOI22xp5_ASAP7_75t_SL g180517 (.A1(n_27315),
    .A2(n_675),
    .B1(n_27316),
    .B2(n_273),
    .Y(n_27317));
 INVx1_ASAP7_75t_SL g180518 (.A(n_273),
    .Y(n_27315));
 INVxp33_ASAP7_75t_R g180519 (.A(n_675),
    .Y(n_27316));
 INVxp67_ASAP7_75t_SL g180521 (.A(n_26428),
    .Y(n_27320));
 AOI22xp33_ASAP7_75t_SL g180534 (.A1(\u3_mem[2] [24]),
    .A2(n_77398),
    .B1(\u3_mem[3] [24]),
    .B2(n_22062),
    .Y(n_27341));
 OAI21xp5_ASAP7_75t_SL g180562 (.A1(n_51041),
    .A2(n_19495),
    .B(n_50293),
    .Y(n_27368));
 NAND4xp25_ASAP7_75t_SL g180564 (.A(n_27368),
    .B(n_27369),
    .C(n_27370),
    .D(n_53369),
    .Y(n_27372));
 NAND2xp5_ASAP7_75t_SL g180565 (.A(n_41491),
    .B(n_50290),
    .Y(n_27369));
 AOI22xp33_ASAP7_75t_L g180566 (.A1(\u7_mem[0] [31]),
    .A2(n_65055),
    .B1(\u7_mem[1] [31]),
    .B2(n_65056),
    .Y(n_27370));
 NAND2xp5_ASAP7_75t_SL g180577 (.A(n_14017),
    .B(n_24350),
    .Y(n_27381));
 AOI22xp33_ASAP7_75t_SL g180578 (.A1(\u4_mem[0] [30]),
    .A2(n_1766),
    .B1(\u4_mem[1] [30]),
    .B2(n_1765),
    .Y(n_27382));
 AOI22xp33_ASAP7_75t_L g180579 (.A1(\u4_mem[2] [30]),
    .A2(n_17624),
    .B1(\u4_mem[3] [30]),
    .B2(n_23531),
    .Y(n_27383));
 NAND4xp25_ASAP7_75t_SL g180714 (.A(n_13824),
    .B(n_35468),
    .C(n_1767),
    .D(n_1807),
    .Y(n_27521));
 AOI22xp5_ASAP7_75t_SL g1809 (.A1(n_58710),
    .A2(n_7285),
    .B1(n_79104),
    .B2(n_43204),
    .Y(n_7288));
 INVxp33_ASAP7_75t_R g181 (.A(wb_data_i[18]),
    .Y(n_65933));
 AOI22xp5_ASAP7_75t_SL g181062 (.A1(\u11_mem[2] [3]),
    .A2(n_61785),
    .B1(n_27878),
    .B2(n_28520),
    .Y(n_27880));
 NAND2xp5_ASAP7_75t_SL g181064 (.A(n_15138),
    .B(n_15139),
    .Y(n_27878));
 NAND3xp33_ASAP7_75t_SL g1811 (.A(n_43205),
    .B(n_7665),
    .C(n_66668),
    .Y(n_7285));
 OAI221xp5_ASAP7_75t_SL g181261 (.A1(n_2523),
    .A2(n_4405),
    .B1(n_46228),
    .B2(n_2524),
    .C(n_28102),
    .Y(n_28103));
 NAND2xp5_ASAP7_75t_SL g181262 (.A(n_47551),
    .B(n_4515),
    .Y(n_28102));
 AOI21xp5_ASAP7_75t_SL g181270 (.A1(n_13899),
    .A2(n_13898),
    .B(n_28110),
    .Y(n_28111));
 XNOR2xp5_ASAP7_75t_SL g181280 (.A(n_65325),
    .B(n_28121),
    .Y(n_28122));
 NAND2xp5_ASAP7_75t_SL g181281 (.A(n_30078),
    .B(n_71392),
    .Y(n_28121));
 AOI22xp5_ASAP7_75t_SL g181393 (.A1(n_46477),
    .A2(\u10_mem[0] [12]),
    .B1(n_46478),
    .B2(n_28747),
    .Y(n_28235));
 NAND2xp5_ASAP7_75t_SL g181397 (.A(n_51051),
    .B(n_31311),
    .Y(n_28239));
 INVx3_ASAP7_75t_SL g181400 (.A(n_9880),
    .Y(n_28240));
 NAND2xp5_ASAP7_75t_SL g181402 (.A(n_78810),
    .B(n_28370),
    .Y(n_28246));
 INVx2_ASAP7_75t_SL g181410 (.A(n_9735),
    .Y(n_28251));
 INVx2_ASAP7_75t_SL g181433 (.A(n_10112),
    .Y(n_28276));
 AOI22xp5_ASAP7_75t_SL g181449 (.A1(n_53101),
    .A2(\u5_mem[0] [2]),
    .B1(\u5_mem[2] [2]),
    .B2(n_65643),
    .Y(n_28294));
 INVx2_ASAP7_75t_SL g181469 (.A(n_10434),
    .Y(n_28316));
 NAND2xp5_ASAP7_75t_SL g181479 (.A(n_78943),
    .B(n_47306),
    .Y(n_28327));
 INVx3_ASAP7_75t_SL g181484 (.A(n_9822),
    .Y(n_28330));
 AOI22xp5_ASAP7_75t_SL g181507 (.A1(n_77853),
    .A2(\u6_mem[2] [15]),
    .B1(\u6_mem[3] [15]),
    .B2(n_41152),
    .Y(n_28364));
 AOI22xp5_ASAP7_75t_SL g181508 (.A1(crac_out[7]),
    .A2(n_28367),
    .B1(n_17578),
    .B2(n_17579),
    .Y(n_28368));
 INVx6_ASAP7_75t_SL g181509 (.A(n_22852),
    .Y(n_28367));
 NAND2xp5_ASAP7_75t_SL g181510 (.A(n_78041),
    .B(n_28370),
    .Y(n_28371));
 NAND2x1_ASAP7_75t_SL g181512 (.A(n_78950),
    .B(n_28364),
    .Y(n_28370));
 INVx2_ASAP7_75t_SL g181523 (.A(n_10303),
    .Y(n_28381));
 AOI22xp33_ASAP7_75t_SL g181532 (.A1(n_58959),
    .A2(\u4_mem[0] [12]),
    .B1(\u4_mem[2] [12]),
    .B2(n_35632),
    .Y(n_28391));
 AND2x2_ASAP7_75t_R g181550 (.A(n_31579),
    .B(n_4042),
    .Y(n_28413));
 INVx2_ASAP7_75t_SL g181557 (.A(n_10408),
    .Y(n_28424));
 AND2x4_ASAP7_75t_SL g181571_dup194251 (.A(n_503),
    .B(n_33100),
    .Y(n_43537));
 NAND2xp67_ASAP7_75t_SL g181574 (.A(n_782),
    .B(n_28391),
    .Y(n_28441));
 NAND4xp25_ASAP7_75t_SL g181575 (.A(n_21996),
    .B(n_35467),
    .C(n_1754),
    .D(n_1809),
    .Y(n_28443));
 AOI22xp5_ASAP7_75t_SL g181634 (.A1(n_31779),
    .A2(n_28520),
    .B1(\u11_mem[2] [14]),
    .B2(n_61785),
    .Y(n_28521));
 INVx5_ASAP7_75t_SL g181635 (.A(n_23289),
    .Y(n_28520));
 OAI21xp33_ASAP7_75t_SL g181642 (.A1(n_78410),
    .A2(n_28528),
    .B(n_179),
    .Y(n_28529));
 NOR2xp33_ASAP7_75t_R g181643 (.A(n_14385),
    .B(n_24741),
    .Y(n_28528));
 AOI21xp5_ASAP7_75t_SL g181705 (.A1(n_41612),
    .A2(u16_u4_dma_req_r1),
    .B(n_28594),
    .Y(n_28595));
 NOR2xp33_ASAP7_75t_R g181707 (.A(dma_ack_i[4]),
    .B(n_83),
    .Y(n_28594));
 AOI21xp5_ASAP7_75t_SL g181757 (.A1(n_31273),
    .A2(u16_u6_dma_req_r1),
    .B(n_28662),
    .Y(n_28663));
 NOR2xp33_ASAP7_75t_R g181759 (.A(dma_ack_i[6]),
    .B(n_86),
    .Y(n_28662));
 NOR3xp33_ASAP7_75t_SL g181760 (.A(n_8186),
    .B(n_26577),
    .C(dma_ack_i[6]),
    .Y(n_28664));
 INVx1_ASAP7_75t_SL g181765 (.A(n_29618),
    .Y(n_28669));
 INVx3_ASAP7_75t_L g181766 (.A(n_10867),
    .Y(n_10889));
 AOI221xp5_ASAP7_75t_SL g181767 (.A1(u13_intm_r[5]),
    .A2(n_7082),
    .B1(n_8174),
    .B2(i4_dout[5]),
    .C(n_28673),
    .Y(n_28674));
 OAI22xp5_ASAP7_75t_SL g181768 (.A1(n_28671),
    .A2(n_28669),
    .B1(n_10889),
    .B2(n_28672),
    .Y(n_28673));
 INVxp67_ASAP7_75t_SL g181769 (.A(oc0_cfg[5]),
    .Y(n_28671));
 INVx1_ASAP7_75t_L g181770 (.A(crac_din[5]),
    .Y(n_28672));
 NOR3xp33_ASAP7_75t_SL g181785 (.A(n_5748),
    .B(n_2596),
    .C(n_28689),
    .Y(n_28690));
 BUFx3_ASAP7_75t_SL g181786 (.A(oc2_cfg[2]),
    .Y(n_28689));
 INVx1_ASAP7_75t_R g181787 (.A(n_28689),
    .Y(n_28691));
 AOI22xp5_ASAP7_75t_SL g181788 (.A1(n_6961),
    .A2(n_28689),
    .B1(n_7083),
    .B2(n_223),
    .Y(n_28692));
 NOR2xp33_ASAP7_75t_SL g181792 (.A(n_79019),
    .B(n_28689),
    .Y(n_28696));
 NAND2xp5_ASAP7_75t_SL g181838 (.A(n_28746),
    .B(n_1209),
    .Y(n_28747));
 AOI22xp5_ASAP7_75t_SL g181839 (.A1(n_1666),
    .A2(in_slt4[14]),
    .B1(in_slt4[12]),
    .B2(n_28745),
    .Y(n_28746));
 INVxp67_ASAP7_75t_SL g181843 (.A(n_17606),
    .Y(n_28745));
 INVx1_ASAP7_75t_R g181864 (.A(u10_rp[2]),
    .Y(n_28774));
 OAI22xp5_ASAP7_75t_SL g181894 (.A1(n_1919),
    .A2(n_28808),
    .B1(n_31535),
    .B2(n_28810),
    .Y(n_28811));
 NOR2x1_ASAP7_75t_SL g181895 (.A(n_1920),
    .B(n_31535),
    .Y(n_28808));
 NAND2xp33_ASAP7_75t_R g181896 (.A(n_1919),
    .B(u2_res_cnt[0]),
    .Y(n_28810));
 NOR3xp33_ASAP7_75t_L g181899 (.A(n_21335),
    .B(n_28926),
    .C(n_15269),
    .Y(n_28814));
 AND2x2_ASAP7_75t_L g181936 (.A(in_valid_s[2]),
    .B(u14_u8_en_out_l_44),
    .Y(n_28848));
 AOI21xp5_ASAP7_75t_SL g181937 (.A1(n_13598),
    .A2(n_13599),
    .B(n_28848),
    .Y(n_28849));
 NAND3xp33_ASAP7_75t_SL g181939 (.A(n_28848),
    .B(n_295),
    .C(n_20426),
    .Y(n_28852));
 NOR3xp33_ASAP7_75t_SL g181964 (.A(n_29934),
    .B(n_34526),
    .C(n_28879),
    .Y(n_28880));
 INVxp67_ASAP7_75t_SL g181966 (.A(n_25294),
    .Y(n_28879));
 OAI21xp5_ASAP7_75t_SL g181968 (.A1(n_19007),
    .A2(n_19006),
    .B(n_64297),
    .Y(n_28881));
 INVx1_ASAP7_75t_SL g181970 (.A(u15_valid_r),
    .Y(n_28884));
 AND2x2_ASAP7_75t_R g181972 (.A(u15_rdd3),
    .B(n_28884),
    .Y(n_28885));
 AO21x1_ASAP7_75t_SL g181979 (.A1(n_1863),
    .A2(n_7414),
    .B(n_176),
    .Y(n_28893));
 AOI22xp5_ASAP7_75t_SL g181981 (.A1(n_10565),
    .A2(n_17687),
    .B1(n_11006),
    .B2(n_47740),
    .Y(n_28901));
 OR2x6_ASAP7_75t_SL g181983 (.A(n_10563),
    .B(wb_addr_i[4]),
    .Y(n_28895));
 INVx1_ASAP7_75t_SL g181986 (.A(n_11011),
    .Y(n_11006));
 BUFx6f_ASAP7_75t_SL g181987 (.A(n_11000),
    .Y(n_11011));
 INVxp33_ASAP7_75t_R g182 (.A(wb_data_i[7]),
    .Y(n_65967));
 NAND2x2_ASAP7_75t_SL g182013 (.A(n_29005),
    .B(u11_wp[1]),
    .Y(n_28952));
 HB1xp67_ASAP7_75t_SL g182015 (.A(u11_wp[1]),
    .Y(n_28948));
 NAND2xp5_ASAP7_75t_SL g182016 (.A(n_23286),
    .B(n_28948),
    .Y(n_28950));
 AND3x4_ASAP7_75t_SL g182018 (.A(n_29005),
    .B(u11_wp[1]),
    .C(n_217),
    .Y(n_28953));
 INVx4_ASAP7_75t_SL g182019 (.A(u11_wp[1]),
    .Y(n_28954));
 OAI22xp5_ASAP7_75t_SL g182020 (.A1(u11_rp[0]),
    .A2(u11_wp[1]),
    .B1(n_28954),
    .B2(n_13027),
    .Y(n_28955));
 HB1xp67_ASAP7_75t_L g182064 (.A(n_11312),
    .Y(n_29003));
 AND2x4_ASAP7_75t_L g182065 (.A(n_29004),
    .B(n_29005),
    .Y(n_29006));
 AND2x2_ASAP7_75t_SL g182066 (.A(u11_wp[1]),
    .B(n_11312),
    .Y(n_29004));
 AND2x4_ASAP7_75t_SL g182067 (.A(n_21226),
    .B(n_7694),
    .Y(n_29005));
 INVx2_ASAP7_75t_SL g182069 (.A(n_29007),
    .Y(n_29008));
 NAND2x1_ASAP7_75t_SL g182070 (.A(n_12908),
    .B(n_29005),
    .Y(n_29007));
 INVx3_ASAP7_75t_SL g182073 (.A(n_29007),
    .Y(n_29011));
 AOI22xp33_ASAP7_75t_SL g182085 (.A1(n_29008),
    .A2(n_26553),
    .B1(\u11_mem[0] [7]),
    .B2(n_4784),
    .Y(n_29024));
 AOI22xp5_ASAP7_75t_SL g182102 (.A1(n_29011),
    .A2(n_4956),
    .B1(\u11_mem[0] [11]),
    .B2(n_4784),
    .Y(n_29041));
 INVx2_ASAP7_75t_SL g182133 (.A(n_29073),
    .Y(n_29074));
 AND4x2_ASAP7_75t_SL g182134 (.A(n_295),
    .B(n_172),
    .C(in_valid_s[2]),
    .D(u14_u8_en_out_l_44),
    .Y(n_29073));
 NOR2xp33_ASAP7_75t_SL g182135 (.A(n_36289),
    .B(n_1701),
    .Y(n_29076));
 NOR2xp33_ASAP7_75t_SL g182138 (.A(n_29074),
    .B(n_14313),
    .Y(n_29078));
 NOR2xp33_ASAP7_75t_SL g182140 (.A(n_36289),
    .B(n_14309),
    .Y(n_29080));
 NOR2xp33_ASAP7_75t_SL g182142 (.A(n_36289),
    .B(n_1704),
    .Y(n_29082));
 NOR2xp33_ASAP7_75t_SL g182148 (.A(n_36289),
    .B(n_1707),
    .Y(n_29088));
 NOR2xp33_ASAP7_75t_SL g182152 (.A(n_36289),
    .B(n_1680),
    .Y(n_29092));
 NOR2xp33_ASAP7_75t_SL g182154 (.A(n_36289),
    .B(n_1681),
    .Y(n_29094));
 NOR2xp33_ASAP7_75t_SL g182156 (.A(n_36289),
    .B(n_21631),
    .Y(n_29096));
 NOR2xp33_ASAP7_75t_SL g182158 (.A(n_36289),
    .B(n_21638),
    .Y(n_29098));
 NOR2xp33_ASAP7_75t_SL g182160 (.A(n_36289),
    .B(n_21646),
    .Y(n_29100));
 NOR2xp33_ASAP7_75t_SL g182162 (.A(n_36289),
    .B(n_21697),
    .Y(n_29102));
 NOR2xp33_ASAP7_75t_SL g182164 (.A(n_36289),
    .B(n_21705),
    .Y(n_29104));
 NOR2xp33_ASAP7_75t_SL g182166 (.A(n_36289),
    .B(n_21709),
    .Y(n_29106));
 INVx1_ASAP7_75t_R g182367 (.A(n_425),
    .Y(n_29310));
 NAND2xp5_ASAP7_75t_SL g182370 (.A(n_31844),
    .B(n_29310),
    .Y(n_29312));
 INVxp67_ASAP7_75t_SL g182371 (.A(n_29312),
    .Y(n_29314));
 AOI22xp33_ASAP7_75t_SL g182412 (.A1(n_32916),
    .A2(n_64861),
    .B1(n_67568),
    .B2(\u6_mem[3] [21]),
    .Y(n_29355));
 AOI22xp5_ASAP7_75t_SL g182413 (.A1(n_10302),
    .A2(n_64861),
    .B1(\u6_mem[3] [22]),
    .B2(n_67568),
    .Y(n_29356));
 AOI22xp5_ASAP7_75t_SL g182414 (.A1(n_10329),
    .A2(n_64861),
    .B1(\u6_mem[3] [23]),
    .B2(n_35215),
    .Y(n_29358));
 INVx1_ASAP7_75t_SL g182417 (.A(n_2663),
    .Y(n_29361));
 INVxp67_ASAP7_75t_SL g182419 (.A(u7_wp[0]),
    .Y(n_29362));
 XOR2xp5_ASAP7_75t_SL g182420 (.A(n_2663),
    .B(n_64714),
    .Y(n_29364));
 NOR5xp2_ASAP7_75t_SL g182421 (.A(n_2753),
    .B(n_503),
    .C(n_29362),
    .D(n_2752),
    .E(u7_wp[2]),
    .Y(n_29365));
 NOR2xp33_ASAP7_75t_SL g182422 (.A(n_29362),
    .B(n_64714),
    .Y(n_29366));
 INVx1_ASAP7_75t_SL g182485 (.A(n_56847),
    .Y(n_29495));
 NOR2xp33_ASAP7_75t_SL g182517 (.A(n_34505),
    .B(n_48056),
    .Y(n_29527));
 NOR2xp33_ASAP7_75t_SL g182520 (.A(n_34505),
    .B(n_14301),
    .Y(n_29529));
 NOR2xp33_ASAP7_75t_SL g182522 (.A(n_34505),
    .B(n_1677),
    .Y(n_29531));
 NOR2xp33_ASAP7_75t_SL g182524 (.A(n_34505),
    .B(n_1678),
    .Y(n_29533));
 NOR2xp33_ASAP7_75t_SL g182534 (.A(n_34505),
    .B(n_48053),
    .Y(n_29543));
 NOR2xp33_ASAP7_75t_SL g182536 (.A(n_34505),
    .B(n_1820),
    .Y(n_29545));
 NOR2xp33_ASAP7_75t_SL g182538 (.A(n_34505),
    .B(n_24886),
    .Y(n_29547));
 NOR2xp33_ASAP7_75t_SL g182540 (.A(n_34505),
    .B(n_1714),
    .Y(n_29549));
 NOR2xp33_ASAP7_75t_SL g182544 (.A(n_34505),
    .B(n_48058),
    .Y(n_29553));
 NOR2xp33_ASAP7_75t_SL g182546 (.A(n_34505),
    .B(n_21665),
    .Y(n_29555));
 NOR2xp33_ASAP7_75t_SL g182548 (.A(n_34505),
    .B(n_21673),
    .Y(n_29557));
 NOR3x1_ASAP7_75t_L g182605 (.A(n_8311),
    .B(wb_addr_i[3]),
    .C(wb_addr_i[4]),
    .Y(n_29618));
 NAND2x1_ASAP7_75t_SL g182607 (.A(rf_we),
    .B(n_29618),
    .Y(n_29619));
 O2A1O1Ixp5_ASAP7_75t_SL g182616 (.A1(n_17626),
    .A2(n_7641),
    .B(n_34475),
    .C(n_38369),
    .Y(n_29630));
 INVx1_ASAP7_75t_SL g182630 (.A(n_195),
    .Y(n_29657));
 AND2x2_ASAP7_75t_SL g182631 (.A(u4_wp[2]),
    .B(n_29658),
    .Y(n_29659));
 INVx1_ASAP7_75t_SL g182632 (.A(n_29657),
    .Y(n_29658));
 AOI22xp5_ASAP7_75t_SL g182633 (.A1(n_28240),
    .A2(n_67247),
    .B1(n_29658),
    .B2(n_67248),
    .Y(n_29661));
 OAI21xp5_ASAP7_75t_SL g182635 (.A1(n_48107),
    .A2(n_17569),
    .B(n_29658),
    .Y(n_29662));
 NAND2xp5_ASAP7_75t_SL g182657 (.A(n_29687),
    .B(n_775),
    .Y(n_29688));
 AOI22xp5_ASAP7_75t_SL g182658 (.A1(n_58959),
    .A2(\u4_mem[0] [3]),
    .B1(\u4_mem[2] [3]),
    .B2(n_35632),
    .Y(n_29687));
 INVx2_ASAP7_75t_SL g182756 (.A(u4_wp[0]),
    .Y(n_29787));
 BUFx12f_ASAP7_75t_SL g182759 (.A(n_33654),
    .Y(n_29790));
 AOI21xp33_ASAP7_75t_SL g182844 (.A1(n_34420),
    .A2(u10_din_tmp1[10]),
    .B(n_29884),
    .Y(n_29885));
 AND4x2_ASAP7_75t_SL g182846 (.A(n_220),
    .B(u14_u7_en_out_l_44),
    .C(in_valid_s[1]),
    .D(n_73),
    .Y(n_29881));
 NOR2xp33_ASAP7_75t_SL g182847 (.A(n_29883),
    .B(n_21669),
    .Y(n_29884));
 INVx4_ASAP7_75t_SL g182848 (.A(n_29881),
    .Y(n_29883));
 AOI21xp33_ASAP7_75t_SL g182851 (.A1(n_34420),
    .A2(u10_din_tmp1[1]),
    .B(n_29888),
    .Y(n_29889));
 NOR2xp33_ASAP7_75t_SL g182852 (.A(n_29883),
    .B(n_26831),
    .Y(n_29888));
 AOI21xp33_ASAP7_75t_SL g182853 (.A1(n_34420),
    .A2(u10_din_tmp1[4]),
    .B(n_29890),
    .Y(n_29891));
 NOR2xp33_ASAP7_75t_SL g182854 (.A(n_29883),
    .B(n_26827),
    .Y(n_29890));
 AOI21xp33_ASAP7_75t_SL g182859 (.A1(n_34420),
    .A2(u10_din_tmp1[5]),
    .B(n_29896),
    .Y(n_29897));
 NOR2xp33_ASAP7_75t_SL g182860 (.A(n_29883),
    .B(n_26815),
    .Y(n_29896));
 AOI21xp33_ASAP7_75t_SL g182861 (.A1(n_34420),
    .A2(u10_din_tmp1[13]),
    .B(n_29898),
    .Y(n_29899));
 NOR2xp33_ASAP7_75t_SL g182862 (.A(n_29883),
    .B(n_26811),
    .Y(n_29898));
 AOI21xp33_ASAP7_75t_SL g182865 (.A1(n_34420),
    .A2(u10_din_tmp1[9]),
    .B(n_29902),
    .Y(n_29903));
 NOR2xp33_ASAP7_75t_SL g182866 (.A(n_29883),
    .B(n_21878),
    .Y(n_29902));
 AOI21xp33_ASAP7_75t_SL g182867 (.A1(n_34420),
    .A2(u10_din_tmp1[2]),
    .B(n_29904),
    .Y(n_29905));
 NOR2xp33_ASAP7_75t_SL g182868 (.A(n_29883),
    .B(n_14292),
    .Y(n_29904));
 AOI21xp33_ASAP7_75t_SL g182869 (.A1(n_34420),
    .A2(u10_din_tmp1[15]),
    .B(n_29906),
    .Y(n_29907));
 NOR2xp33_ASAP7_75t_SL g182870 (.A(n_29883),
    .B(n_1699),
    .Y(n_29906));
 AOI21xp33_ASAP7_75t_SL g182871 (.A1(n_34420),
    .A2(u10_din_tmp1[14]),
    .B(n_29908),
    .Y(n_29909));
 NOR2xp33_ASAP7_75t_SL g182872 (.A(n_29883),
    .B(n_11693),
    .Y(n_29908));
 AOI21xp33_ASAP7_75t_SL g182873 (.A1(n_34420),
    .A2(u10_din_tmp1[7]),
    .B(n_29910),
    .Y(n_29911));
 NOR2xp33_ASAP7_75t_SL g182874 (.A(n_29883),
    .B(n_14280),
    .Y(n_29910));
 AOI21xp33_ASAP7_75t_SL g182877 (.A1(n_34420),
    .A2(u10_din_tmp1[3]),
    .B(n_29914),
    .Y(n_29915));
 NOR2xp33_ASAP7_75t_SL g182878 (.A(n_29883),
    .B(n_64696),
    .Y(n_29914));
 INVx2_ASAP7_75t_SL g182896 (.A(ic1_cfg[0]),
    .Y(n_29934));
 OAI211xp5_ASAP7_75t_L g182899 (.A1(n_34524),
    .A2(n_34525),
    .B(n_17687),
    .C(n_25294),
    .Y(n_29938));
 OAI21xp33_ASAP7_75t_SL g182901 (.A1(n_34524),
    .A2(n_34525),
    .B(n_17687),
    .Y(n_29939));
 O2A1O1Ixp5_ASAP7_75t_SL g182902 (.A1(n_14820),
    .A2(n_14821),
    .B(n_17687),
    .C(n_17690),
    .Y(n_29940));
 AOI221xp5_ASAP7_75t_SL g182911 (.A1(n_36361),
    .A2(out_slt7[7]),
    .B1(n_37341),
    .B2(n_25954),
    .C(n_4415),
    .Y(n_29949));
 INVxp67_ASAP7_75t_L g182917 (.A(u5_rp[0]),
    .Y(n_13405));
 INVxp33_ASAP7_75t_R g183 (.A(wb_data_i[2]),
    .Y(n_65998));
 AOI21xp33_ASAP7_75t_SL g183006 (.A1(n_30059),
    .A2(n_30060),
    .B(n_30061),
    .Y(n_30062));
 INVx1_ASAP7_75t_SL g183007 (.A(n_2980),
    .Y(n_30059));
 INVx1_ASAP7_75t_SL g183008 (.A(n_2522),
    .Y(n_30060));
 NAND2xp5_ASAP7_75t_SL g183009 (.A(n_43083),
    .B(n_15020),
    .Y(n_30061));
 AND2x6_ASAP7_75t_SL g183025 (.A(u4_rp[1]),
    .B(u4_rp[2]),
    .Y(n_30078));
 OAI22xp5_ASAP7_75t_SL g183172 (.A1(n_10659),
    .A2(n_35911),
    .B1(n_47390),
    .B2(\u4_mem[3] [30]),
    .Y(n_30235));
 AOI22xp5_ASAP7_75t_SL g183188 (.A1(n_65975),
    .A2(n_30253),
    .B1(\u4_mem[3] [10]),
    .B2(n_35911),
    .Y(n_30254));
 OAI211xp5_ASAP7_75t_SL g183255 (.A1(n_37051),
    .A2(n_35463),
    .B(n_30330),
    .C(n_30331),
    .Y(n_30332));
 AOI22xp33_ASAP7_75t_L g183256 (.A1(\u4_mem[2] [25]),
    .A2(n_17624),
    .B1(\u4_mem[3] [25]),
    .B2(n_23531),
    .Y(n_30330));
 AOI21xp33_ASAP7_75t_SL g183257 (.A1(n_26733),
    .A2(n_24350),
    .B(n_24351),
    .Y(n_30331));
 AND2x2_ASAP7_75t_SL g183349 (.A(u14_u6_en_out_l_44),
    .B(in_valid_s[0]),
    .Y(n_17399));
 AND2x2_ASAP7_75t_SL g183362 (.A(u7_wp[0]),
    .B(o8_we),
    .Y(n_30452));
 NAND2x1_ASAP7_75t_SL g183363 (.A(o8_we),
    .B(u7_wp[0]),
    .Y(n_30453));
 AOI22xp33_ASAP7_75t_L g183375 (.A1(\u6_mem[1] [29]),
    .A2(n_48415),
    .B1(\u6_mem[3] [29]),
    .B2(n_17704),
    .Y(n_30469));
 NAND2xp5_ASAP7_75t_SL g183377 (.A(n_31107),
    .B(n_78810),
    .Y(n_30471));
 AOI22xp33_ASAP7_75t_SL g183378 (.A1(\u6_mem[0] [29]),
    .A2(n_79305),
    .B1(\u6_mem[2] [29]),
    .B2(n_79306),
    .Y(n_30472));
 AOI22xp5_ASAP7_75t_SL g183511 (.A1(n_71972),
    .A2(\u3_mem[3] [2]),
    .B1(n_50388),
    .B2(\u3_mem[2] [2]),
    .Y(n_30616));
 NAND2xp5_ASAP7_75t_SL g183901 (.A(n_31056),
    .B(n_31057),
    .Y(n_31058));
 AOI22xp33_ASAP7_75t_SL g183902 (.A1(\u3_mem[1] [3]),
    .A2(n_43317),
    .B1(\u3_mem[0] [3]),
    .B2(n_43318),
    .Y(n_31056));
 AOI22xp5_ASAP7_75t_SL g183903 (.A1(\u3_mem[3] [3]),
    .A2(n_71972),
    .B1(\u3_mem[2] [3]),
    .B2(n_50388),
    .Y(n_31057));
 OAI211xp5_ASAP7_75t_L g183923 (.A1(n_4318),
    .A2(n_7665),
    .B(n_43201),
    .C(n_66682),
    .Y(n_31078));
 NAND2xp5_ASAP7_75t_SL g183946 (.A(n_78956),
    .B(n_63778),
    .Y(n_31107));
 AOI21xp5_ASAP7_75t_SL g183967 (.A1(n_31127),
    .A2(u16_u2_dma_req_r1),
    .B(n_31128),
    .Y(n_31129));
 INVx1_ASAP7_75t_SL g183968 (.A(n_28881),
    .Y(n_31127));
 NOR2xp33_ASAP7_75t_R g183969 (.A(dma_ack_i[2]),
    .B(n_33),
    .Y(n_31128));
 INVxp33_ASAP7_75t_R g184 (.A(wb_data_i[24]),
    .Y(n_65911));
 AOI21xp5_ASAP7_75t_SL g184025 (.A1(n_79205),
    .A2(n_79177),
    .B(n_31190),
    .Y(n_31191));
 OAI22xp33_ASAP7_75t_SL g184027 (.A1(n_13266),
    .A2(n_21876),
    .B1(n_2689),
    .B2(n_3996),
    .Y(n_31190));
 INVx1_ASAP7_75t_SL g184056 (.A(u9_wp[0]),
    .Y(n_113));
 INVx1_ASAP7_75t_SL g184057 (.A(u14_u6_en_out_l2),
    .Y(n_31227));
 AND4x2_ASAP7_75t_SL g184059 (.A(n_31227),
    .B(n_113),
    .C(u14_u6_en_out_l_44),
    .D(in_valid_s[0]),
    .Y(n_31228));
 OAI21xp5_ASAP7_75t_SL g184089 (.A1(n_2546),
    .A2(n_2373),
    .B(n_28664),
    .Y(n_31272));
 AOI22xp5_ASAP7_75t_SL g184114 (.A1(\u7_mem[1] [0]),
    .A2(n_49617),
    .B1(\u7_mem[3] [0]),
    .B2(n_49618),
    .Y(n_31311));
 NAND3xp33_ASAP7_75t_SL g184164 (.A(n_59763),
    .B(n_31396),
    .C(u2_res_cnt[2]),
    .Y(n_31397));
 NAND2xp5_ASAP7_75t_SL g184212 (.A(n_31890),
    .B(n_56855),
    .Y(n_31445));
 NAND2xp5_ASAP7_75t_SL g184219 (.A(n_16858),
    .B(n_79176),
    .Y(n_31455));
 NAND2xp5_ASAP7_75t_L g184294 (.A(u2_res_cnt[1]),
    .B(u2_res_cnt[0]),
    .Y(n_31534));
 OR2x6_ASAP7_75t_SL g184295 (.A(n_50091),
    .B(n_20783),
    .Y(n_31535));
 XOR2xp5_ASAP7_75t_SL g184298 (.A(n_27317),
    .B(n_26428),
    .Y(n_31538));
 INVx1_ASAP7_75t_SL g184324 (.A(u14_u3_en_out_l2),
    .Y(n_31579));
 AND2x4_ASAP7_75t_L g184483 (.A(n_523),
    .B(n_21261),
    .Y(n_31720));
 NOR2xp33_ASAP7_75t_L g184487 (.A(u2_sync_beat),
    .B(u2_sync_resume),
    .Y(n_31724));
 AND3x1_ASAP7_75t_R g184489 (.A(n_47740),
    .B(n_387),
    .C(n_35655),
    .Y(n_31726));
 OA22x2_ASAP7_75t_SL g184495 (.A1(n_17584),
    .A2(n_28895),
    .B1(n_176),
    .B2(n_6960),
    .Y(n_31732));
 AND2x2_ASAP7_75t_SL g184496 (.A(n_56848),
    .B(n_52880),
    .Y(n_31733));
 OR2x2_ASAP7_75t_SL g184503 (.A(n_4280),
    .B(n_18857),
    .Y(n_31740));
 OR2x6_ASAP7_75t_SL g184504 (.A(n_47787),
    .B(n_18964),
    .Y(n_31741));
 AOI22xp33_ASAP7_75t_R g184505 (.A1(\u7_mem[0] [24]),
    .A2(n_65055),
    .B1(\u7_mem[1] [24]),
    .B2(n_65056),
    .Y(n_31742));
 AOI22xp33_ASAP7_75t_R g184506 (.A1(\u7_mem[0] [26]),
    .A2(n_65055),
    .B1(n_65056),
    .B2(\u7_mem[1] [26]),
    .Y(n_31743));
 AO22x1_ASAP7_75t_SL g184510 (.A1(\u10_mem[0] [23]),
    .A2(n_11548),
    .B1(\u10_mem[1] [23]),
    .B2(n_14825),
    .Y(n_31747));
 OR2x2_ASAP7_75t_L g184511 (.A(n_35632),
    .B(n_50709),
    .Y(n_31748));
 XNOR2xp5_ASAP7_75t_SL g184513 (.A(n_321),
    .B(n_146),
    .Y(n_31750));
 XNOR2xp5_ASAP7_75t_SL g184517 (.A(u5_wp[2]),
    .B(n_37311),
    .Y(n_31754));
 NOR4xp25_ASAP7_75t_SL g184533 (.A(n_29657),
    .B(n_24632),
    .C(u4_wp[2]),
    .D(n_14546),
    .Y(n_31770));
 AO21x1_ASAP7_75t_SL g184540 (.A1(u11_din_tmp1[9]),
    .A2(n_13236),
    .B(n_16436),
    .Y(n_31777));
 AO21x1_ASAP7_75t_SL g184542 (.A1(u11_din_tmp1[14]),
    .A2(n_13236),
    .B(n_18089),
    .Y(n_31779));
 AO21x1_ASAP7_75t_SL g184544 (.A1(u11_din_tmp1[12]),
    .A2(n_13236),
    .B(n_18480),
    .Y(n_31781));
 AO221x1_ASAP7_75t_SL g184549 (.A1(n_24336),
    .A2(u10_din_tmp1[8]),
    .B1(n_1666),
    .B2(in_slt4[10]),
    .C(n_17608),
    .Y(n_31786));
 AO22x1_ASAP7_75t_SL g184558 (.A1(n_14821),
    .A2(\u10_mem[2] [23]),
    .B1(n_21092),
    .B2(\u10_mem[3] [23]),
    .Y(n_31795));
 AND2x2_ASAP7_75t_SL g184562 (.A(n_25438),
    .B(n_234),
    .Y(n_31801));
 NOR4xp25_ASAP7_75t_SL g184582 (.A(n_2235),
    .B(n_7231),
    .C(n_8299),
    .D(n_8256),
    .Y(n_31821));
 XOR2xp5_ASAP7_75t_L g184595 (.A(n_2462),
    .B(n_23508),
    .Y(n_31834));
 NOR3xp33_ASAP7_75t_SL g184605 (.A(n_19133),
    .B(n_34539),
    .C(n_43082),
    .Y(n_31844));
 NAND2x1_ASAP7_75t_SL g184610 (.A(n_31849),
    .B(n_33788),
    .Y(n_31850));
 AOI211xp5_ASAP7_75t_SL g184613 (.A1(n_8124),
    .A2(n_25405),
    .B(n_4401),
    .C(n_31864),
    .Y(n_31865));
 AND2x2_ASAP7_75t_R g184614 (.A(out_slt3[14]),
    .B(n_5024),
    .Y(n_31864));
 AOI211xp5_ASAP7_75t_SL g184615 (.A1(n_46336),
    .A2(n_25405),
    .B(n_4404),
    .C(n_31866),
    .Y(n_31867));
 AND2x2_ASAP7_75t_R g184616 (.A(out_slt3[15]),
    .B(n_4513),
    .Y(n_31866));
 AND2x4_ASAP7_75t_SL g184622 (.A(u5_rp[1]),
    .B(n_14010),
    .Y(n_31888));
 AOI22xp5_ASAP7_75t_SL g184623 (.A1(\u5_mem[0] [11]),
    .A2(n_53101),
    .B1(n_64833),
    .B2(\u5_mem[1] [11]),
    .Y(n_31890));
 AOI22xp5_ASAP7_75t_SL g184625 (.A1(n_53101),
    .A2(\u5_mem[0] [5]),
    .B1(n_64833),
    .B2(\u5_mem[1] [5]),
    .Y(n_31891));
 AOI22xp5_ASAP7_75t_SL g184626 (.A1(n_53101),
    .A2(\u5_mem[0] [7]),
    .B1(n_64833),
    .B2(\u5_mem[1] [7]),
    .Y(n_31892));
 BUFx3_ASAP7_75t_SL g184630 (.A(n_31888),
    .Y(n_31895));
 AOI22xp33_ASAP7_75t_SL g184634 (.A1(n_65642),
    .A2(\u5_mem[0] [13]),
    .B1(n_64833),
    .B2(\u5_mem[1] [13]),
    .Y(n_31900));
 AOI22xp5_ASAP7_75t_SL g184641 (.A1(n_64833),
    .A2(\u5_mem[1] [4]),
    .B1(n_53101),
    .B2(\u5_mem[0] [4]),
    .Y(n_31907));
 AND2x4_ASAP7_75t_L g184750 (.A(n_675),
    .B(n_32162),
    .Y(n_32163));
 INVx2_ASAP7_75t_SL g184751 (.A(n_379),
    .Y(n_675));
 AND2x2_ASAP7_75t_SL g184752 (.A(u5_wp[0]),
    .B(o6_we),
    .Y(n_32162));
 NAND2x1p5_ASAP7_75t_SL g184861 (.A(n_33604),
    .B(u10_wp[1]),
    .Y(n_32299));
 INVx1_ASAP7_75t_SL g184862 (.A(n_234),
    .Y(n_32300));
 NAND3x2_ASAP7_75t_SL g184873 (.B(wb_addr_i[4]),
    .C(wb_addr_i[2]),
    .Y(n_32317),
    .A(n_8177));
 AOI22xp5_ASAP7_75t_SL g184874 (.A1(n_66842),
    .A2(n_6732),
    .B1(n_290),
    .B2(n_32319),
    .Y(n_32320));
 OR2x6_ASAP7_75t_SL g184875 (.A(n_32318),
    .B(n_32317),
    .Y(n_32319));
 INVx2_ASAP7_75t_SL g184876 (.A(rf_we),
    .Y(n_32318));
 AOI22xp5_ASAP7_75t_SL g184877 (.A1(n_10924),
    .A2(n_6732),
    .B1(u13_intm_r[0]),
    .B2(n_32319),
    .Y(n_32321));
 AOI22xp5_ASAP7_75t_SL g184878 (.A1(n_78044),
    .A2(n_6732),
    .B1(n_19002),
    .B2(n_32319),
    .Y(n_32322));
 AOI22xp5_ASAP7_75t_SL g184879 (.A1(n_65908),
    .A2(n_6748),
    .B1(u13_intm_r[27]),
    .B2(n_32319),
    .Y(n_32323));
 AOI22xp5_ASAP7_75t_SL g184880 (.A1(n_66010),
    .A2(n_6748),
    .B1(n_24637),
    .B2(n_32319),
    .Y(n_32324));
 AOI22xp5_ASAP7_75t_SL g184881 (.A1(n_28316),
    .A2(n_6748),
    .B1(u13_intm_r[25]),
    .B2(n_32319),
    .Y(n_32325));
 AOI22xp5_ASAP7_75t_SL g184882 (.A1(n_28424),
    .A2(n_6748),
    .B1(n_227),
    .B2(n_32319),
    .Y(n_32326));
 AOI22xp5_ASAP7_75t_SL g184883 (.A1(n_22640),
    .A2(n_6748),
    .B1(u13_intm_r[28]),
    .B2(n_32319),
    .Y(n_32327));
 AOI22xp5_ASAP7_75t_SL g184884 (.A1(n_65930),
    .A2(n_6748),
    .B1(n_312),
    .B2(n_32319),
    .Y(n_32328));
 AOI22xp5_ASAP7_75t_SL g184886 (.A1(n_73996),
    .A2(n_6748),
    .B1(u13_intm_r[21]),
    .B2(n_32319),
    .Y(n_32330));
 AOI22xp5_ASAP7_75t_SL g184887 (.A1(n_66026),
    .A2(n_6748),
    .B1(u13_intm_r[20]),
    .B2(n_32319),
    .Y(n_32331));
 AOI22xp5_ASAP7_75t_SL g184888 (.A1(n_10196),
    .A2(n_6748),
    .B1(n_291),
    .B2(n_32319),
    .Y(n_32332));
 AOI22xp5_ASAP7_75t_SL g184889 (.A1(n_65934),
    .A2(n_6748),
    .B1(n_223),
    .B2(n_32319),
    .Y(n_32333));
 AOI22xp5_ASAP7_75t_SL g184890 (.A1(n_65952),
    .A2(n_6748),
    .B1(u13_intm_r[17]),
    .B2(n_32319),
    .Y(n_32334));
 AOI22xp5_ASAP7_75t_SL g184891 (.A1(n_28276),
    .A2(n_6748),
    .B1(u13_intm_r[16]),
    .B2(n_32335),
    .Y(n_32336));
 AOI22xp5_ASAP7_75t_SL g184892 (.A1(n_65955),
    .A2(n_6732),
    .B1(n_319),
    .B2(n_32335),
    .Y(n_32337));
 AOI22xp5_ASAP7_75t_SL g184893 (.A1(n_66868),
    .A2(n_6732),
    .B1(u13_intm_r[5]),
    .B2(n_32335),
    .Y(n_32338));
 AOI22xp5_ASAP7_75t_SL g184894 (.A1(n_10026),
    .A2(n_6732),
    .B1(u13_intm_r[12]),
    .B2(n_32335),
    .Y(n_32339));
 AOI22xp5_ASAP7_75t_SL g184896 (.A1(n_79971),
    .A2(n_6732),
    .B1(n_206),
    .B2(n_32335),
    .Y(n_32341));
 AOI22xp5_ASAP7_75t_SL g184898 (.A1(n_28240),
    .A2(n_6732),
    .B1(n_301),
    .B2(n_32335),
    .Y(n_32343));
 AOI22xp5_ASAP7_75t_SL g184899 (.A1(n_28330),
    .A2(n_6732),
    .B1(u13_intm_r[2]),
    .B2(n_32335),
    .Y(n_32344));
 AOI22xp5_ASAP7_75t_SL g184900 (.A1(n_17578),
    .A2(n_6732),
    .B1(u13_intm_r[7]),
    .B2(n_32335),
    .Y(n_32345));
 AOI22xp5_ASAP7_75t_SL g184901 (.A1(n_65990),
    .A2(n_6748),
    .B1(u13_intm_r[15]),
    .B2(n_32335),
    .Y(n_32346));
 AOI22xp5_ASAP7_75t_SL g184903 (.A1(n_32650),
    .A2(n_6732),
    .B1(n_310),
    .B2(n_32335),
    .Y(n_32348));
 AOI22xp5_ASAP7_75t_SL g184904 (.A1(n_66856),
    .A2(n_6732),
    .B1(n_317),
    .B2(n_32335),
    .Y(n_32349));
 AND2x2_ASAP7_75t_SL g184935 (.A(u9_rp[0]),
    .B(u9_rp[1]),
    .Y(n_32381));
 AOI22xp33_ASAP7_75t_SL g184936 (.A1(n_1171),
    .A2(\u9_mem[1] [17]),
    .B1(n_32382),
    .B2(\u9_mem[3] [17]),
    .Y(n_32383));
 AOI22xp33_ASAP7_75t_SL g184938 (.A1(n_1171),
    .A2(\u9_mem[1] [11]),
    .B1(n_32382),
    .B2(\u9_mem[3] [11]),
    .Y(n_32384));
 AOI22xp33_ASAP7_75t_SL g184939 (.A1(n_1171),
    .A2(\u9_mem[1] [1]),
    .B1(n_32382),
    .B2(\u9_mem[3] [1]),
    .Y(n_32385));
 AOI22xp33_ASAP7_75t_SL g184940 (.A1(n_1171),
    .A2(\u9_mem[1] [15]),
    .B1(n_32382),
    .B2(\u9_mem[3] [15]),
    .Y(n_32386));
 AOI22xp33_ASAP7_75t_SL g184941 (.A1(n_1171),
    .A2(\u9_mem[1] [3]),
    .B1(n_32382),
    .B2(\u9_mem[3] [3]),
    .Y(n_32387));
 AOI22xp33_ASAP7_75t_SL g184942 (.A1(n_1171),
    .A2(\u9_mem[1] [29]),
    .B1(n_32382),
    .B2(\u9_mem[3] [29]),
    .Y(n_32388));
 AOI22xp33_ASAP7_75t_SL g184943 (.A1(n_1171),
    .A2(\u9_mem[1] [2]),
    .B1(n_32382),
    .B2(\u9_mem[3] [2]),
    .Y(n_32389));
 AOI22xp33_ASAP7_75t_SL g184944 (.A1(n_1171),
    .A2(\u9_mem[1] [30]),
    .B1(n_32382),
    .B2(\u9_mem[3] [30]),
    .Y(n_32390));
 AOI22xp33_ASAP7_75t_SL g184945 (.A1(n_1171),
    .A2(\u9_mem[1] [21]),
    .B1(n_32382),
    .B2(\u9_mem[3] [21]),
    .Y(n_32391));
 AOI22xp33_ASAP7_75t_SL g184946 (.A1(n_1171),
    .A2(\u9_mem[1] [18]),
    .B1(n_32382),
    .B2(\u9_mem[3] [18]),
    .Y(n_32392));
 AOI22xp33_ASAP7_75t_SL g184947 (.A1(n_1171),
    .A2(\u9_mem[1] [4]),
    .B1(n_32382),
    .B2(\u9_mem[3] [4]),
    .Y(n_32393));
 AOI22xp33_ASAP7_75t_SL g184948 (.A1(n_1171),
    .A2(\u9_mem[1] [25]),
    .B1(n_32382),
    .B2(\u9_mem[3] [25]),
    .Y(n_32394));
 AOI22xp33_ASAP7_75t_SL g184949 (.A1(n_1171),
    .A2(\u9_mem[1] [9]),
    .B1(n_32382),
    .B2(\u9_mem[3] [9]),
    .Y(n_32395));
 AOI22xp33_ASAP7_75t_SL g184950 (.A1(n_1171),
    .A2(\u9_mem[1] [24]),
    .B1(n_32382),
    .B2(\u9_mem[3] [24]),
    .Y(n_32396));
 AOI22xp33_ASAP7_75t_SL g184951 (.A1(n_1171),
    .A2(\u9_mem[1] [28]),
    .B1(n_22780),
    .B2(\u9_mem[3] [28]),
    .Y(n_32398));
 AOI22xp33_ASAP7_75t_SL g184952 (.A1(n_1171),
    .A2(\u9_mem[1] [6]),
    .B1(n_22780),
    .B2(\u9_mem[3] [6]),
    .Y(n_32399));
 AOI22xp33_ASAP7_75t_SL g184953 (.A1(n_1171),
    .A2(\u9_mem[1] [31]),
    .B1(n_22780),
    .B2(\u9_mem[3] [31]),
    .Y(n_32400));
 AOI22xp33_ASAP7_75t_SL g184954 (.A1(n_1171),
    .A2(\u9_mem[1] [23]),
    .B1(n_22780),
    .B2(\u9_mem[3] [23]),
    .Y(n_32401));
 AOI22xp33_ASAP7_75t_SL g184955 (.A1(n_1171),
    .A2(\u9_mem[1] [5]),
    .B1(n_22780),
    .B2(\u9_mem[3] [5]),
    .Y(n_32402));
 AOI22xp33_ASAP7_75t_SL g184956 (.A1(n_1171),
    .A2(\u9_mem[1] [20]),
    .B1(n_22780),
    .B2(\u9_mem[3] [20]),
    .Y(n_32403));
 AOI22xp33_ASAP7_75t_SL g184957 (.A1(n_1171),
    .A2(\u9_mem[1] [13]),
    .B1(n_22780),
    .B2(\u9_mem[3] [13]),
    .Y(n_32404));
 AOI22xp33_ASAP7_75t_SL g184958 (.A1(n_1171),
    .A2(\u9_mem[1] [26]),
    .B1(n_22780),
    .B2(\u9_mem[3] [26]),
    .Y(n_32405));
 AOI22xp33_ASAP7_75t_SL g184959 (.A1(n_1171),
    .A2(\u9_mem[1] [12]),
    .B1(n_22780),
    .B2(\u9_mem[3] [12]),
    .Y(n_32406));
 AOI22xp33_ASAP7_75t_SL g184960 (.A1(n_1171),
    .A2(\u9_mem[1] [27]),
    .B1(n_22780),
    .B2(\u9_mem[3] [27]),
    .Y(n_32407));
 AOI22xp33_ASAP7_75t_SL g184961 (.A1(n_1171),
    .A2(\u9_mem[1] [10]),
    .B1(n_22780),
    .B2(\u9_mem[3] [10]),
    .Y(n_32408));
 AOI22xp33_ASAP7_75t_SL g184962 (.A1(n_1171),
    .A2(\u9_mem[1] [8]),
    .B1(n_22780),
    .B2(\u9_mem[3] [8]),
    .Y(n_32409));
 AOI22xp33_ASAP7_75t_SL g184963 (.A1(n_1171),
    .A2(\u9_mem[1] [16]),
    .B1(n_22780),
    .B2(\u9_mem[3] [16]),
    .Y(n_32410));
 AOI22xp33_ASAP7_75t_SL g184964 (.A1(n_1171),
    .A2(\u9_mem[1] [0]),
    .B1(n_22780),
    .B2(\u9_mem[3] [0]),
    .Y(n_32411));
 INVxp33_ASAP7_75t_R g185 (.A(wb_data_i[11]),
    .Y(n_65964));
 AND2x4_ASAP7_75t_SL g185112 (.A(n_26379),
    .B(n_7766),
    .Y(n_32582));
 AOI211xp5_ASAP7_75t_SL g185115 (.A1(n_16743),
    .A2(n_32582),
    .B(n_4562),
    .C(n_7788),
    .Y(n_32587));
 AOI21xp5_ASAP7_75t_SL g185116 (.A1(n_28443),
    .A2(n_32585),
    .B(n_14917),
    .Y(n_32588));
 AOI211xp5_ASAP7_75t_SL g185119 (.A1(n_36014),
    .A2(n_32582),
    .B(n_4557),
    .C(n_7502),
    .Y(n_32591));
 AOI211xp5_ASAP7_75t_SL g185120 (.A1(n_36010),
    .A2(n_32582),
    .B(n_4549),
    .C(n_7426),
    .Y(n_32592));
 AOI22xp5_ASAP7_75t_SL g185123 (.A1(n_32582),
    .A2(n_27521),
    .B1(n_14926),
    .B2(n_14925),
    .Y(n_32595));
 AOI211xp5_ASAP7_75t_SL g185125 (.A1(n_30332),
    .A2(n_32582),
    .B(n_7800),
    .C(n_7725),
    .Y(n_32597));
 AOI211xp5_ASAP7_75t_SL g185127 (.A1(n_46486),
    .A2(n_32582),
    .B(n_15082),
    .C(n_7586),
    .Y(n_32599));
 AOI211xp5_ASAP7_75t_SL g185129 (.A1(n_7588),
    .A2(n_32582),
    .B(n_4574),
    .C(n_7589),
    .Y(n_32601));
 AND2x2_ASAP7_75t_SL g185545 (.A(u7_wp[0]),
    .B(o8_we),
    .Y(n_33100));
 OAI21xp5_ASAP7_75t_SL g185556 (.A1(n_43535),
    .A2(n_23504),
    .B(n_549),
    .Y(n_33112));
 AND2x2_ASAP7_75t_SL g185961 (.A(u10_wp[1]),
    .B(n_32300),
    .Y(n_33603));
 AND2x4_ASAP7_75t_SL g185962 (.A(n_709),
    .B(n_41767),
    .Y(n_33604));
 INVxp33_ASAP7_75t_R g186 (.A(wb_data_i[27]),
    .Y(n_65905));
 INVx1_ASAP7_75t_SL g186001 (.A(u14_u4_en_out_l2),
    .Y(n_33644));
 AND3x4_ASAP7_75t_SL g186009 (.A(n_29787),
    .B(n_35902),
    .C(o4_we),
    .Y(n_33654));
 AOI22xp5_ASAP7_75t_SL g186010 (.A1(n_29790),
    .A2(n_65915),
    .B1(\u4_mem[0] [24]),
    .B2(n_33655),
    .Y(n_33656));
 INVx3_ASAP7_75t_SL g186011 (.A(n_33654),
    .Y(n_33655));
 AOI22xp5_ASAP7_75t_SL g186012 (.A1(n_29790),
    .A2(n_10194),
    .B1(\u4_mem[0] [18]),
    .B2(n_33657),
    .Y(n_33658));
 INVx3_ASAP7_75t_SL g186013 (.A(n_33654),
    .Y(n_33657));
 AOI22xp5_ASAP7_75t_SL g186014 (.A1(n_29790),
    .A2(n_35041),
    .B1(\u4_mem[0] [13]),
    .B2(n_33657),
    .Y(n_33659));
 AOI22xp5_ASAP7_75t_SL g186015 (.A1(n_29790),
    .A2(n_66000),
    .B1(\u4_mem[0] [2]),
    .B2(n_33657),
    .Y(n_33660));
 AOI22xp33_ASAP7_75t_SL g186016 (.A1(n_29790),
    .A2(n_28251),
    .B1(\u4_mem[0] [14]),
    .B2(n_33657),
    .Y(n_33661));
 AOI22xp5_ASAP7_75t_SL g186017 (.A1(n_29790),
    .A2(n_28381),
    .B1(\u4_mem[0] [23]),
    .B2(n_33657),
    .Y(n_33662));
 AOI22xp5_ASAP7_75t_SL g186018 (.A1(n_29790),
    .A2(n_10247),
    .B1(\u4_mem[0] [20]),
    .B2(n_33657),
    .Y(n_33663));
 AOI22xp5_ASAP7_75t_SL g186019 (.A1(n_29790),
    .A2(n_10143),
    .B1(\u4_mem[0] [17]),
    .B2(n_33657),
    .Y(n_33664));
 AOI22xp5_ASAP7_75t_SL g186020 (.A1(n_65949),
    .A2(n_29790),
    .B1(\u4_mem[0] [16]),
    .B2(n_33657),
    .Y(n_33665));
 AOI22xp5_ASAP7_75t_SL g186021 (.A1(n_29790),
    .A2(n_65997),
    .B1(\u4_mem[0] [12]),
    .B2(n_33657),
    .Y(n_33666));
 AOI22xp5_ASAP7_75t_SL g186022 (.A1(n_66843),
    .A2(n_29790),
    .B1(\u4_mem[0] [11]),
    .B2(n_33657),
    .Y(n_33667));
 AOI22xp5_ASAP7_75t_SL g186023 (.A1(n_29790),
    .A2(n_79971),
    .B1(\u4_mem[0] [9]),
    .B2(n_33657),
    .Y(n_33668));
 AOI22xp5_ASAP7_75t_SL g186025 (.A1(n_29790),
    .A2(n_28240),
    .B1(\u4_mem[0] [8]),
    .B2(n_33657),
    .Y(n_33670));
 AOI22xp5_ASAP7_75t_SL g186026 (.A1(n_29790),
    .A2(n_66855),
    .B1(\u4_mem[0] [3]),
    .B2(n_33657),
    .Y(n_33671));
 AOI22xp5_ASAP7_75t_SL g186027 (.A1(n_29790),
    .A2(n_17578),
    .B1(\u4_mem[0] [7]),
    .B2(n_33657),
    .Y(n_33672));
 AOI22xp5_ASAP7_75t_SL g186028 (.A1(n_29790),
    .A2(n_28913),
    .B1(\u4_mem[0] [15]),
    .B2(n_33657),
    .Y(n_33673));
 AOI22xp5_ASAP7_75t_SL g186029 (.A1(n_29790),
    .A2(n_10640),
    .B1(\u4_mem[0] [30]),
    .B2(n_33655),
    .Y(n_33674));
 AOI22xp5_ASAP7_75t_SL g186030 (.A1(n_29790),
    .A2(n_62940),
    .B1(\u4_mem[0] [27]),
    .B2(n_33655),
    .Y(n_33675));
 AOI22xp5_ASAP7_75t_SL g186031 (.A1(n_29790),
    .A2(n_35437),
    .B1(\u4_mem[0] [26]),
    .B2(n_33655),
    .Y(n_33676));
 AOI22xp5_ASAP7_75t_SL g186032 (.A1(n_29790),
    .A2(n_28316),
    .B1(\u4_mem[0] [25]),
    .B2(n_33655),
    .Y(n_33677));
 AOI22xp5_ASAP7_75t_SL g186033 (.A1(n_29790),
    .A2(n_22640),
    .B1(\u4_mem[0] [28]),
    .B2(n_33655),
    .Y(n_33678));
 AOI22xp5_ASAP7_75t_SL g186034 (.A1(n_29790),
    .A2(n_65902),
    .B1(\u4_mem[0] [31]),
    .B2(n_33655),
    .Y(n_33679));
 AOI22xp5_ASAP7_75t_SL g186036 (.A1(n_29790),
    .A2(n_66016),
    .B1(\u4_mem[0] [21]),
    .B2(n_33655),
    .Y(n_33681));
 AOI22xp5_ASAP7_75t_SL g186037 (.A1(n_29790),
    .A2(n_10196),
    .B1(\u4_mem[0] [19]),
    .B2(n_33655),
    .Y(n_33682));
 AOI22xp5_ASAP7_75t_SL g186038 (.A1(n_29790),
    .A2(n_10058),
    .B1(\u4_mem[0] [5]),
    .B2(n_33655),
    .Y(n_33683));
 AOI22xp5_ASAP7_75t_SL g186039 (.A1(n_29790),
    .A2(n_10924),
    .B1(\u4_mem[0] [0]),
    .B2(n_33655),
    .Y(n_33684));
 AOI22xp5_ASAP7_75t_SL g186040 (.A1(n_29790),
    .A2(n_10891),
    .B1(\u4_mem[0] [1]),
    .B2(n_33655),
    .Y(n_33685));
 AOI22xp5_ASAP7_75t_SL g186041 (.A1(n_29790),
    .A2(n_15952),
    .B1(\u4_mem[0] [29]),
    .B2(n_33655),
    .Y(n_33686));
 AOI22xp5_ASAP7_75t_SL g186042 (.A1(n_29790),
    .A2(n_66004),
    .B1(\u4_mem[0] [6]),
    .B2(n_33655),
    .Y(n_33687));
 OR2x6_ASAP7_75t_SL g186104 (.A(n_30453),
    .B(n_33771),
    .Y(n_33772));
 INVx2_ASAP7_75t_SL g186105 (.A(u7_wp[1]),
    .Y(n_33771));
 INVx2_ASAP7_75t_SL g186107 (.A(n_33771),
    .Y(n_33774));
 OR2x6_ASAP7_75t_SL g186110 (.A(n_33771),
    .B(n_30453),
    .Y(n_33777));
 AOI22xp33_ASAP7_75t_SL g186118 (.A1(\u3_mem[1] [5]),
    .A2(n_71971),
    .B1(\u3_mem[3] [5]),
    .B2(n_71972),
    .Y(n_33786));
 AOI22xp5_ASAP7_75t_SL g186120 (.A1(\u3_mem[0] [11]),
    .A2(n_43318),
    .B1(n_71971),
    .B2(\u3_mem[1] [11]),
    .Y(n_33787));
 AOI22xp5_ASAP7_75t_SL g186121 (.A1(\u3_mem[1] [14]),
    .A2(n_71971),
    .B1(\u3_mem[0] [14]),
    .B2(n_43318),
    .Y(n_33788));
 AOI22xp5_ASAP7_75t_SL g186122 (.A1(\u3_mem[0] [1]),
    .A2(n_43318),
    .B1(\u3_mem[1] [1]),
    .B2(n_71971),
    .Y(n_33789));
 AOI22xp5_ASAP7_75t_SL g186123 (.A1(\u3_mem[0] [15]),
    .A2(n_43318),
    .B1(\u3_mem[1] [15]),
    .B2(n_71971),
    .Y(n_33790));
 AOI22xp5_ASAP7_75t_SL g186124 (.A1(\u3_mem[1] [10]),
    .A2(n_71971),
    .B1(\u3_mem[3] [10]),
    .B2(n_71972),
    .Y(n_33791));
 AOI22xp5_ASAP7_75t_SL g186125 (.A1(\u3_mem[1] [12]),
    .A2(n_71971),
    .B1(\u3_mem[3] [12]),
    .B2(n_71972),
    .Y(n_33792));
 AOI22xp5_ASAP7_75t_SL g186126 (.A1(n_71971),
    .A2(\u3_mem[1] [13]),
    .B1(\u3_mem[3] [13]),
    .B2(n_71972),
    .Y(n_33793));
 HB1xp67_ASAP7_75t_SL g186129 (.A(n_71971),
    .Y(n_33795));
 AOI211xp5_ASAP7_75t_SL g186369 (.A1(n_357),
    .A2(in_slt1[10]),
    .B(n_34081),
    .C(n_388),
    .Y(n_34082));
 INVx1_ASAP7_75t_SL g186370 (.A(n_195),
    .Y(n_34081));
 AOI22xp33_ASAP7_75t_SL g186388 (.A1(n_58959),
    .A2(\u4_mem[0] [13]),
    .B1(n_50709),
    .B2(\u4_mem[1] [13]),
    .Y(n_34098));
 AOI22xp5_ASAP7_75t_SL g186389 (.A1(n_35632),
    .A2(\u4_mem[2] [13]),
    .B1(\u4_mem[3] [13]),
    .B2(n_30078),
    .Y(n_34099));
 NAND2xp5_ASAP7_75t_SL g186390 (.A(n_37052),
    .B(n_24350),
    .Y(n_34102));
 NAND2x1_ASAP7_75t_SL g186474 (.A(n_78945),
    .B(n_48405),
    .Y(n_34190));
 NAND2x1_ASAP7_75t_SL g186487 (.A(n_78940),
    .B(n_12053),
    .Y(n_34203));
 AND2x2_ASAP7_75t_SL g186515 (.A(n_34234),
    .B(n_4027),
    .Y(n_34235));
 NOR3x1_ASAP7_75t_SL g186516 (.A(n_43082),
    .B(n_3468),
    .C(n_57965),
    .Y(n_34234));
 AOI21xp33_ASAP7_75t_SL g186598 (.A1(u10_din_tmp1[8]),
    .A2(n_34420),
    .B(n_34362),
    .Y(n_34363));
 NOR2xp33_ASAP7_75t_SL g186599 (.A(n_29883),
    .B(n_26819),
    .Y(n_34362));
 AOI21xp33_ASAP7_75t_SL g186613 (.A1(u10_din_tmp1[12]),
    .A2(n_34420),
    .B(n_34377),
    .Y(n_34378));
 NOR2xp33_ASAP7_75t_SL g186614 (.A(n_29883),
    .B(n_26807),
    .Y(n_34377));
 AOI21xp33_ASAP7_75t_SL g186648 (.A1(u10_din_tmp1[11]),
    .A2(n_34420),
    .B(n_34412),
    .Y(n_34413));
 NOR2xp33_ASAP7_75t_SL g186649 (.A(n_29883),
    .B(n_14288),
    .Y(n_34412));
 INVx3_ASAP7_75t_SL g186656 (.A(n_29881),
    .Y(n_34420));
 AOI21xp33_ASAP7_75t_SL g186657 (.A1(u10_din_tmp1[6]),
    .A2(n_34420),
    .B(n_34421),
    .Y(n_34422));
 NOR2xp33_ASAP7_75t_SL g186658 (.A(n_29883),
    .B(n_26823),
    .Y(n_34421));
 AND2x2_ASAP7_75t_SL g186669 (.A(n_51032),
    .B(n_34433),
    .Y(n_34434));
 AOI22xp33_ASAP7_75t_SL g186670 (.A1(n_49129),
    .A2(\u7_mem[0] [6]),
    .B1(n_49617),
    .B2(\u7_mem[1] [6]),
    .Y(n_34433));
 AND2x4_ASAP7_75t_SL g186702 (.A(out_slt0[9]),
    .B(n_31581),
    .Y(n_34472));
 INVx1_ASAP7_75t_L g186703 (.A(oc2_cfg[2]),
    .Y(n_34473));
 HB1xp67_ASAP7_75t_L g186708 (.A(n_58649),
    .Y(n_34475));
 INVxp33_ASAP7_75t_R g186709 (.A(n_58649),
    .Y(n_34479));
 INVx1_ASAP7_75t_R g186710 (.A(in_slt6[5]),
    .Y(n_34480));
 NOR2xp33_ASAP7_75t_SL g186713 (.A(n_36289),
    .B(n_34480),
    .Y(n_34482));
 INVxp67_ASAP7_75t_L g186714 (.A(in_slt6[7]),
    .Y(n_34484));
 NOR2xp33_ASAP7_75t_SL g186717 (.A(n_36289),
    .B(n_34484),
    .Y(n_34486));
 INVx1_ASAP7_75t_L g186718 (.A(in_slt3[8]),
    .Y(n_34488));
 NOR2xp33_ASAP7_75t_SL g186721 (.A(n_34505),
    .B(n_34488),
    .Y(n_34490));
 INVx1_ASAP7_75t_R g186722 (.A(in_slt3[13]),
    .Y(n_34492));
 NOR2xp33_ASAP7_75t_SL g186725 (.A(n_34505),
    .B(n_34492),
    .Y(n_34494));
 NOR2xp33_ASAP7_75t_SL g186729 (.A(n_34505),
    .B(n_48052),
    .Y(n_34498));
 INVx1_ASAP7_75t_L g186730 (.A(in_slt3[15]),
    .Y(n_34500));
 NOR2xp33_ASAP7_75t_SL g186733 (.A(n_34505),
    .B(n_34500),
    .Y(n_34502));
 INVx1_ASAP7_75t_R g186734 (.A(in_slt3[17]),
    .Y(n_34504));
 INVx5_ASAP7_75t_SL g186735 (.A(n_31228),
    .Y(n_34505));
 NOR2xp33_ASAP7_75t_SL g186737 (.A(n_34505),
    .B(n_34504),
    .Y(n_34506));
 INVx2_ASAP7_75t_SL g186753 (.A(oc0_cfg[0]),
    .Y(n_34532));
 NAND2xp5_ASAP7_75t_L g186754 (.A(n_34533),
    .B(n_15026),
    .Y(n_34534));
 INVx2_ASAP7_75t_SL g186755 (.A(n_34532),
    .Y(n_34533));
 OAI21xp33_ASAP7_75t_SL g186756 (.A1(n_14432),
    .A2(n_19069),
    .B(n_34535),
    .Y(n_34536));
 INVx1_ASAP7_75t_L g186757 (.A(n_34532),
    .Y(n_34535));
 AND3x1_ASAP7_75t_R g186758 (.A(n_34533),
    .B(n_390),
    .C(n_269),
    .Y(n_34537));
 INVx1_ASAP7_75t_L g186759 (.A(n_34533),
    .Y(n_34538));
 NAND2xp33_ASAP7_75t_L g186760 (.A(n_34533),
    .B(n_608),
    .Y(n_34539));
 INVx1_ASAP7_75t_SL g186761 (.A(n_34535),
    .Y(n_34540));
 OAI21x1_ASAP7_75t_SL g186762 (.A1(n_19133),
    .A2(n_43082),
    .B(n_34535),
    .Y(n_34541));
 AOI21xp33_ASAP7_75t_SL g186830 (.A1(n_34420),
    .A2(u10_din_tmp1[0]),
    .B(n_34613),
    .Y(n_34614));
 NOR2xp67_ASAP7_75t_SL g186831 (.A(n_26859),
    .B(n_34420),
    .Y(n_34613));
 AOI221xp5_ASAP7_75t_SL g186849 (.A1(n_34633),
    .A2(n_32582),
    .B1(n_43087),
    .B2(out_slt4[18]),
    .C(n_4573),
    .Y(n_34634));
 NAND4xp25_ASAP7_75t_SL g186850 (.A(n_50712),
    .B(n_27381),
    .C(n_27382),
    .D(n_27383),
    .Y(n_34633));
 NAND2xp5_ASAP7_75t_SL g186856 (.A(n_34644),
    .B(n_63786),
    .Y(n_34645));
 AOI22xp33_ASAP7_75t_SL g186857 (.A1(n_49129),
    .A2(\u7_mem[0] [14]),
    .B1(\u7_mem[1] [14]),
    .B2(n_49617),
    .Y(n_34644));
 AND2x2_ASAP7_75t_SL g186860 (.A(n_51042),
    .B(n_34648),
    .Y(n_34649));
 AOI22xp33_ASAP7_75t_SL g186861 (.A1(n_49617),
    .A2(\u7_mem[1] [5]),
    .B1(n_49129),
    .B2(\u7_mem[0] [5]),
    .Y(n_34648));
 A2O1A1Ixp33_ASAP7_75t_SL g187013 (.A1(n_34837),
    .A2(n_37136),
    .B(n_48223),
    .C(n_46190),
    .Y(n_34841));
 INVx2_ASAP7_75t_SL g187014 (.A(n_79326),
    .Y(n_34837));
 INVx4_ASAP7_75t_SL g187152 (.A(n_10083),
    .Y(n_35041));
 NOR2x1_ASAP7_75t_L g187220 (.A(n_14280),
    .B(n_1365),
    .Y(n_35120));
 OR2x6_ASAP7_75t_SL g187222 (.A(n_24975),
    .B(n_534),
    .Y(n_35121));
 OR2x6_ASAP7_75t_SL g187310 (.A(n_47780),
    .B(n_29352),
    .Y(n_35215));
 AOI22xp5_ASAP7_75t_SL g187476 (.A1(n_61242),
    .A2(n_35392),
    .B1(\u10_mem[3] [3]),
    .B2(n_61244),
    .Y(n_35393));
 NAND2x1_ASAP7_75t_SL g187477 (.A(n_35390),
    .B(n_35391),
    .Y(n_35392));
 AOI22xp5_ASAP7_75t_SL g187478 (.A1(in_slt4[5]),
    .A2(n_1666),
    .B1(u10_din_tmp1[3]),
    .B2(n_24336),
    .Y(n_35390));
 NAND2xp5_ASAP7_75t_SL g187479 (.A(in_slt4[3]),
    .B(n_1667),
    .Y(n_35391));
 AOI21xp5_ASAP7_75t_SL g187484 (.A1(n_35398),
    .A2(n_28848),
    .B(ic2_int_set[2]),
    .Y(n_35399));
 NOR2xp33_ASAP7_75t_SL g187485 (.A(n_2227),
    .B(n_14319),
    .Y(n_35398));
 NAND2x1_ASAP7_75t_SL g187491 (.A(n_51039),
    .B(n_6295),
    .Y(n_35407));
 INVx3_ASAP7_75t_SL g187520 (.A(n_10460),
    .Y(n_35437));
 INVx2_ASAP7_75t_SL g187538 (.A(n_35457),
    .Y(n_35458));
 BUFx3_ASAP7_75t_SL g187539 (.A(oc1_cfg[3]),
    .Y(n_35457));
 AOI22xp5_ASAP7_75t_SL g187540 (.A1(n_10000),
    .A2(n_67247),
    .B1(n_35459),
    .B2(n_29621),
    .Y(n_35460));
 INVx1_ASAP7_75t_L g187541 (.A(n_35458),
    .Y(n_35459));
 INVx1_ASAP7_75t_SL g187542 (.A(n_35461),
    .Y(n_35462));
 BUFx3_ASAP7_75t_SL g187543 (.A(n_35457),
    .Y(n_35461));
 INVxp67_ASAP7_75t_R g187544 (.A(n_35461),
    .Y(n_35463));
 NAND2xp5_ASAP7_75t_SL g187547 (.A(n_1828),
    .B(n_35459),
    .Y(n_35466));
 NAND2xp5_ASAP7_75t_SL g187548 (.A(n_28441),
    .B(n_35459),
    .Y(n_35467));
 NAND2xp5_ASAP7_75t_SL g187549 (.A(n_35459),
    .B(n_13547),
    .Y(n_35468));
 AOI22xp33_ASAP7_75t_SL g187550 (.A1(n_24350),
    .A2(n_7990),
    .B1(n_35459),
    .B2(n_13822),
    .Y(n_35469));
 OR2x2_ASAP7_75t_R g187553 (.A(u2_res_cnt[2]),
    .B(n_31534),
    .Y(n_35474));
 NAND2xp5_ASAP7_75t_SL g187623 (.A(n_51483),
    .B(n_7538),
    .Y(n_35550));
 INVxp67_ASAP7_75t_R g187653 (.A(n_43100),
    .Y(n_35577));
 NOR5xp2_ASAP7_75t_SL g187654 (.A(n_374),
    .B(n_675),
    .C(n_43100),
    .D(n_2746),
    .E(u5_wp[2]),
    .Y(n_35578));
 AOI22xp5_ASAP7_75t_SL g187708 (.A1(\u4_mem[2] [16]),
    .A2(n_35632),
    .B1(\u4_mem[3] [16]),
    .B2(n_30078),
    .Y(n_35633));
 AND2x6_ASAP7_75t_SL g187709 (.A(u4_rp[2]),
    .B(n_50809),
    .Y(n_35632));
 INVxp67_ASAP7_75t_SL g187711 (.A(n_42621),
    .Y(n_35634));
 INVx1_ASAP7_75t_SL g187712 (.A(u12_re2),
    .Y(n_35636));
 OR3x1_ASAP7_75t_R g187713 (.A(n_35637),
    .B(n_670),
    .C(n_18887),
    .Y(n_35638));
 HB1xp67_ASAP7_75t_SL g187714 (.A(u12_re2),
    .Y(n_35637));
 NAND2xp5_ASAP7_75t_R g187725 (.A(in_slt1[5]),
    .B(oc5_cfg[1]),
    .Y(n_35655));
 AOI22xp5_ASAP7_75t_SL g187726 (.A1(n_79972),
    .A2(n_21311),
    .B1(n_35653),
    .B2(n_26541),
    .Y(n_35654));
 HB1xp67_ASAP7_75t_R g187727 (.A(oc5_cfg[1]),
    .Y(n_35653));
 INVxp67_ASAP7_75t_SL g187728 (.A(oc5_cfg[1]),
    .Y(n_35656));
 INVx2_ASAP7_75t_SL g187960 (.A(u4_wp[1]),
    .Y(n_35902));
 BUFx2_ASAP7_75t_SL g187963 (.A(n_35902),
    .Y(n_35904));
 OR2x6_ASAP7_75t_SL g187966 (.A(n_26050),
    .B(n_35904),
    .Y(n_35908));
 AND2x4_ASAP7_75t_SL g187970_dup198303 (.A(n_48106),
    .B(n_37935),
    .Y(n_48107));
 INVx2_ASAP7_75t_SL g188042 (.A(n_36007),
    .Y(n_36008));
 OR2x2_ASAP7_75t_SL g188043 (.A(oc1_cfg[3]),
    .B(n_71390),
    .Y(n_36007));
 OAI222xp33_ASAP7_75t_SL g188044 (.A1(n_7756),
    .A2(n_26801),
    .B1(n_43305),
    .B2(n_8113),
    .C1(n_50711),
    .C2(n_36007),
    .Y(n_36010));
 OR2x2_ASAP7_75t_SL g188046 (.A(n_415),
    .B(n_36007),
    .Y(n_36011));
 OAI22xp33_ASAP7_75t_R g188047 (.A1(n_8113),
    .A2(n_5691),
    .B1(n_36007),
    .B2(n_5687),
    .Y(n_36012));
 OAI222xp33_ASAP7_75t_SL g188048 (.A1(n_4540),
    .A2(n_26801),
    .B1(n_8111),
    .B2(n_8113),
    .C1(n_2393),
    .C2(n_36007),
    .Y(n_36013));
 OAI222xp33_ASAP7_75t_SL g188049 (.A1(n_46697),
    .A2(n_26801),
    .B1(n_36007),
    .B2(n_13787),
    .C1(n_18679),
    .C2(n_8113),
    .Y(n_36014));
 OR2x2_ASAP7_75t_SL g188058 (.A(n_37456),
    .B(out_slt0[6]),
    .Y(n_36071));
 AOI31xp33_ASAP7_75t_SL g188060 (.A1(n_37456),
    .A2(n_14328),
    .A3(n_1042),
    .B(oc0_int_set[1]),
    .Y(n_36072));
 AND2x2_ASAP7_75t_SL g188061 (.A(n_37457),
    .B(n_37456),
    .Y(n_36073));
 NAND2xp5_ASAP7_75t_SL g188063 (.A(n_37457),
    .B(n_62919),
    .Y(n_36076));
 MAJIxp5_ASAP7_75t_SL g188065 (.A(n_37456),
    .B(n_517),
    .C(n_34082),
    .Y(n_36077));
 AOI22xp33_ASAP7_75t_SL g188066 (.A1(n_3937),
    .A2(n_36078),
    .B1(n_62919),
    .B2(u14_u2_full_empty_r),
    .Y(n_36079));
 MAJIxp5_ASAP7_75t_SL g188068 (.A(n_62919),
    .B(n_181),
    .C(n_1051),
    .Y(n_36080));
 AOI22xp5_ASAP7_75t_SL g188069 (.A1(u14_u1_full_empty_r),
    .A2(n_62919),
    .B1(n_4040),
    .B2(n_36078),
    .Y(n_36081));
 AOI22xp5_ASAP7_75t_SL g188070 (.A1(u14_u3_full_empty_r),
    .A2(n_62919),
    .B1(n_4042),
    .B2(n_36082),
    .Y(n_36083));
 AO21x1_ASAP7_75t_SL g188072 (.A1(n_62919),
    .A2(n_22774),
    .B(n_22775),
    .Y(n_36084));
 AND2x2_ASAP7_75t_SL g188073 (.A(n_62919),
    .B(n_28885),
    .Y(n_36085));
 AOI22xp33_ASAP7_75t_SL g188074 (.A1(u14_u5_full_empty_r),
    .A2(n_62919),
    .B1(o9_empty),
    .B2(n_36078),
    .Y(n_36086));
 NAND2xp5_ASAP7_75t_SL g188077 (.A(out_slt0[11]),
    .B(n_62919),
    .Y(n_36089));
 AOI21xp5_ASAP7_75t_SL g188078 (.A1(n_62919),
    .A2(n_14324),
    .B(n_14326),
    .Y(n_36090));
 AOI31xp33_ASAP7_75t_SL g188079 (.A1(n_62919),
    .A2(n_14345),
    .A3(n_35645),
    .B(oc4_int_set[1]),
    .Y(n_36091));
 NAND2xp5_ASAP7_75t_SL g188080 (.A(n_35645),
    .B(n_62919),
    .Y(n_36092));
 NAND2xp5_ASAP7_75t_SL g188082 (.A(out_slt0[8]),
    .B(n_62919),
    .Y(n_36094));
 AND2x2_ASAP7_75t_SL g188084 (.A(n_1042),
    .B(n_37456),
    .Y(n_36095));
 AOI22xp5_ASAP7_75t_SL g188085 (.A1(out_slt0[13]),
    .A2(n_36078),
    .B1(n_62919),
    .B2(crac_wr),
    .Y(n_36097));
 MAJIxp5_ASAP7_75t_SL g188086 (.A(n_62919),
    .B(n_62918),
    .C(n_43099),
    .Y(n_36098));
 AOI31xp33_ASAP7_75t_SL g188087 (.A1(n_62919),
    .A2(out_slt0[8]),
    .A3(n_28413),
    .B(oc3_int_set[1]),
    .Y(n_36099));
 AOI31xp33_ASAP7_75t_SL g188088 (.A1(n_62919),
    .A2(n_62918),
    .A3(n_14343),
    .B(oc2_int_set[1]),
    .Y(n_36100));
 AOI22xp5_ASAP7_75t_SL g188089 (.A1(u14_u4_full_empty_r),
    .A2(n_62919),
    .B1(n_14350),
    .B2(n_36078),
    .Y(n_36101));
 AOI22xp5_ASAP7_75t_SL g188090 (.A1(u14_u0_full_empty_r),
    .A2(n_62919),
    .B1(n_14333),
    .B2(n_36078),
    .Y(n_36102));
 NAND2xp5_ASAP7_75t_SL g188091 (.A(n_1042),
    .B(n_62919),
    .Y(n_36103));
 NAND2x1_ASAP7_75t_SL g188094 (.A(n_51037),
    .B(n_19501),
    .Y(n_36107));
 NAND2xp5_ASAP7_75t_L g188211 (.A(n_56845),
    .B(n_28294),
    .Y(n_36224));
 INVxp67_ASAP7_75t_R g188258 (.A(in_slt6[11]),
    .Y(n_36288));
 NOR2xp33_ASAP7_75t_SL g188261 (.A(n_36289),
    .B(n_36288),
    .Y(n_36290));
 BUFx3_ASAP7_75t_SL g188330 (.A(n_46182),
    .Y(n_36361));
 NAND2xp5_ASAP7_75t_SL g188331 (.A(out_slt7[5]),
    .B(n_36361),
    .Y(n_36363));
 AND2x2_ASAP7_75t_R g188332 (.A(n_36361),
    .B(out_slt7[16]),
    .Y(n_36364));
 NAND2xp5_ASAP7_75t_SL g188349 (.A(n_36382),
    .B(n_78951),
    .Y(n_36383));
 AOI22xp33_ASAP7_75t_SL g188350 (.A1(n_77853),
    .A2(\u6_mem[2] [2]),
    .B1(n_41152),
    .B2(\u6_mem[3] [2]),
    .Y(n_36382));
 NAND2xp5_ASAP7_75t_SL g188352 (.A(n_12070),
    .B(n_78957),
    .Y(n_36385));
 OA22x2_ASAP7_75t_SL g188414 (.A1(n_26827),
    .A2(n_330),
    .B1(n_14292),
    .B2(n_17606),
    .Y(n_36478));
 NAND2xp5_ASAP7_75t_SL g188460 (.A(n_48412),
    .B(n_78944),
    .Y(n_36525));
 AND2x4_ASAP7_75t_SL g188463 (.A(n_497),
    .B(n_79192),
    .Y(n_36528));
 NAND4xp25_ASAP7_75t_SL g188465 (.A(n_1444),
    .B(n_2444),
    .C(n_1391),
    .D(n_36530),
    .Y(n_36531));
 NAND2xp5_ASAP7_75t_SL g188466 (.A(n_48974),
    .B(n_36528),
    .Y(n_36530));
 INVxp67_ASAP7_75t_SL g188517 (.A(n_24316),
    .Y(n_36580));
 OAI21xp5_ASAP7_75t_SL g188518 (.A1(n_36580),
    .A2(n_36581),
    .B(n_36582),
    .Y(n_36583));
 HB1xp67_ASAP7_75t_SL g188519 (.A(n_33771),
    .Y(n_36581));
 INVxp33_ASAP7_75t_R g188520 (.A(\u7_mem[3] [16]),
    .Y(n_36582));
 AOI22xp5_ASAP7_75t_SL g188525 (.A1(\u4_mem[1] [9]),
    .A2(n_50709),
    .B1(\u4_mem[3] [9]),
    .B2(n_30078),
    .Y(n_36613));
 NAND2xp5_ASAP7_75t_SL g188533 (.A(n_78953),
    .B(n_13974),
    .Y(n_36628));
 AOI22xp5_ASAP7_75t_SL g188542 (.A1(n_64833),
    .A2(\u5_mem[1] [14]),
    .B1(\u5_mem[0] [14]),
    .B2(n_65642),
    .Y(n_36635));
 OAI21xp5_ASAP7_75t_SL g188567 (.A1(n_31535),
    .A2(n_31534),
    .B(u2_res_cnt[2]),
    .Y(n_36662));
 NAND2xp33_ASAP7_75t_SL g188672 (.A(n_78810),
    .B(n_65395),
    .Y(n_36769));
 INVxp33_ASAP7_75t_SL g188676 (.A(n_65395),
    .Y(n_36770));
 NAND2xp5_ASAP7_75t_SL g188677 (.A(n_65395),
    .B(n_78041),
    .Y(n_36771));
 OAI221xp5_ASAP7_75t_SL g188727 (.A1(n_50292),
    .A2(n_34434),
    .B1(n_14959),
    .B2(n_64715),
    .C(n_14961),
    .Y(n_36843));
 NAND2x1_ASAP7_75t_SL g188803 (.A(n_36968),
    .B(n_56860),
    .Y(n_36969));
 AOI22xp5_ASAP7_75t_SL g188804 (.A1(n_65642),
    .A2(\u5_mem[0] [6]),
    .B1(n_64833),
    .B2(\u5_mem[1] [6]),
    .Y(n_36968));
 AND2x2_ASAP7_75t_SL g188886 (.A(n_34098),
    .B(n_34099),
    .Y(n_37051));
 NAND2xp5_ASAP7_75t_SL g188887 (.A(n_34098),
    .B(n_34099),
    .Y(n_37052));
 AOI21x1_ASAP7_75t_SL g188937 (.A1(n_37110),
    .A2(n_34537),
    .B(n_36095),
    .Y(n_37111));
 OR2x2_ASAP7_75t_SL g188938 (.A(n_62919),
    .B(out_slt0[12]),
    .Y(n_37110));
 NAND2xp5_ASAP7_75t_SL g188953 (.A(n_73154),
    .B(n_78041),
    .Y(n_37136));
 NAND4xp25_ASAP7_75t_SL g188955 (.A(n_37137),
    .B(n_37138),
    .C(n_37139),
    .D(n_37136),
    .Y(n_37140));
 AOI22xp33_ASAP7_75t_SL g188956 (.A1(\u6_mem[1] [21]),
    .A2(n_48415),
    .B1(\u6_mem[3] [21]),
    .B2(n_17704),
    .Y(n_37137));
 NAND2xp5_ASAP7_75t_SL g188957 (.A(n_36525),
    .B(n_78810),
    .Y(n_37138));
 AOI22xp33_ASAP7_75t_L g188958 (.A1(\u6_mem[0] [21]),
    .A2(n_79305),
    .B1(\u6_mem[2] [21]),
    .B2(n_79306),
    .Y(n_37139));
 AND2x2_ASAP7_75t_SL g189005 (.A(n_7671),
    .B(n_13405),
    .Y(n_37200));
 INVx2_ASAP7_75t_SL g189094 (.A(n_37336),
    .Y(n_37337));
 NAND2x1_ASAP7_75t_SL g189095 (.A(u6_rp[0]),
    .B(n_37335),
    .Y(n_37336));
 NOR2xp33_ASAP7_75t_R g189097 (.A(n_37336),
    .B(n_77796),
    .Y(n_37338));
 OAI21xp33_ASAP7_75t_SL g189098 (.A1(n_4027),
    .A2(n_37339),
    .B(n_12227),
    .Y(n_37340));
 INVx2_ASAP7_75t_L g189099 (.A(n_37337),
    .Y(n_37339));
 OAI222xp33_ASAP7_75t_SL g189100 (.A1(n_34837),
    .A2(n_6122),
    .B1(n_41154),
    .B2(n_37339),
    .C1(n_31886),
    .C2(n_7442),
    .Y(n_37341));
 OAI211xp5_ASAP7_75t_SL g189101 (.A1(n_70415),
    .A2(n_37339),
    .B(n_14966),
    .C(n_19672),
    .Y(n_37342));
 OAI222xp33_ASAP7_75t_SL g189103 (.A1(n_77855),
    .A2(n_37339),
    .B1(n_37367),
    .B2(n_6138),
    .C1(n_2375),
    .C2(n_7442),
    .Y(n_37344));
 AOI22xp33_ASAP7_75t_L g189110 (.A1(n_79305),
    .A2(\u6_mem[0] [26]),
    .B1(\u6_mem[2] [26]),
    .B2(n_79306),
    .Y(n_37350));
 NAND2x1_ASAP7_75t_SL g189113 (.A(n_78949),
    .B(n_12066),
    .Y(n_37355));
 AND2x2_ASAP7_75t_SL g189123 (.A(n_48407),
    .B(n_78947),
    .Y(n_37367));
 NAND2xp33_ASAP7_75t_SL g189125 (.A(n_78947),
    .B(n_48407),
    .Y(n_37368));
 OAI21xp5_ASAP7_75t_SL g189137 (.A1(n_37381),
    .A2(n_65029),
    .B(n_37383),
    .Y(n_37384));
 INVxp67_ASAP7_75t_R g189138 (.A(\u7_mem[2] [25]),
    .Y(n_37381));
 NAND2xp5_ASAP7_75t_L g189140 (.A(\u7_mem[3] [25]),
    .B(n_73175),
    .Y(n_37383));
 AND2x2_ASAP7_75t_SL g189142 (.A(n_37386),
    .B(n_33604),
    .Y(n_37387));
 INVx1_ASAP7_75t_SL g189143 (.A(n_47767),
    .Y(n_37386));
 AOI21xp5_ASAP7_75t_SL g189208 (.A1(n_37456),
    .A2(n_37459),
    .B(oc5_int_set[1]),
    .Y(n_37460));
 INVx2_ASAP7_75t_SL g189209 (.A(n_43082),
    .Y(n_37456));
 NOR3xp33_ASAP7_75t_L g189210 (.A(n_37458),
    .B(n_2964),
    .C(n_67328),
    .Y(n_37459));
 INVx1_ASAP7_75t_SL g189211 (.A(n_37457),
    .Y(n_37458));
 BUFx3_ASAP7_75t_SL g189212 (.A(out_slt0[6]),
    .Y(n_37457));
 AOI21xp33_ASAP7_75t_SL g189273 (.A1(in_slt1[6]),
    .A2(oc4_cfg[1]),
    .B(n_70326),
    .Y(n_37521));
 AND2x2_ASAP7_75t_SL g189476 (.A(u4_wp[0]),
    .B(o4_we),
    .Y(n_37935));
 AND2x4_ASAP7_75t_SL g189837 (.A(n_28689),
    .B(n_79103),
    .Y(n_38363));
 NAND2xp33_ASAP7_75t_R g189838 (.A(n_66666),
    .B(n_38364),
    .Y(n_38365));
 INVx3_ASAP7_75t_SL g189839 (.A(n_38363),
    .Y(n_38364));
 NAND2xp33_ASAP7_75t_R g189840 (.A(n_66680),
    .B(n_38364),
    .Y(n_38366));
 OAI22xp33_ASAP7_75t_SL g189841 (.A1(n_7270),
    .A2(n_66670),
    .B1(n_4316),
    .B2(n_38364),
    .Y(n_38367));
 NAND2xp33_ASAP7_75t_R g189842 (.A(n_38364),
    .B(n_66682),
    .Y(n_38368));
 A2O1A1Ixp33_ASAP7_75t_SL g189843 (.A1(n_65000),
    .A2(n_65646),
    .B(n_38364),
    .C(n_66677),
    .Y(n_38369));
 NAND2xp33_ASAP7_75t_R g189845 (.A(n_66667),
    .B(n_38364),
    .Y(n_38371));
 NOR2xp33_ASAP7_75t_R g189847 (.A(n_4318),
    .B(n_38364),
    .Y(n_38373));
 A2O1A1Ixp33_ASAP7_75t_SL g189855 (.A1(n_7689),
    .A2(n_73169),
    .B(n_38374),
    .C(n_66669),
    .Y(n_38382));
 AND2x4_ASAP7_75t_SL g19 (.A(n_22851),
    .B(rf_we),
    .Y(n_22852));
 XNOR2xp5_ASAP7_75t_L g190134 (.A(n_13898),
    .B(u6_wp[2]),
    .Y(n_38705));
 A2O1A1Ixp33_ASAP7_75t_SL g190187 (.A1(n_16672),
    .A2(n_2524),
    .B(n_4485),
    .C(n_13955),
    .Y(n_38758));
 MAJIxp5_ASAP7_75t_SL g190188 (.A(n_38759),
    .B(n_62919),
    .C(n_35645),
    .Y(n_38760));
 AND2x2_ASAP7_75t_SL g190189 (.A(n_37521),
    .B(n_491),
    .Y(n_38759));
 AOI21xp5_ASAP7_75t_SL g190190 (.A1(n_49618),
    .A2(u7_rp[0]),
    .B(n_2691),
    .Y(n_38761));
 NAND2x1_ASAP7_75t_SL g191422 (.A(n_40286),
    .B(n_6051),
    .Y(n_40287));
 AOI22xp5_ASAP7_75t_SL g191423 (.A1(\u3_mem[3] [8]),
    .A2(n_71972),
    .B1(\u3_mem[1] [8]),
    .B2(n_43317),
    .Y(n_40286));
 AOI21xp5_ASAP7_75t_SL g191486 (.A1(n_24336),
    .A2(u10_din_tmp1[4]),
    .B(n_40371),
    .Y(n_40372));
 NOR2xp33_ASAP7_75t_L g191487 (.A(n_14292),
    .B(n_330),
    .Y(n_40371));
 AOI21xp5_ASAP7_75t_SL g191491 (.A1(n_24336),
    .A2(u10_din_tmp1[5]),
    .B(n_64697),
    .Y(n_40379));
 INVx1_ASAP7_75t_SL g191527 (.A(u3_wp[0]),
    .Y(n_24373));
 INVx1_ASAP7_75t_SL g191530 (.A(n_24373),
    .Y(n_40418));
 OAI22xp33_ASAP7_75t_SL g191531 (.A1(n_40420),
    .A2(u3_rp[0]),
    .B1(n_417),
    .B2(n_40419),
    .Y(n_40421));
 INVx1_ASAP7_75t_SL g191532 (.A(n_40419),
    .Y(n_40420));
 AOI22xp5_ASAP7_75t_SL g191533 (.A1(n_24373),
    .A2(n_40417),
    .B1(n_40418),
    .B2(n_40416),
    .Y(n_40419));
 NAND2xp5_ASAP7_75t_SL g191781 (.A(n_48631),
    .B(n_50454),
    .Y(n_40712));
 NAND2xp5_ASAP7_75t_SL g191893 (.A(n_40900),
    .B(n_51481),
    .Y(n_40902));
 AOI22xp33_ASAP7_75t_SL g191894 (.A1(n_59474),
    .A2(\u8_mem[0] [0]),
    .B1(n_78274),
    .B2(\u8_mem[1] [0]),
    .Y(n_40900));
 INVxp67_ASAP7_75t_L g191896 (.A(n_40902),
    .Y(n_40904));
 NAND2x1_ASAP7_75t_SL g191944 (.A(n_40954),
    .B(n_40955),
    .Y(n_40956));
 AOI22xp5_ASAP7_75t_SL g191945 (.A1(u10_din_tmp1[0]),
    .A2(n_24336),
    .B1(in_slt4[2]),
    .B2(n_1666),
    .Y(n_40954));
 NAND2xp5_ASAP7_75t_SL g191946 (.A(n_1667),
    .B(in_slt4[0]),
    .Y(n_40955));
 AND2x2_ASAP7_75t_SL g191966 (.A(u8_wp[0]),
    .B(o9_we),
    .Y(n_40978));
 INVx2_ASAP7_75t_L g191967 (.A(n_64814),
    .Y(n_14763));
 AOI22xp5_ASAP7_75t_SL g191970 (.A1(n_28913),
    .A2(n_75734),
    .B1(\u8_mem[1] [15]),
    .B2(n_73399),
    .Y(n_40982));
 AOI22xp5_ASAP7_75t_SL g191971 (.A1(n_10026),
    .A2(n_75734),
    .B1(\u8_mem[1] [12]),
    .B2(n_73399),
    .Y(n_40983));
 AOI22xp5_ASAP7_75t_SL g191973 (.A1(\u8_mem[1] [13]),
    .A2(n_31464),
    .B1(n_65955),
    .B2(n_75734),
    .Y(n_40985));
 AOI22xp5_ASAP7_75t_SL g191974 (.A1(\u8_mem[1] [2]),
    .A2(n_31464),
    .B1(n_66000),
    .B2(n_75734),
    .Y(n_40986));
 AOI22xp5_ASAP7_75t_SL g191975 (.A1(\u8_mem[1] [7]),
    .A2(n_31464),
    .B1(n_17578),
    .B2(n_75734),
    .Y(n_40987));
 AOI22xp5_ASAP7_75t_SL g191976 (.A1(\u8_mem[1] [8]),
    .A2(n_31460),
    .B1(n_65980),
    .B2(n_75734),
    .Y(n_40988));
 AOI22xp5_ASAP7_75t_SL g191977 (.A1(\u8_mem[1] [14]),
    .A2(n_31460),
    .B1(n_28251),
    .B2(n_75734),
    .Y(n_40989));
 AOI22xp5_ASAP7_75t_SL g191978 (.A1(\u8_mem[1] [5]),
    .A2(n_73399),
    .B1(n_66868),
    .B2(n_75734),
    .Y(n_40990));
 AOI22xp5_ASAP7_75t_SL g191980 (.A1(n_66842),
    .A2(n_75734),
    .B1(\u8_mem[1] [11]),
    .B2(n_75735),
    .Y(n_40992));
 AOI22xp5_ASAP7_75t_SL g191981 (.A1(n_75734),
    .A2(n_3815),
    .B1(\u8_mem[1] [1]),
    .B2(n_73399),
    .Y(n_40993));
 OAI21xp5_ASAP7_75t_SL g191982 (.A1(n_75734),
    .A2(n_17545),
    .B(n_556),
    .Y(n_40994));
 AOI22xp5_ASAP7_75t_L g192019 (.A1(\u3_mem[1] [6]),
    .A2(n_43317),
    .B1(\u3_mem[3] [6]),
    .B2(n_71972),
    .Y(n_41034));
 AND2x6_ASAP7_75t_SL g192138 (.A(u6_rp[1]),
    .B(u6_rp[2]),
    .Y(n_41152));
 AND2x2_ASAP7_75t_SL g192139 (.A(n_78946),
    .B(n_48423),
    .Y(n_41154));
 NAND2xp5_ASAP7_75t_SL g192278 (.A(n_31445),
    .B(n_37200),
    .Y(n_41323));
 OAI22xp33_ASAP7_75t_SL g192329 (.A1(n_1892),
    .A2(n_41376),
    .B1(n_23529),
    .B2(n_41377),
    .Y(n_41378));
 INVx1_ASAP7_75t_SL g192330 (.A(n_41375),
    .Y(n_41376));
 HB1xp67_ASAP7_75t_SL g192331 (.A(n_48105),
    .Y(n_41375));
 HB1xp67_ASAP7_75t_L g192332 (.A(n_41375),
    .Y(n_41377));
 AOI22xp33_ASAP7_75t_SL g192333 (.A1(n_31770),
    .A2(n_41377),
    .B1(n_29659),
    .B2(n_35910),
    .Y(n_41379));
 NAND2xp5_ASAP7_75t_SL g192383 (.A(n_36528),
    .B(n_78276),
    .Y(n_41435));
 INVx1_ASAP7_75t_SL g192437 (.A(n_41491),
    .Y(n_41492));
 NAND2x1_ASAP7_75t_SL g192438 (.A(n_6297),
    .B(n_51033),
    .Y(n_41491));
 AOI22xp5_ASAP7_75t_SL g192552 (.A1(n_50388),
    .A2(\u3_mem[2] [11]),
    .B1(\u3_mem[3] [11]),
    .B2(n_71972),
    .Y(n_41606));
 INVx1_ASAP7_75t_SL g192553 (.A(n_70326),
    .Y(n_41608));
 AO21x1_ASAP7_75t_SL g192554 (.A1(n_24523),
    .A2(n_24524),
    .B(n_41610),
    .Y(n_41611));
 NAND2xp5_ASAP7_75t_SL g192555 (.A(n_41608),
    .B(n_41609),
    .Y(n_41610));
 AND2x2_ASAP7_75t_L g192556 (.A(n_15037),
    .B(oc4_cfg[6]),
    .Y(n_41609));
 AOI21xp33_ASAP7_75t_SL g192557 (.A1(n_24523),
    .A2(n_24524),
    .B(n_41610),
    .Y(n_41612));
 NAND2x1_ASAP7_75t_SL g192579 (.A(n_41636),
    .B(n_56856),
    .Y(n_41637));
 AOI22xp5_ASAP7_75t_SL g192581 (.A1(n_64833),
    .A2(\u5_mem[1] [10]),
    .B1(n_65642),
    .B2(\u5_mem[0] [10]),
    .Y(n_41636));
 AOI21xp5_ASAP7_75t_SL g192700 (.A1(n_41758),
    .A2(n_41759),
    .B(n_43100),
    .Y(n_41761));
 NAND2xp5_ASAP7_75t_SL g192701 (.A(n_19617),
    .B(n_2746),
    .Y(n_41758));
 NAND2xp33_ASAP7_75t_SL g192702 (.A(n_19615),
    .B(o6_we),
    .Y(n_41759));
 NOR2xp33_ASAP7_75t_SL g192709 (.A(n_41767),
    .B(n_41768),
    .Y(n_41769));
 INVx1_ASAP7_75t_SL g192710 (.A(n_12116),
    .Y(n_41767));
 NOR4xp25_ASAP7_75t_SL g192711 (.A(n_2965),
    .B(n_29934),
    .C(u14_u7_full_empty_r),
    .D(n_4075),
    .Y(n_41768));
 INVx2_ASAP7_75t_SL g192845 (.A(u3_wp[0]),
    .Y(n_41910));
 NAND2xp5_ASAP7_75t_SL g192950 (.A(n_42030),
    .B(n_56853),
    .Y(n_42031));
 INVx2_ASAP7_75t_SL g193147 (.A(n_42248),
    .Y(n_42249));
 OA21x2_ASAP7_75t_SL g193148 (.A1(n_70322),
    .A2(n_70325),
    .B(n_331),
    .Y(n_42248));
 NAND2xp5_ASAP7_75t_SL g193149 (.A(out_slt8[10]),
    .B(n_51158),
    .Y(n_42251));
 NAND2xp5_ASAP7_75t_L g193151 (.A(out_slt8[8]),
    .B(n_51158),
    .Y(n_42252));
 NAND2xp5_ASAP7_75t_L g193152 (.A(out_slt8[9]),
    .B(n_42253),
    .Y(n_42254));
 INVx2_ASAP7_75t_SL g193153 (.A(n_42249),
    .Y(n_42253));
 NAND2xp5_ASAP7_75t_SL g193154 (.A(out_slt8[14]),
    .B(n_51158),
    .Y(n_42255));
 NAND2xp5_ASAP7_75t_L g193155 (.A(out_slt8[16]),
    .B(n_51158),
    .Y(n_42256));
 NAND2xp5_ASAP7_75t_L g193156 (.A(out_slt8[17]),
    .B(n_51158),
    .Y(n_42257));
 NAND2xp5_ASAP7_75t_SL g193157 (.A(out_slt8[12]),
    .B(n_51158),
    .Y(n_42258));
 AOI22xp5_ASAP7_75t_SL g193159 (.A1(n_28239),
    .A2(n_49719),
    .B1(out_slt8[0]),
    .B2(n_42253),
    .Y(n_42260));
 AOI221xp5_ASAP7_75t_SL g193162 (.A1(n_22250),
    .A2(n_5077),
    .B1(out_slt8[18]),
    .B2(n_42253),
    .C(n_4384),
    .Y(n_42263));
 HB1xp67_ASAP7_75t_SL g193484 (.A(u26_ps_cnt[0]),
    .Y(n_42613));
 NAND3xp33_ASAP7_75t_SL g193485 (.A(n_42617),
    .B(n_31535),
    .C(n_76054),
    .Y(n_42618));
 OAI22xp33_ASAP7_75t_SL g193486 (.A1(n_42615),
    .A2(n_42613),
    .B1(n_42616),
    .B2(n_76055),
    .Y(n_42617));
 HB1xp67_ASAP7_75t_SL g193487 (.A(n_171),
    .Y(n_42615));
 INVxp67_ASAP7_75t_SL g193488 (.A(n_42615),
    .Y(n_42616));
 AND2x2_ASAP7_75t_SL g193489 (.A(n_42620),
    .B(n_26254),
    .Y(n_42621));
 NOR2xp33_ASAP7_75t_SL g193490 (.A(u12_re2),
    .B(n_42619),
    .Y(n_42620));
 INVxp67_ASAP7_75t_SL g193491 (.A(u12_re1),
    .Y(n_42619));
 AOI22xp5_ASAP7_75t_SL g193552 (.A1(crac_din[6]),
    .A2(n_42722),
    .B1(in_slt2[10]),
    .B2(crac_rd_done),
    .Y(n_42723));
 INVx3_ASAP7_75t_SL g193553 (.A(crac_rd_done),
    .Y(n_42722));
 AOI22xp5_ASAP7_75t_SL g193554 (.A1(crac_din[8]),
    .A2(n_42722),
    .B1(in_slt2[12]),
    .B2(crac_rd_done),
    .Y(n_42724));
 AOI22xp5_ASAP7_75t_SL g193555 (.A1(crac_din[12]),
    .A2(n_42722),
    .B1(in_slt2[16]),
    .B2(crac_rd_done),
    .Y(n_42725));
 AOI22xp5_ASAP7_75t_SL g193556 (.A1(crac_din[14]),
    .A2(n_42722),
    .B1(in_slt2[18]),
    .B2(crac_rd_done),
    .Y(n_42726));
 AOI22xp5_ASAP7_75t_SL g193557 (.A1(crac_din[5]),
    .A2(n_42722),
    .B1(in_slt2[9]),
    .B2(crac_rd_done),
    .Y(n_42727));
 OAI22xp5_ASAP7_75t_SL g193558 (.A1(crac_din[7]),
    .A2(crac_rd_done),
    .B1(n_42722),
    .B2(in_slt2[11]),
    .Y(n_42728));
 AOI22xp33_ASAP7_75t_SL g193559 (.A1(crac_din[13]),
    .A2(n_42729),
    .B1(in_slt2[17]),
    .B2(crac_rd_done),
    .Y(n_42730));
 INVx5_ASAP7_75t_SL g193560 (.A(crac_rd_done),
    .Y(n_42729));
 AOI22xp33_ASAP7_75t_SL g193561 (.A1(crac_din[0]),
    .A2(n_42729),
    .B1(in_slt2[4]),
    .B2(crac_rd_done),
    .Y(n_42731));
 AOI22xp33_ASAP7_75t_SL g193562 (.A1(crac_din[15]),
    .A2(n_42729),
    .B1(in_slt2[19]),
    .B2(crac_rd_done),
    .Y(n_42732));
 AOI22xp33_ASAP7_75t_SL g193563 (.A1(crac_din[1]),
    .A2(n_42729),
    .B1(crac_rd_done),
    .B2(in_slt2[5]),
    .Y(n_42733));
 AOI22xp5_ASAP7_75t_SL g193564 (.A1(crac_din[11]),
    .A2(n_42729),
    .B1(in_slt2[15]),
    .B2(crac_rd_done),
    .Y(n_42734));
 AOI22xp5_ASAP7_75t_SL g193565 (.A1(crac_din[3]),
    .A2(n_42729),
    .B1(in_slt2[7]),
    .B2(crac_rd_done),
    .Y(n_42735));
 INVxp67_ASAP7_75t_SL g193566 (.A(n_42729),
    .Y(n_42736));
 AOI22xp33_ASAP7_75t_SL g193567 (.A1(crac_din[4]),
    .A2(n_42729),
    .B1(in_slt2[8]),
    .B2(crac_rd_done),
    .Y(n_42737));
 AOI22xp33_ASAP7_75t_SL g193568 (.A1(crac_din[10]),
    .A2(n_42729),
    .B1(in_slt2[14]),
    .B2(crac_rd_done),
    .Y(n_42738));
 AOI22xp33_ASAP7_75t_SL g193569 (.A1(crac_din[2]),
    .A2(n_42729),
    .B1(in_slt2[6]),
    .B2(crac_rd_done),
    .Y(n_42739));
 AOI22xp33_ASAP7_75t_SL g193570 (.A1(crac_din[9]),
    .A2(n_42729),
    .B1(in_slt2[13]),
    .B2(crac_rd_done),
    .Y(n_42740));
 INVx2_ASAP7_75t_SL g193607 (.A(n_23526),
    .Y(n_42779));
 OR2x2_ASAP7_75t_R g193622 (.A(n_26815),
    .B(n_330),
    .Y(n_42799));
 AOI31xp33_ASAP7_75t_SL g193853 (.A1(n_43077),
    .A2(n_2692),
    .A3(n_29364),
    .B(oc4_int_set[2]),
    .Y(n_43078));
 AO22x1_ASAP7_75t_SL g193854 (.A1(u7_rp[2]),
    .A2(n_43531),
    .B1(n_33771),
    .B2(n_7656),
    .Y(n_43077));
 INVx4_ASAP7_75t_SL g193857 (.A(n_36068),
    .Y(n_43082));
 INVx1_ASAP7_75t_SL g193858 (.A(n_201),
    .Y(n_43083));
 NAND2xp33_ASAP7_75t_R g193859 (.A(n_43085),
    .B(out_slt4[8]),
    .Y(n_43086));
 OA21x2_ASAP7_75t_SL g193860 (.A1(n_43082),
    .A2(n_43084),
    .B(n_43083),
    .Y(n_43085));
 INVxp67_ASAP7_75t_L g193861 (.A(n_519),
    .Y(n_43084));
 BUFx2_ASAP7_75t_SL g193862 (.A(n_43085),
    .Y(n_43087));
 AOI22xp33_ASAP7_75t_SL g193863 (.A1(n_23129),
    .A2(n_7772),
    .B1(n_43088),
    .B2(out_slt4[12]),
    .Y(n_43089));
 INVx1_ASAP7_75t_SL g193865 (.A(n_43085),
    .Y(n_43090));
 AOI222xp33_ASAP7_75t_SL g193869 (.A1(n_26802),
    .A2(n_29688),
    .B1(n_7772),
    .B2(n_18684),
    .C1(out_slt4[3]),
    .C2(n_43088),
    .Y(n_43094));
 AOI222xp33_ASAP7_75t_SL g193870 (.A1(n_7772),
    .A2(n_8112),
    .B1(n_26802),
    .B2(n_43306),
    .C1(n_43088),
    .C2(out_slt4[2]),
    .Y(n_43095));
 AND2x2_ASAP7_75t_L g193873 (.A(n_78094),
    .B(n_43098),
    .Y(n_43099));
 AOI211xp5_ASAP7_75t_SL g193874 (.A1(oc2_cfg[1]),
    .A2(in_slt1[8]),
    .B(u14_u2_full_empty_r),
    .C(n_4075),
    .Y(n_43098));
 INVx2_ASAP7_75t_SL g193875 (.A(n_78094),
    .Y(n_43100));
 OAI211xp5_ASAP7_75t_SL g193966 (.A1(n_59639),
    .A2(n_43201),
    .B(n_43202),
    .C(n_43203),
    .Y(n_43204));
 AND2x2_ASAP7_75t_L g193968 (.A(n_56845),
    .B(n_28294),
    .Y(n_43201));
 NAND2xp5_ASAP7_75t_SL g193969 (.A(n_7672),
    .B(n_36969),
    .Y(n_43202));
 NAND2xp5_ASAP7_75t_L g193970 (.A(n_49203),
    .B(n_698),
    .Y(n_43203));
 INVx1_ASAP7_75t_SL g193971 (.A(n_36969),
    .Y(n_43205));
 AND2x2_ASAP7_75t_L g194 (.A(n_51048),
    .B(n_19503),
    .Y(n_14959));
 AOI221xp5_ASAP7_75t_SL g194035 (.A1(n_43281),
    .A2(n_5091),
    .B1(n_4988),
    .B2(out_slt9[10]),
    .C(n_4364),
    .Y(n_43282));
 NAND4xp25_ASAP7_75t_SL g194036 (.A(n_2009),
    .B(n_2057),
    .C(n_1389),
    .D(n_1439),
    .Y(n_43281));
 AOI221xp5_ASAP7_75t_SL g194039 (.A1(n_43290),
    .A2(n_25956),
    .B1(n_5062),
    .B2(out_slt7[17]),
    .C(n_4434),
    .Y(n_43291));
 NAND4xp25_ASAP7_75t_SL g194040 (.A(n_30472),
    .B(n_30471),
    .C(n_70414),
    .D(n_30469),
    .Y(n_43290));
 AND2x2_ASAP7_75t_SL g194048 (.A(n_27305),
    .B(n_811),
    .Y(n_43305));
 NAND2xp5_ASAP7_75t_SL g194049 (.A(n_27305),
    .B(n_811),
    .Y(n_43306));
 INVx3_ASAP7_75t_SL g194060 (.A(n_7567),
    .Y(n_43317));
 AND2x4_ASAP7_75t_SL g194061 (.A(n_24586),
    .B(n_40416),
    .Y(n_43318));
 NAND2xp5_ASAP7_75t_SL g194062 (.A(n_43319),
    .B(n_30616),
    .Y(n_43320));
 AOI22xp33_ASAP7_75t_SL g194063 (.A1(n_43317),
    .A2(\u3_mem[1] [2]),
    .B1(n_43318),
    .B2(\u3_mem[0] [2]),
    .Y(n_43319));
 AOI22xp33_ASAP7_75t_SL g194136 (.A1(n_50341),
    .A2(\u3_mem[0] [12]),
    .B1(n_43394),
    .B2(\u3_mem[2] [12]),
    .Y(n_43395));
 OAI21xp5_ASAP7_75t_SL g194197 (.A1(n_1290),
    .A2(n_43467),
    .B(n_43468),
    .Y(n_43469));
 AND2x2_ASAP7_75t_L g194198 (.A(n_178),
    .B(n_1289),
    .Y(n_43467));
 AND2x2_ASAP7_75t_SL g194199 (.A(n_2286),
    .B(n_19578),
    .Y(n_43468));
 INVx2_ASAP7_75t_L g194244 (.A(n_43530),
    .Y(n_43531));
 INVx2_ASAP7_75t_SL g194245 (.A(u7_wp[1]),
    .Y(n_43530));
 OAI31xp33_ASAP7_75t_SL g194246 (.A1(n_36580),
    .A2(n_503),
    .A3(n_65949),
    .B(n_36583),
    .Y(n_43533));
 INVx2_ASAP7_75t_SL g194247 (.A(n_43531),
    .Y(n_503));
 AND3x4_ASAP7_75t_SL g194248 (.A(n_136),
    .B(o8_we),
    .C(n_43530),
    .Y(n_43534));
 AND2x2_ASAP7_75t_SL g194249 (.A(n_503),
    .B(n_33100),
    .Y(n_43535));
 AND2x4_ASAP7_75t_L g194250 (.A(n_503),
    .B(n_33100),
    .Y(n_43536));
 AO21x1_ASAP7_75t_SL g194315 (.A1(n_49618),
    .A2(n_25398),
    .B(n_38761),
    .Y(n_43604));
 NAND2xp5_ASAP7_75t_SL g194374 (.A(n_36528),
    .B(n_35550),
    .Y(n_43665));
 AOI22xp33_ASAP7_75t_SL g194375 (.A1(\u8_mem[2] [31]),
    .A2(n_51488),
    .B1(\u8_mem[3] [31]),
    .B2(n_14001),
    .Y(n_43666));
 AOI22xp33_ASAP7_75t_SL g194376 (.A1(\u8_mem[0] [31]),
    .A2(n_27133),
    .B1(\u8_mem[1] [31]),
    .B2(n_27134),
    .Y(n_43667));
 OR2x2_ASAP7_75t_SL g194404 (.A(n_4448),
    .B(n_15100),
    .Y(n_43720));
 AOI22xp5_ASAP7_75t_SL g194437 (.A1(n_79104),
    .A2(n_43760),
    .B1(n_7430),
    .B2(n_38366),
    .Y(n_43761));
 NAND4xp25_ASAP7_75t_SL g194438 (.A(n_2185),
    .B(n_2193),
    .C(n_64794),
    .D(n_1461),
    .Y(n_43760));
 NAND2xp5_ASAP7_75t_SL g195 (.A(n_50290),
    .B(n_49131),
    .Y(n_14961));
 AOI22xp5_ASAP7_75t_SL g195056 (.A1(\u6_mem[3] [11]),
    .A2(n_77233),
    .B1(n_66843),
    .B2(n_61228),
    .Y(n_44440));
 AOI22xp5_ASAP7_75t_SL g195063 (.A1(\u6_mem[3] [8]),
    .A2(n_77233),
    .B1(n_65980),
    .B2(n_61228),
    .Y(n_44447));
 AOI22xp5_ASAP7_75t_SL g195068 (.A1(\u6_mem[3] [5]),
    .A2(n_77233),
    .B1(n_66869),
    .B2(n_61228),
    .Y(n_44452));
 AOI22xp5_ASAP7_75t_SL g195072 (.A1(\u6_mem[3] [0]),
    .A2(n_77233),
    .B1(n_75733),
    .B2(n_61228),
    .Y(n_44456));
 AOI22xp5_ASAP7_75t_SL g195169 (.A1(\u10_mem[1] [6]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_65879),
    .Y(n_44556));
 AOI22xp5_ASAP7_75t_SL g195458 (.A1(\u6_mem[3] [9]),
    .A2(n_77233),
    .B1(n_79971),
    .B2(n_61228),
    .Y(n_44864));
 INVx8_ASAP7_75t_SL g195911 (.A(n_24739),
    .Y(n_45330));
 AOI22xp5_ASAP7_75t_SL g195965 (.A1(\u6_mem[3] [3]),
    .A2(n_77233),
    .B1(n_66856),
    .B2(n_61228),
    .Y(n_45388));
 AOI22xp5_ASAP7_75t_SL g196136 (.A1(\u11_mem[2] [25]),
    .A2(n_61785),
    .B1(n_4909),
    .B2(n_45625),
    .Y(n_45569));
 AOI22xp5_ASAP7_75t_SL g196171 (.A1(\u11_mem[2] [31]),
    .A2(n_61785),
    .B1(n_30483),
    .B2(n_45625),
    .Y(n_45607));
 OAI22xp5_ASAP7_75t_SL g196187 (.A1(n_1701),
    .A2(n_1679),
    .B1(n_34484),
    .B2(n_10937),
    .Y(n_45624));
 INVx5_ASAP7_75t_SL g196188 (.A(n_23287),
    .Y(n_45625));
 OAI22xp33_ASAP7_75t_SL g196605 (.A1(n_432),
    .A2(n_11011),
    .B1(n_185),
    .B2(n_10576),
    .Y(n_46110));
 AOI22xp5_ASAP7_75t_SL g196639 (.A1(crac_out[18]),
    .A2(n_56881),
    .B1(n_10171),
    .B2(n_12219),
    .Y(n_46163));
 OA21x2_ASAP7_75t_SL g196651 (.A1(n_70322),
    .A2(n_3468),
    .B(n_198),
    .Y(n_46182));
 INVx1_ASAP7_75t_SL g196652 (.A(n_46182),
    .Y(n_46183));
 AND2x2_ASAP7_75t_R g196653 (.A(n_46184),
    .B(out_slt7[19]),
    .Y(n_46185));
 BUFx3_ASAP7_75t_SL g196654 (.A(n_46182),
    .Y(n_46184));
 NAND2xp5_ASAP7_75t_SL g196655 (.A(n_46186),
    .B(out_slt7[18]),
    .Y(n_46187));
 INVxp67_ASAP7_75t_SL g196656 (.A(n_46183),
    .Y(n_46186));
 NAND2xp5_ASAP7_75t_L g196658 (.A(n_46184),
    .B(out_slt7[8]),
    .Y(n_46189));
 NAND2xp5_ASAP7_75t_L g196659 (.A(out_slt7[9]),
    .B(n_46184),
    .Y(n_46190));
 AOI22xp33_ASAP7_75t_SL g196660 (.A1(n_4527),
    .A2(n_27129),
    .B1(n_46184),
    .B2(out_slt7[1]),
    .Y(n_46191));
 INVxp67_ASAP7_75t_SL g196661 (.A(n_263),
    .Y(n_46192));
 BUFx3_ASAP7_75t_SL g196662 (.A(n_263),
    .Y(n_1679));
 INVx2_ASAP7_75t_SL g196696 (.A(n_47551),
    .Y(n_46227));
 AND2x2_ASAP7_75t_SL g196697 (.A(n_7418),
    .B(n_33786),
    .Y(n_46228));
 NOR2xp33_ASAP7_75t_SL g196698 (.A(n_24511),
    .B(n_1781),
    .Y(n_46229));
 AND2x2_ASAP7_75t_SL g196700 (.A(u11_rp[0]),
    .B(u11_rp[1]),
    .Y(n_46232));
 NAND2xp5_ASAP7_75t_SL g196701 (.A(n_46234),
    .B(i6_re),
    .Y(n_46235));
 AOI22xp33_ASAP7_75t_SL g196703 (.A1(n_1167),
    .A2(\u11_mem[1] [15]),
    .B1(n_46234),
    .B2(\u11_mem[3] [15]),
    .Y(n_46236));
 AOI22xp33_ASAP7_75t_SL g196704 (.A1(n_1167),
    .A2(\u11_mem[1] [9]),
    .B1(n_46234),
    .B2(\u11_mem[3] [9]),
    .Y(n_46237));
 AOI22xp33_ASAP7_75t_SL g196705 (.A1(n_1167),
    .A2(\u11_mem[1] [24]),
    .B1(n_46234),
    .B2(\u11_mem[3] [24]),
    .Y(n_46238));
 AOI22xp33_ASAP7_75t_SL g196706 (.A1(n_1167),
    .A2(\u11_mem[1] [2]),
    .B1(n_46234),
    .B2(\u11_mem[3] [2]),
    .Y(n_46239));
 AOI22xp33_ASAP7_75t_SL g196707 (.A1(n_1167),
    .A2(\u11_mem[1] [10]),
    .B1(n_46234),
    .B2(\u11_mem[3] [10]),
    .Y(n_46240));
 AOI22xp33_ASAP7_75t_SL g196708 (.A1(n_1167),
    .A2(\u11_mem[1] [3]),
    .B1(n_46234),
    .B2(\u11_mem[3] [3]),
    .Y(n_46241));
 AOI22xp33_ASAP7_75t_SL g196709 (.A1(n_1167),
    .A2(\u11_mem[1] [12]),
    .B1(n_46234),
    .B2(\u11_mem[3] [12]),
    .Y(n_46242));
 AOI22xp33_ASAP7_75t_SL g196710 (.A1(n_1167),
    .A2(\u11_mem[1] [8]),
    .B1(n_46234),
    .B2(\u11_mem[3] [8]),
    .Y(n_46243));
 AOI22xp33_ASAP7_75t_SL g196711 (.A1(n_1167),
    .A2(\u11_mem[1] [20]),
    .B1(n_46234),
    .B2(\u11_mem[3] [20]),
    .Y(n_46244));
 AOI22xp33_ASAP7_75t_SL g196712 (.A1(n_1167),
    .A2(\u11_mem[1] [4]),
    .B1(n_46234),
    .B2(\u11_mem[3] [4]),
    .Y(n_46245));
 AOI22xp33_ASAP7_75t_SL g196713 (.A1(n_1167),
    .A2(\u11_mem[1] [0]),
    .B1(n_46234),
    .B2(\u11_mem[3] [0]),
    .Y(n_46246));
 AOI22xp33_ASAP7_75t_SL g196714 (.A1(n_1167),
    .A2(\u11_mem[1] [22]),
    .B1(n_46234),
    .B2(\u11_mem[3] [22]),
    .Y(n_46247));
 AOI22xp33_ASAP7_75t_SL g196715 (.A1(n_1167),
    .A2(\u11_mem[1] [23]),
    .B1(n_46234),
    .B2(\u11_mem[3] [23]),
    .Y(n_46248));
 AOI22xp33_ASAP7_75t_SL g196716 (.A1(n_1167),
    .A2(\u11_mem[1] [25]),
    .B1(n_46234),
    .B2(\u11_mem[3] [25]),
    .Y(n_46249));
 AOI22xp33_ASAP7_75t_SL g196717 (.A1(n_1167),
    .A2(\u11_mem[1] [6]),
    .B1(n_46234),
    .B2(\u11_mem[3] [6]),
    .Y(n_46250));
 AOI22xp33_ASAP7_75t_SL g196718 (.A1(n_1167),
    .A2(\u11_mem[1] [14]),
    .B1(n_46234),
    .B2(\u11_mem[3] [14]),
    .Y(n_46251));
 AOI22xp33_ASAP7_75t_SL g196719 (.A1(n_1167),
    .A2(\u11_mem[1] [19]),
    .B1(n_46234),
    .B2(\u11_mem[3] [19]),
    .Y(n_46252));
 AOI22xp33_ASAP7_75t_SL g196720 (.A1(n_1167),
    .A2(\u11_mem[1] [1]),
    .B1(n_46234),
    .B2(\u11_mem[3] [1]),
    .Y(n_46253));
 AOI22xp33_ASAP7_75t_SL g196721 (.A1(n_1167),
    .A2(\u11_mem[1] [17]),
    .B1(n_46234),
    .B2(\u11_mem[3] [17]),
    .Y(n_46254));
 AOI22xp33_ASAP7_75t_SL g196722 (.A1(n_1167),
    .A2(\u11_mem[1] [5]),
    .B1(n_46234),
    .B2(\u11_mem[3] [5]),
    .Y(n_46255));
 AOI22xp33_ASAP7_75t_SL g196723 (.A1(n_1167),
    .A2(\u11_mem[1] [29]),
    .B1(n_46234),
    .B2(\u11_mem[3] [29]),
    .Y(n_46256));
 AOI22xp33_ASAP7_75t_SL g196724 (.A1(n_1167),
    .A2(\u11_mem[1] [27]),
    .B1(n_46234),
    .B2(\u11_mem[3] [27]),
    .Y(n_46257));
 AOI22xp33_ASAP7_75t_SL g196725 (.A1(n_1167),
    .A2(\u11_mem[1] [30]),
    .B1(n_46234),
    .B2(\u11_mem[3] [30]),
    .Y(n_46258));
 AOI22xp33_ASAP7_75t_SL g196726 (.A1(n_1167),
    .A2(\u11_mem[1] [18]),
    .B1(n_46234),
    .B2(\u11_mem[3] [18]),
    .Y(n_46259));
 AOI22xp33_ASAP7_75t_SL g196727 (.A1(n_1167),
    .A2(\u11_mem[1] [11]),
    .B1(n_46234),
    .B2(\u11_mem[3] [11]),
    .Y(n_46260));
 AOI22xp33_ASAP7_75t_SL g196728 (.A1(n_1167),
    .A2(\u11_mem[1] [31]),
    .B1(n_46234),
    .B2(\u11_mem[3] [31]),
    .Y(n_46261));
 AOI22xp33_ASAP7_75t_SL g196729 (.A1(n_1167),
    .A2(\u11_mem[1] [21]),
    .B1(n_46234),
    .B2(\u11_mem[3] [21]),
    .Y(n_46262));
 AOI22xp33_ASAP7_75t_SL g196730 (.A1(n_1167),
    .A2(\u11_mem[1] [7]),
    .B1(n_46234),
    .B2(\u11_mem[3] [7]),
    .Y(n_46263));
 AOI22xp5_ASAP7_75t_SL g196753 (.A1(\u8_mem[1] [17]),
    .A2(n_73399),
    .B1(n_10143),
    .B2(n_73997),
    .Y(n_46289));
 NAND2x1_ASAP7_75t_SL g196789 (.A(n_33787),
    .B(n_41606),
    .Y(n_46334));
 NAND4xp25_ASAP7_75t_SL g196790 (.A(n_15084),
    .B(n_46335),
    .C(n_15085),
    .D(n_15087),
    .Y(n_46336));
 NAND2xp5_ASAP7_75t_SL g196791 (.A(n_46334),
    .B(n_47551),
    .Y(n_46335));
 AOI22xp5_ASAP7_75t_SL g196865 (.A1(\u6_mem[3] [15]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_28913),
    .Y(n_46422));
 AOI22xp5_ASAP7_75t_SL g196914 (.A1(n_46477),
    .A2(\u10_mem[0] [10]),
    .B1(n_46478),
    .B2(n_46479),
    .Y(n_46480));
 INVx6_ASAP7_75t_SL g196915 (.A(n_26250),
    .Y(n_46477));
 AND2x6_ASAP7_75t_SL g196916 (.A(n_31801),
    .B(n_33604),
    .Y(n_46478));
 NAND2xp5_ASAP7_75t_SL g196917 (.A(n_18524),
    .B(n_1228),
    .Y(n_46479));
 AOI22xp5_ASAP7_75t_SL g196922 (.A1(\u4_mem[1] [26]),
    .A2(n_1765),
    .B1(\u4_mem[0] [26]),
    .B2(n_1766),
    .Y(n_46485));
 NAND2xp5_ASAP7_75t_SL g196982 (.A(n_48630),
    .B(n_50461),
    .Y(n_46558));
 AOI22xp5_ASAP7_75t_SL g196984 (.A1(n_24735),
    .A2(n_46562),
    .B1(\u9_mem[3] [3]),
    .B2(n_45330),
    .Y(n_46563));
 NAND2xp5_ASAP7_75t_SL g196985 (.A(n_48629),
    .B(n_50460),
    .Y(n_46562));
 NAND2xp5_ASAP7_75t_SL g196989 (.A(n_46564),
    .B(n_56059),
    .Y(n_46566));
 NOR2xp67_ASAP7_75t_SL g196990 (.A(n_37384),
    .B(n_24516),
    .Y(n_46564));
 AOI22xp33_ASAP7_75t_SL g197007 (.A1(\u9_mem[0] [0]),
    .A2(n_46587),
    .B1(n_31720),
    .B2(n_40712),
    .Y(n_46588));
 INVx8_ASAP7_75t_SL g197008 (.A(n_17925),
    .Y(n_46587));
 AOI21xp5_ASAP7_75t_SL g197057 (.A1(n_46639),
    .A2(n_46638),
    .B(oc1_int_set[1]),
    .Y(n_46640));
 AND2x2_ASAP7_75t_R g197058 (.A(n_43),
    .B(n_4040),
    .Y(n_46638));
 INVxp67_ASAP7_75t_SL g197059 (.A(n_36089),
    .Y(n_46639));
 NAND2xp5_ASAP7_75t_SL g197061 (.A(n_78955),
    .B(n_47357),
    .Y(n_46642));
 NAND4xp25_ASAP7_75t_SL g197062 (.A(n_37350),
    .B(n_46643),
    .C(n_27219),
    .D(n_23079),
    .Y(n_46644));
 NAND2xp5_ASAP7_75t_SL g197063 (.A(n_46642),
    .B(n_78041),
    .Y(n_46643));
 A2O1A1Ixp33_ASAP7_75t_SL g197105 (.A1(n_46697),
    .A2(n_46698),
    .B(n_64852),
    .C(n_46700),
    .Y(n_46701));
 INVx2_ASAP7_75t_SL g197106 (.A(n_7990),
    .Y(n_46697));
 NAND2xp5_ASAP7_75t_SL g197107 (.A(n_1932),
    .B(n_26733),
    .Y(n_46698));
 NAND2xp5_ASAP7_75t_L g197109 (.A(out_slt4[9]),
    .B(n_4253),
    .Y(n_46700));
 AOI22xp5_ASAP7_75t_SL g197155 (.A1(\u10_mem[1] [9]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_18707),
    .Y(n_46750));
 AOI22xp5_ASAP7_75t_SL g197482 (.A1(n_10660),
    .A2(n_64818),
    .B1(\u8_mem[3] [30]),
    .B2(n_72908),
    .Y(n_47121));
 AOI22xp5_ASAP7_75t_SL g197487 (.A1(n_28316),
    .A2(n_64861),
    .B1(\u6_mem[3] [25]),
    .B2(n_72084),
    .Y(n_47127));
 AOI22xp5_ASAP7_75t_SL g197522 (.A1(n_28424),
    .A2(n_64861),
    .B1(\u6_mem[3] [24]),
    .B2(n_72084),
    .Y(n_47164));
 AOI22xp5_ASAP7_75t_SL g197539 (.A1(n_65927),
    .A2(n_64819),
    .B1(\u8_mem[3] [25]),
    .B2(n_11204),
    .Y(n_47184));
 AOI22xp5_ASAP7_75t_SL g197544 (.A1(n_65908),
    .A2(n_64818),
    .B1(\u8_mem[3] [27]),
    .B2(n_11204),
    .Y(n_47192));
 AOI22xp5_ASAP7_75t_SL g197567 (.A1(n_65900),
    .A2(n_64818),
    .B1(\u8_mem[3] [31]),
    .B2(n_72908),
    .Y(n_47217));
 AOI22xp5_ASAP7_75t_SL g197605 (.A1(n_32644),
    .A2(n_47390),
    .B1(\u4_mem[3] [6]),
    .B2(n_35908),
    .Y(n_47255));
 AOI22xp5_ASAP7_75t_SL g197608 (.A1(n_73996),
    .A2(n_64818),
    .B1(\u8_mem[3] [21]),
    .B2(n_11204),
    .Y(n_47261));
 AOI22xp5_ASAP7_75t_SL g197613 (.A1(n_10684),
    .A2(n_64819),
    .B1(\u8_mem[3] [29]),
    .B2(n_72908),
    .Y(n_47266));
 AOI22xp5_ASAP7_75t_SL g197631 (.A1(n_66010),
    .A2(n_64818),
    .B1(\u8_mem[3] [26]),
    .B2(n_11204),
    .Y(n_47287));
 AOI22xp5_ASAP7_75t_SL g197647 (.A1(\u6_mem[2] [10]),
    .A2(n_77853),
    .B1(\u6_mem[3] [10]),
    .B2(n_41152),
    .Y(n_47306));
 AOI22xp5_ASAP7_75t_SL g197661 (.A1(n_66868),
    .A2(n_47390),
    .B1(\u4_mem[3] [5]),
    .B2(n_35908),
    .Y(n_47322));
 AOI22xp5_ASAP7_75t_SL g197673 (.A1(n_33024),
    .A2(n_47390),
    .B1(\u4_mem[3] [20]),
    .B2(n_35909),
    .Y(n_47334));
 AOI22xp5_ASAP7_75t_SL g197679 (.A1(n_28381),
    .A2(n_64819),
    .B1(\u8_mem[3] [23]),
    .B2(n_72908),
    .Y(n_47340));
 AOI22xp5_ASAP7_75t_SL g197686 (.A1(n_65941),
    .A2(n_64818),
    .B1(\u8_mem[3] [22]),
    .B2(n_11204),
    .Y(n_47348));
 AOI22xp5_ASAP7_75t_SL g197695 (.A1(\u6_mem[2] [14]),
    .A2(n_77853),
    .B1(\u6_mem[3] [14]),
    .B2(n_41152),
    .Y(n_47357));
 AOI22xp5_ASAP7_75t_SL g197708 (.A1(n_65917),
    .A2(n_64818),
    .B1(\u8_mem[3] [24]),
    .B2(n_11204),
    .Y(n_47373));
 AOI22xp5_ASAP7_75t_SL g197726 (.A1(n_65969),
    .A2(n_47390),
    .B1(\u4_mem[3] [7]),
    .B2(n_35908),
    .Y(n_47391));
 INVx6_ASAP7_75t_SL g197727 (.A(n_35911),
    .Y(n_47390));
 AOI22xp5_ASAP7_75t_SL g197738 (.A1(n_10638),
    .A2(n_73997),
    .B1(\u8_mem[1] [30]),
    .B2(n_75735),
    .Y(n_47403));
 AOI22xp5_ASAP7_75t_SL g197748 (.A1(n_10247),
    .A2(n_64819),
    .B1(\u8_mem[3] [20]),
    .B2(n_11204),
    .Y(n_47415));
 OAI21xp5_ASAP7_75t_SL g197826 (.A1(n_50808),
    .A2(n_47498),
    .B(n_17687),
    .Y(n_47500));
 AOI21xp33_ASAP7_75t_SL g197827 (.A1(n_21092),
    .A2(i4_re),
    .B(n_28774),
    .Y(n_47498));
 AOI21xp33_ASAP7_75t_R g197863 (.A1(n_19013),
    .A2(n_47538),
    .B(n_24725),
    .Y(n_47539));
 AND2x2_ASAP7_75t_SL g197864 (.A(u26_ps_cnt[1]),
    .B(u26_ps_cnt[0]),
    .Y(n_47538));
 NAND3xp33_ASAP7_75t_SL g197865 (.A(n_47538),
    .B(n_19013),
    .C(n_24726),
    .Y(n_47540));
 INVx1_ASAP7_75t_SL g197866 (.A(n_47538),
    .Y(n_47541));
 AND2x4_ASAP7_75t_SL g197875 (.A(n_417),
    .B(n_176),
    .Y(n_47551));
 NAND2x1_ASAP7_75t_SL g197876 (.A(n_41034),
    .B(n_13557),
    .Y(n_47552));
 NAND4xp25_ASAP7_75t_SL g197877 (.A(n_2176),
    .B(n_1780),
    .C(n_1747),
    .D(n_47553),
    .Y(n_47554));
 NAND2xp5_ASAP7_75t_SL g197878 (.A(n_47552),
    .B(n_47551),
    .Y(n_47553));
 NAND2xp5_ASAP7_75t_SL g197927 (.A(n_48628),
    .B(n_48627),
    .Y(n_47616));
 INVx1_ASAP7_75t_R g197929 (.A(n_399),
    .Y(n_47613));
 NAND2xp5_ASAP7_75t_SL g197943 (.A(n_12070),
    .B(n_78957),
    .Y(n_47631));
 INVxp67_ASAP7_75t_L g197944 (.A(n_47631),
    .Y(n_47632));
 NAND4xp25_ASAP7_75t_SL g197985 (.A(n_31871),
    .B(n_41323),
    .C(n_14859),
    .D(n_1455),
    .Y(n_47682));
 INVxp33_ASAP7_75t_SL g198008 (.A(n_31895),
    .Y(n_47706));
 INVxp33_ASAP7_75t_L g198009 (.A(n_65643),
    .Y(n_47707));
 INVxp33_ASAP7_75t_L g198038 (.A(oc5_cfg[0]),
    .Y(n_47739));
 BUFx3_ASAP7_75t_SL g198039 (.A(oc5_cfg[0]),
    .Y(n_47740));
 NAND2xp5_ASAP7_75t_SL g198064 (.A(n_25438),
    .B(u10_wp[2]),
    .Y(n_47767));
 INVx3_ASAP7_75t_SL g198065 (.A(n_33604),
    .Y(n_47768));
 AOI21xp5_ASAP7_75t_SL g198066 (.A1(n_36975),
    .A2(n_4667),
    .B(n_47771),
    .Y(n_47772));
 NAND2xp5_ASAP7_75t_L g198067 (.A(n_47769),
    .B(n_47770),
    .Y(n_47771));
 NAND2xp33_ASAP7_75t_R g198068 (.A(n_47767),
    .B(\u10_mem[2] [24]),
    .Y(n_47769));
 NAND2xp33_ASAP7_75t_L g198069 (.A(n_47768),
    .B(\u10_mem[2] [24]),
    .Y(n_47770));
 NOR2xp33_ASAP7_75t_SL g198075 (.A(n_27061),
    .B(n_10576),
    .Y(n_47778));
 NAND2xp5_ASAP7_75t_SL g198076 (.A(u6_wp[0]),
    .B(o7_we),
    .Y(n_47780));
 AND3x4_ASAP7_75t_SL g198082 (.A(n_20669),
    .B(o7_we),
    .C(n_24745),
    .Y(n_47786));
 NAND2xp67_ASAP7_75t_SL g198083 (.A(o7_we),
    .B(n_24745),
    .Y(n_47787));
 AOI221xp5_ASAP7_75t_SL g198086 (.A1(n_7082),
    .A2(u13_intm_r[14]),
    .B1(i4_dout[14]),
    .B2(n_8173),
    .C(n_14908),
    .Y(n_47793));
 AOI22xp5_ASAP7_75t_SL g198087 (.A1(n_66032),
    .A2(n_6732),
    .B1(n_47791),
    .B2(n_32335),
    .Y(n_47792));
 HB1xp67_ASAP7_75t_R g198088 (.A(u13_intm_r[14]),
    .Y(n_47791));
 AOI22xp5_ASAP7_75t_SL g198089 (.A1(u13_intm_r[15]),
    .A2(u13_ints_r[15]),
    .B1(u13_intm_r[14]),
    .B2(u13_ints_r[14]),
    .Y(n_47794));
 OAI221xp5_ASAP7_75t_SL g198251 (.A1(n_48057),
    .A2(n_48052),
    .B1(n_50452),
    .B2(n_48053),
    .C(n_48626),
    .Y(n_48055));
 INVx1_ASAP7_75t_SL g198253 (.A(in_slt3[14]),
    .Y(n_48052));
 INVx1_ASAP7_75t_SL g198254 (.A(in_slt3[12]),
    .Y(n_48053));
 OAI22xp5_ASAP7_75t_SL g198256 (.A1(n_48056),
    .A2(n_48057),
    .B1(n_48058),
    .B2(n_50452),
    .Y(n_48060));
 BUFx6f_ASAP7_75t_SL g198257 (.A(n_329),
    .Y(n_48057));
 INVx1_ASAP7_75t_L g198258 (.A(in_slt3[4]),
    .Y(n_48058));
 INVx2_ASAP7_75t_SL g198302 (.A(n_35902),
    .Y(n_48105));
 INVx2_ASAP7_75t_L g198304 (.A(n_48105),
    .Y(n_48106));
 AND2x4_ASAP7_75t_SL g198305 (.A(n_48106),
    .B(n_37935),
    .Y(n_48109));
 INVx1_ASAP7_75t_SL g198308 (.A(n_48106),
    .Y(n_48110));
 NOR2x2_ASAP7_75t_SL g198342 (.A(n_47768),
    .B(n_47767),
    .Y(n_48145));
 AOI22xp5_ASAP7_75t_SL g198369 (.A1(n_65879),
    .A2(n_36975),
    .B1(n_48153),
    .B2(\u10_mem[2] [6]),
    .Y(n_48174));
 AOI22xp5_ASAP7_75t_SL g198372 (.A1(n_36975),
    .A2(n_40956),
    .B1(\u10_mem[2] [0]),
    .B2(n_48153),
    .Y(n_48177));
 INVx4_ASAP7_75t_SL g198416 (.A(n_34235),
    .Y(n_48223));
 AOI211x1_ASAP7_75t_SL g198417 (.A1(n_2350),
    .A2(n_25954),
    .B(n_48224),
    .C(n_46185),
    .Y(n_48225));
 AOI22xp5_ASAP7_75t_SL g198570 (.A1(\u6_mem[1] [18]),
    .A2(n_76763),
    .B1(\u6_mem[3] [18]),
    .B2(n_41152),
    .Y(n_48404));
 AOI22xp5_ASAP7_75t_SL g198572 (.A1(\u6_mem[1] [12]),
    .A2(n_76763),
    .B1(\u6_mem[3] [12]),
    .B2(n_41152),
    .Y(n_48405));
 AOI22xp5_ASAP7_75t_SL g198574 (.A1(\u6_mem[3] [6]),
    .A2(n_41152),
    .B1(n_76763),
    .B2(\u6_mem[1] [6]),
    .Y(n_48407));
 AOI22xp33_ASAP7_75t_SL g198579 (.A1(n_76763),
    .A2(\u6_mem[1] [5]),
    .B1(n_41152),
    .B2(\u6_mem[3] [5]),
    .Y(n_48412));
 AOI22xp5_ASAP7_75t_SL g198580 (.A1(\u6_mem[3] [7]),
    .A2(n_41152),
    .B1(n_76763),
    .B2(\u6_mem[1] [7]),
    .Y(n_48413));
 AND2x4_ASAP7_75t_SL g198582 (.A(n_37337),
    .B(n_76763),
    .Y(n_48415));
 AOI22xp5_ASAP7_75t_SL g198590 (.A1(n_76763),
    .A2(\u6_mem[1] [19]),
    .B1(\u6_mem[3] [19]),
    .B2(n_41152),
    .Y(n_48423));
 HB1xp67_ASAP7_75t_L g198593 (.A(n_76763),
    .Y(n_48425));
 INVx2_ASAP7_75t_SL g198594 (.A(n_48427),
    .Y(n_48428));
 INVx1_ASAP7_75t_SL g198595 (.A(u3_wp[1]),
    .Y(n_48427));
 OAI31xp33_ASAP7_75t_SL g198596 (.A1(n_21543),
    .A2(n_48429),
    .A3(n_65952),
    .B(n_48430),
    .Y(n_48431));
 INVx1_ASAP7_75t_L g198597 (.A(n_48428),
    .Y(n_48429));
 OAI21xp5_ASAP7_75t_SL g198598 (.A1(n_48429),
    .A2(n_21543),
    .B(n_21546),
    .Y(n_48430));
 OAI31xp33_ASAP7_75t_SL g198599 (.A1(n_21521),
    .A2(n_48429),
    .A3(n_32916),
    .B(n_48433),
    .Y(n_48434));
 OAI21xp5_ASAP7_75t_SL g198600 (.A1(n_48432),
    .A2(n_21521),
    .B(n_8),
    .Y(n_48433));
 INVx1_ASAP7_75t_SL g198601 (.A(u3_wp[1]),
    .Y(n_48432));
 AND3x4_ASAP7_75t_SL g198603 (.A(n_41910),
    .B(n_48432),
    .C(o3_we),
    .Y(n_48436));
 AO22x1_ASAP7_75t_SL g198604 (.A1(n_48432),
    .A2(n_24588),
    .B1(n_24587),
    .B2(n_48676),
    .Y(n_48437));
 NAND2x1_ASAP7_75t_SL g198621 (.A(n_48454),
    .B(n_48455),
    .Y(n_48456));
 AOI22xp5_ASAP7_75t_SL g198622 (.A1(u10_din_tmp1[1]),
    .A2(n_24336),
    .B1(in_slt4[3]),
    .B2(n_1666),
    .Y(n_48454));
 NAND2xp5_ASAP7_75t_SL g198623 (.A(in_slt4[1]),
    .B(n_1667),
    .Y(n_48455));
 NAND2xp5_ASAP7_75t_SL g198735 (.A(u9_din_tmp1[12]),
    .B(n_48625),
    .Y(n_48626));
 NOR2x1_ASAP7_75t_SL g198737 (.A(n_427),
    .B(n_286),
    .Y(n_48624));
 AO21x1_ASAP7_75t_SL g198738 (.A1(n_48625),
    .A2(n_17402),
    .B(n_47613),
    .Y(n_48627));
 NAND3xp33_ASAP7_75t_L g198739 (.A(n_48625),
    .B(n_17402),
    .C(n_47613),
    .Y(n_48628));
 AOI22xp33_ASAP7_75t_SL g198740 (.A1(in_slt3[5]),
    .A2(n_1692),
    .B1(u9_din_tmp1[3]),
    .B2(n_48625),
    .Y(n_48629));
 AOI22xp33_ASAP7_75t_SL g198741 (.A1(in_slt3[4]),
    .A2(n_1692),
    .B1(u9_din_tmp1[2]),
    .B2(n_48625),
    .Y(n_48630));
 AOI22xp5_ASAP7_75t_SL g198742 (.A1(u9_din_tmp1[0]),
    .A2(n_48625),
    .B1(in_slt3[2]),
    .B2(n_1692),
    .Y(n_48631));
 NAND4xp25_ASAP7_75t_SL g198743 (.A(n_48625),
    .B(n_24738),
    .C(n_50426),
    .D(n_21600),
    .Y(n_48632));
 NAND2xp5_ASAP7_75t_L g198744 (.A(n_48633),
    .B(u9_din_tmp1[5]),
    .Y(n_48634));
 NAND2xp5_ASAP7_75t_SL g198746 (.A(n_48625),
    .B(u9_din_tmp1[10]),
    .Y(n_48635));
 NAND2xp5_ASAP7_75t_L g198747 (.A(u9_din_tmp1[9]),
    .B(n_48625),
    .Y(n_48636));
 NAND2xp5_ASAP7_75t_SL g198749 (.A(u9_din_tmp1[6]),
    .B(n_48625),
    .Y(n_48638));
 AOI22xp5_ASAP7_75t_SL g198750 (.A1(u9_din_tmp1[1]),
    .A2(n_48625),
    .B1(in_slt3[3]),
    .B2(n_1692),
    .Y(n_48639));
 NAND2xp5_ASAP7_75t_L g198751 (.A(u9_din_tmp1[8]),
    .B(n_48625),
    .Y(n_48640));
 AO21x1_ASAP7_75t_L g198753 (.A1(u9_din_tmp1[4]),
    .A2(n_48633),
    .B(n_48060),
    .Y(n_48642));
 NAND2xp33_ASAP7_75t_SL g198754 (.A(u9_din_tmp1[11]),
    .B(n_48633),
    .Y(n_48643));
 NAND2xp5_ASAP7_75t_L g198755 (.A(u9_din_tmp1[15]),
    .B(n_48633),
    .Y(n_48644));
 NAND2xp5_ASAP7_75t_SL g198756 (.A(n_48633),
    .B(u9_din_tmp1[7]),
    .Y(n_48645));
 NAND2xp5_ASAP7_75t_L g198757 (.A(u9_din_tmp1[14]),
    .B(n_48633),
    .Y(n_48646));
 NAND2xp5_ASAP7_75t_L g198758 (.A(u9_din_tmp1[13]),
    .B(n_48633),
    .Y(n_48647));
 BUFx3_ASAP7_75t_SL g198781 (.A(n_190),
    .Y(n_48675));
 INVxp33_ASAP7_75t_L g198782 (.A(n_190),
    .Y(n_48676));
 NAND2x1_ASAP7_75t_SL g198833 (.A(n_27038),
    .B(n_50389),
    .Y(n_48729));
 INVxp33_ASAP7_75t_SL g199 (.A(n_49131),
    .Y(n_14963));
 AND2x6_ASAP7_75t_SL g199173 (.A(n_7653),
    .B(n_51030),
    .Y(n_49129));
 NAND2xp5_ASAP7_75t_SL g199174 (.A(n_51034),
    .B(n_19502),
    .Y(n_49131));
 AOI31xp33_ASAP7_75t_SL g199186 (.A1(n_48437),
    .A2(n_40419),
    .A3(n_2688),
    .B(oc0_int_set[2]),
    .Y(n_49143));
 NOR3xp33_ASAP7_75t_SL g199211 (.A(n_49172),
    .B(n_49173),
    .C(n_50794),
    .Y(n_49175));
 OAI21xp5_ASAP7_75t_SL g199212 (.A1(n_68),
    .A2(n_10613),
    .B(n_7132),
    .Y(n_49172));
 OAI21xp5_ASAP7_75t_SL g199213 (.A1(n_65897),
    .A2(n_8340),
    .B(n_7174),
    .Y(n_49173));
 AND2x2_ASAP7_75t_SL g199216 (.A(n_78958),
    .B(n_49177),
    .Y(n_49178));
 AOI22xp33_ASAP7_75t_SL g199218 (.A1(n_77853),
    .A2(\u6_mem[2] [16]),
    .B1(n_41152),
    .B2(\u6_mem[3] [16]),
    .Y(n_49177));
 OAI211xp5_ASAP7_75t_SL g199219 (.A1(n_6122),
    .A2(n_49178),
    .B(n_1422),
    .C(n_7569),
    .Y(n_49180));
 A2O1A1Ixp33_ASAP7_75t_SL g199220 (.A1(n_49178),
    .A2(n_77964),
    .B(n_48223),
    .C(n_46187),
    .Y(n_49181));
 OAI221xp5_ASAP7_75t_SL g199221 (.A1(n_7442),
    .A2(n_13978),
    .B1(n_49178),
    .B2(n_37339),
    .C(n_36771),
    .Y(n_49182));
 NAND2xp5_ASAP7_75t_SL g199240 (.A(n_64834),
    .B(n_7883),
    .Y(n_49203));
 AND2x2_ASAP7_75t_L g199334 (.A(n_47740),
    .B(n_432),
    .Y(n_49309));
 OAI211xp5_ASAP7_75t_SL g199344 (.A1(n_8113),
    .A2(n_23671),
    .B(n_49319),
    .C(n_46698),
    .Y(n_49320));
 AOI22xp5_ASAP7_75t_SL g199410 (.A1(n_32650),
    .A2(n_75734),
    .B1(\u8_mem[1] [6]),
    .B2(n_31460),
    .Y(n_49387));
 OAI211xp5_ASAP7_75t_SL g199521 (.A1(n_46227),
    .A2(n_16672),
    .B(n_49499),
    .C(n_18841),
    .Y(n_49500));
 NAND2xp5_ASAP7_75t_SL g199522 (.A(n_425),
    .B(n_40287),
    .Y(n_49499));
 AND2x6_ASAP7_75t_SL g199621 (.A(u7_rp[1]),
    .B(n_7653),
    .Y(n_49617));
 AND2x6_ASAP7_75t_SL g199622 (.A(u7_rp[1]),
    .B(u7_rp[2]),
    .Y(n_49618));
 NAND2xp5_ASAP7_75t_SL g199623 (.A(n_51045),
    .B(n_49619),
    .Y(n_49620));
 AOI22xp5_ASAP7_75t_SL g199624 (.A1(n_49617),
    .A2(\u7_mem[1] [11]),
    .B1(\u7_mem[3] [11]),
    .B2(n_49618),
    .Y(n_49619));
 AOI22xp5_ASAP7_75t_SL g199637 (.A1(\u6_mem[3] [13]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_65955),
    .Y(n_49641));
 NOR3xp33_ASAP7_75t_SL g199705 (.A(n_50292),
    .B(n_4116),
    .C(n_247),
    .Y(n_49719));
 XNOR2xp5_ASAP7_75t_SL g2 (.A(u9_rp[2]),
    .B(n_13751),
    .Y(n_64133));
 NOR3x2_ASAP7_75t_SL g20 (.B(wb_addr_i[2]),
    .C(wb_addr_i[3]),
    .Y(n_22851),
    .A(n_8228));
 INVxp33_ASAP7_75t_R g200045 (.A(u26_ps_cnt[4]),
    .Y(n_50088));
 NAND2xp33_ASAP7_75t_L g200047 (.A(n_22837),
    .B(u26_ps_cnt[4]),
    .Y(n_50090));
 NAND3xp33_ASAP7_75t_SL g200049 (.A(u26_ps_cnt[5]),
    .B(u26_ps_cnt[4]),
    .C(u26_ps_cnt[0]),
    .Y(n_50091));
 AOI22xp5_ASAP7_75t_SL g200140 (.A1(n_3815),
    .A2(n_43537),
    .B1(\u7_mem[1] [1]),
    .B2(n_50218),
    .Y(n_50219));
 INVx4_ASAP7_75t_SL g200141 (.A(n_50217),
    .Y(n_50218));
 AND3x4_ASAP7_75t_SL g200142 (.A(u7_wp[0]),
    .B(o8_we),
    .C(n_33771),
    .Y(n_50217));
 AOI22xp5_ASAP7_75t_SL g200143 (.A1(n_50220),
    .A2(\u7_mem[1] [21]),
    .B1(n_73996),
    .B2(n_43536),
    .Y(n_50221));
 INVx5_ASAP7_75t_SL g200144 (.A(n_50217),
    .Y(n_50220));
 AOI22xp5_ASAP7_75t_SL g200145 (.A1(n_50218),
    .A2(\u7_mem[1] [29]),
    .B1(n_22715),
    .B2(n_43536),
    .Y(n_50222));
 AOI22xp5_ASAP7_75t_SL g200146 (.A1(n_50218),
    .A2(\u7_mem[1] [5]),
    .B1(n_10058),
    .B2(n_43537),
    .Y(n_50223));
 AOI22xp5_ASAP7_75t_SL g200147 (.A1(n_50218),
    .A2(\u7_mem[1] [27]),
    .B1(n_62940),
    .B2(n_43537),
    .Y(n_50224));
 AOI22xp5_ASAP7_75t_SL g200148 (.A1(n_33203),
    .A2(n_43535),
    .B1(\u7_mem[1] [0]),
    .B2(n_50218),
    .Y(n_50225));
 AOI22xp5_ASAP7_75t_SL g200149 (.A1(n_10640),
    .A2(n_43537),
    .B1(n_50218),
    .B2(\u7_mem[1] [30]),
    .Y(n_50226));
 AOI22xp5_ASAP7_75t_SL g200150 (.A1(n_28316),
    .A2(n_43537),
    .B1(n_50218),
    .B2(\u7_mem[1] [25]),
    .Y(n_50227));
 AOI22xp5_ASAP7_75t_SL g200151 (.A1(\u7_mem[1] [18]),
    .A2(n_50218),
    .B1(n_10194),
    .B2(n_43537),
    .Y(n_50228));
 AOI22xp5_ASAP7_75t_SL g200152 (.A1(n_50218),
    .A2(\u7_mem[1] [11]),
    .B1(n_66842),
    .B2(n_43537),
    .Y(n_50229));
 AOI22xp5_ASAP7_75t_SL g200153 (.A1(n_50218),
    .A2(\u7_mem[1] [9]),
    .B1(n_9942),
    .B2(n_43536),
    .Y(n_50230));
 AOI22xp5_ASAP7_75t_SL g200154 (.A1(n_50218),
    .A2(\u7_mem[1] [12]),
    .B1(n_10026),
    .B2(n_43537),
    .Y(n_50231));
 AOI22xp5_ASAP7_75t_SL g200155 (.A1(n_50218),
    .A2(\u7_mem[1] [19]),
    .B1(n_10196),
    .B2(n_43536),
    .Y(n_50232));
 AOI22xp5_ASAP7_75t_SL g200156 (.A1(n_50218),
    .A2(\u7_mem[1] [15]),
    .B1(n_28913),
    .B2(n_43536),
    .Y(n_50233));
 AOI22xp5_ASAP7_75t_SL g200157 (.A1(n_65969),
    .A2(n_43537),
    .B1(\u7_mem[1] [7]),
    .B2(n_50218),
    .Y(n_50234));
 AOI22xp33_ASAP7_75t_SL g200158 (.A1(n_50220),
    .A2(\u7_mem[1] [17]),
    .B1(n_65952),
    .B2(n_43536),
    .Y(n_50235));
 AOI22xp5_ASAP7_75t_SL g200159 (.A1(n_66004),
    .A2(n_43535),
    .B1(\u7_mem[1] [6]),
    .B2(n_50220),
    .Y(n_50236));
 AOI22xp5_ASAP7_75t_SL g200160 (.A1(n_50220),
    .A2(\u7_mem[1] [20]),
    .B1(n_66026),
    .B2(n_43535),
    .Y(n_50237));
 AOI22xp5_ASAP7_75t_SL g200161 (.A1(n_50220),
    .A2(\u7_mem[1] [23]),
    .B1(n_28381),
    .B2(n_43535),
    .Y(n_50238));
 AOI22xp5_ASAP7_75t_SL g200162 (.A1(\u7_mem[1] [2]),
    .A2(n_50220),
    .B1(n_28330),
    .B2(n_43535),
    .Y(n_50239));
 AOI22xp5_ASAP7_75t_SL g200163 (.A1(n_28251),
    .A2(n_43537),
    .B1(\u7_mem[1] [14]),
    .B2(n_50220),
    .Y(n_50240));
 AOI22xp5_ASAP7_75t_SL g200164 (.A1(n_28424),
    .A2(n_43537),
    .B1(\u7_mem[1] [24]),
    .B2(n_50220),
    .Y(n_50241));
 AOI22xp5_ASAP7_75t_SL g200165 (.A1(n_35041),
    .A2(n_43535),
    .B1(\u7_mem[1] [13]),
    .B2(n_50220),
    .Y(n_50242));
 AOI22xp5_ASAP7_75t_SL g200166 (.A1(n_35437),
    .A2(n_43536),
    .B1(\u7_mem[1] [26]),
    .B2(n_50220),
    .Y(n_50243));
 AOI22xp5_ASAP7_75t_SL g200168 (.A1(n_28276),
    .A2(n_43537),
    .B1(\u7_mem[1] [16]),
    .B2(n_50220),
    .Y(n_50245));
 AOI22xp5_ASAP7_75t_SL g200169 (.A1(n_28240),
    .A2(n_43537),
    .B1(\u7_mem[1] [8]),
    .B2(n_50220),
    .Y(n_50246));
 AOI22xp5_ASAP7_75t_SL g200170 (.A1(n_66855),
    .A2(n_43537),
    .B1(\u7_mem[1] [3]),
    .B2(n_50220),
    .Y(n_50247));
 AOI22xp5_ASAP7_75t_SL g200173 (.A1(n_50220),
    .A2(\u7_mem[1] [31]),
    .B1(n_15920),
    .B2(n_43536),
    .Y(n_50250));
 AOI22xp5_ASAP7_75t_SL g200174 (.A1(n_50220),
    .A2(\u7_mem[1] [28]),
    .B1(n_22640),
    .B2(n_43536),
    .Y(n_50251));
 INVx2_ASAP7_75t_SL g200191 (.A(oc4_cfg[3]),
    .Y(n_50287));
 OAI22xp5_ASAP7_75t_SL g200192 (.A1(n_11011),
    .A2(n_50287),
    .B1(n_14909),
    .B2(n_42),
    .Y(n_50289));
 AND2x2_ASAP7_75t_SL g200193 (.A(n_419),
    .B(n_50287),
    .Y(n_50290));
 AO21x1_ASAP7_75t_SL g200194 (.A1(n_51048),
    .A2(n_19503),
    .B(n_50287),
    .Y(n_50291));
 BUFx3_ASAP7_75t_SL g200195 (.A(n_50287),
    .Y(n_50292));
 INVx3_ASAP7_75t_SL g200196 (.A(n_50287),
    .Y(n_50293));
 OAI222xp33_ASAP7_75t_SL g200197 (.A1(n_2424),
    .A2(n_15100),
    .B1(n_16880),
    .B2(n_64715),
    .C1(n_4448),
    .C2(n_50292),
    .Y(n_50295));
 AND2x2_ASAP7_75t_L g200217 (.A(n_71350),
    .B(n_71351),
    .Y(n_50319));
 AND2x4_ASAP7_75t_SL g200239 (.A(n_40416),
    .B(n_6248),
    .Y(n_50341));
 NAND2x1_ASAP7_75t_SL g200241 (.A(n_50343),
    .B(n_33791),
    .Y(n_50344));
 AOI22xp5_ASAP7_75t_SL g200242 (.A1(\u3_mem[0] [10]),
    .A2(n_50341),
    .B1(n_50342),
    .B2(\u3_mem[2] [10]),
    .Y(n_50343));
 AOI22xp5_ASAP7_75t_SL g200276 (.A1(\u3_mem[2] [9]),
    .A2(n_50388),
    .B1(\u3_mem[3] [9]),
    .B2(n_71972),
    .Y(n_50389));
 NOR2xp33_ASAP7_75t_R g200312 (.A(n_399),
    .B(n_66054),
    .Y(n_50426));
 NAND3xp33_ASAP7_75t_SL g200315 (.A(n_21600),
    .B(n_24738),
    .C(n_66054),
    .Y(n_50427));
 BUFx3_ASAP7_75t_SL g200340 (.A(n_17584),
    .Y(n_50452));
 NAND2xp5_ASAP7_75t_SL g200341 (.A(in_slt3[0]),
    .B(n_50453),
    .Y(n_50454));
 INVx2_ASAP7_75t_SL g200342 (.A(n_50452),
    .Y(n_50453));
 NAND2xp5_ASAP7_75t_SL g200343 (.A(n_50455),
    .B(in_slt3[1]),
    .Y(n_50456));
 INVx1_ASAP7_75t_SL g200344 (.A(n_50452),
    .Y(n_50455));
 AOI22xp5_ASAP7_75t_SL g200345 (.A1(in_slt3[17]),
    .A2(n_50453),
    .B1(in_slt3[19]),
    .B2(n_1692),
    .Y(n_50457));
 INVx1_ASAP7_75t_SL g200346 (.A(n_50453),
    .Y(n_50458));
 AOI22xp5_ASAP7_75t_SL g200347 (.A1(in_slt3[16]),
    .A2(n_50453),
    .B1(in_slt3[18]),
    .B2(n_1692),
    .Y(n_50459));
 NAND2xp5_ASAP7_75t_SL g200348 (.A(in_slt3[3]),
    .B(n_50455),
    .Y(n_50460));
 NAND2xp5_ASAP7_75t_SL g200349 (.A(in_slt3[2]),
    .B(n_50455),
    .Y(n_50461));
 BUFx3_ASAP7_75t_SL g200411 (.A(n_17600),
    .Y(n_50546));
 INVx2_ASAP7_75t_SL g200412 (.A(n_50546),
    .Y(n_1667));
 OAI22xp5_ASAP7_75t_SL g200413 (.A1(n_14292),
    .A2(n_1534),
    .B1(n_50548),
    .B2(n_11693),
    .Y(n_50549));
 BUFx2_ASAP7_75t_SL g200414 (.A(n_50546),
    .Y(n_50548));
 OAI22xp5_ASAP7_75t_SL g200415 (.A1(n_64696),
    .A2(n_1534),
    .B1(n_50546),
    .B2(n_1699),
    .Y(n_50551));
 OAI211xp5_ASAP7_75t_SL g200417 (.A1(n_64696),
    .A2(n_50548),
    .B(n_1358),
    .C(n_42799),
    .Y(n_50552));
 OAI21xp5_ASAP7_75t_SL g200418 (.A1(n_26831),
    .A2(n_50548),
    .B(n_40379),
    .Y(n_50553));
 OAI211xp5_ASAP7_75t_L g200419 (.A1(n_64696),
    .A2(n_50548),
    .B(n_1358),
    .C(n_42799),
    .Y(n_50554));
 OAI21xp5_ASAP7_75t_SL g200420 (.A1(n_50548),
    .A2(n_26859),
    .B(n_40372),
    .Y(n_50555));
 OAI221xp5_ASAP7_75t_SL g200463 (.A1(n_5687),
    .A2(n_4496),
    .B1(n_5691),
    .B2(n_50601),
    .C(n_32583),
    .Y(n_50602));
 INVx1_ASAP7_75t_SL g200464 (.A(n_43088),
    .Y(n_50601));
 AOI22xp5_ASAP7_75t_SL g200520 (.A1(\u10_mem[1] [4]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_50555),
    .Y(n_50660));
 AOI221xp5_ASAP7_75t_SL g200558 (.A1(n_50706),
    .A2(n_5091),
    .B1(n_4988),
    .B2(out_slt9[11]),
    .C(n_4363),
    .Y(n_50707));
 NAND4xp25_ASAP7_75t_SL g200559 (.A(n_50702),
    .B(n_50703),
    .C(n_50704),
    .D(n_50705),
    .Y(n_50706));
 NAND2xp5_ASAP7_75t_L g200560 (.A(n_36528),
    .B(n_17618),
    .Y(n_50702));
 NAND2xp5_ASAP7_75t_SL g200561 (.A(n_16458),
    .B(n_2013),
    .Y(n_50703));
 AOI22xp33_ASAP7_75t_L g200562 (.A1(\u8_mem[2] [23]),
    .A2(n_51488),
    .B1(\u8_mem[3] [23]),
    .B2(n_14001),
    .Y(n_50704));
 AOI22xp33_ASAP7_75t_L g200563 (.A1(\u8_mem[0] [23]),
    .A2(n_27133),
    .B1(\u8_mem[1] [23]),
    .B2(n_27134),
    .Y(n_50705));
 AND2x6_ASAP7_75t_SL g200565 (.A(u4_rp[1]),
    .B(n_23524),
    .Y(n_50709));
 NOR2xp33_ASAP7_75t_SL g200566 (.A(n_50710),
    .B(n_1643),
    .Y(n_50711));
 AO22x1_ASAP7_75t_SL g200567 (.A1(n_58959),
    .A2(\u4_mem[0] [18]),
    .B1(\u4_mem[1] [18]),
    .B2(n_50709),
    .Y(n_50710));
 OAI21xp5_ASAP7_75t_SL g200568 (.A1(n_1643),
    .A2(n_50710),
    .B(n_35461),
    .Y(n_50712));
 NAND2xp5_ASAP7_75t_SL g200637 (.A(n_50792),
    .B(n_50793),
    .Y(n_50794));
 AOI22xp5_ASAP7_75t_SL g200638 (.A1(i4_dout[16]),
    .A2(n_8173),
    .B1(n_7082),
    .B2(u13_intm_r[16]),
    .Y(n_50792));
 NAND2xp5_ASAP7_75t_SL g200639 (.A(n_8212),
    .B(n_78094),
    .Y(n_50793));
 AND3x1_ASAP7_75t_SL g200646 (.A(i4_re),
    .B(n_28774),
    .C(n_21092),
    .Y(n_50808));
 NOR2xp33_ASAP7_75t_R g200650 (.A(n_29787),
    .B(n_50810),
    .Y(n_50812));
 NAND2xp5_ASAP7_75t_SL g200652 (.A(n_50810),
    .B(n_71392),
    .Y(n_50814));
 AOI22xp33_ASAP7_75t_SL g200830 (.A1(n_63785),
    .A2(\u7_mem[2] [6]),
    .B1(\u7_mem[3] [6]),
    .B2(n_49618),
    .Y(n_51032));
 AOI22xp5_ASAP7_75t_SL g200832 (.A1(n_63785),
    .A2(\u7_mem[2] [15]),
    .B1(\u7_mem[3] [15]),
    .B2(n_49618),
    .Y(n_51033));
 AOI22xp33_ASAP7_75t_SL g200833 (.A1(n_63785),
    .A2(\u7_mem[2] [2]),
    .B1(n_49129),
    .B2(\u7_mem[0] [2]),
    .Y(n_51034));
 HB1xp67_ASAP7_75t_SL g200835 (.A(n_63785),
    .Y(n_51035));
 AOI22xp5_ASAP7_75t_SL g200836 (.A1(n_49129),
    .A2(\u7_mem[0] [3]),
    .B1(\u7_mem[2] [3]),
    .B2(n_63785),
    .Y(n_51037));
 AOI22xp33_ASAP7_75t_SL g200837 (.A1(n_63785),
    .A2(\u7_mem[2] [7]),
    .B1(\u7_mem[3] [7]),
    .B2(n_49618),
    .Y(n_51038));
 AOI22xp5_ASAP7_75t_SL g200838 (.A1(n_63785),
    .A2(\u7_mem[2] [12]),
    .B1(\u7_mem[3] [12]),
    .B2(n_49618),
    .Y(n_51039));
 AOI22xp33_ASAP7_75t_SL g200839 (.A1(\u7_mem[0] [16]),
    .A2(n_49129),
    .B1(n_63785),
    .B2(\u7_mem[2] [16]),
    .Y(n_51040));
 AO22x1_ASAP7_75t_SL g200840 (.A1(n_49129),
    .A2(\u7_mem[0] [19]),
    .B1(n_63785),
    .B2(\u7_mem[2] [19]),
    .Y(n_51041));
 AOI22xp33_ASAP7_75t_SL g200841 (.A1(n_49618),
    .A2(\u7_mem[3] [5]),
    .B1(n_63785),
    .B2(\u7_mem[2] [5]),
    .Y(n_51042));
 AOI22xp33_ASAP7_75t_SL g200844 (.A1(n_49129),
    .A2(\u7_mem[0] [11]),
    .B1(\u7_mem[2] [11]),
    .B2(n_63785),
    .Y(n_51045));
 AOI22xp5_ASAP7_75t_SL g200845 (.A1(\u7_mem[0] [9]),
    .A2(n_49129),
    .B1(\u7_mem[2] [9]),
    .B2(n_63785),
    .Y(n_51046));
 AOI22xp5_ASAP7_75t_SL g200846 (.A1(\u7_mem[0] [8]),
    .A2(n_49129),
    .B1(\u7_mem[2] [8]),
    .B2(n_63785),
    .Y(n_51047));
 AOI22xp5_ASAP7_75t_SL g200847 (.A1(\u7_mem[0] [18]),
    .A2(n_49129),
    .B1(\u7_mem[2] [18]),
    .B2(n_63785),
    .Y(n_51048));
 AOI22xp5_ASAP7_75t_SL g200848 (.A1(\u7_mem[0] [10]),
    .A2(n_49129),
    .B1(\u7_mem[2] [10]),
    .B2(n_63785),
    .Y(n_51049));
 AOI22xp5_ASAP7_75t_SL g200850 (.A1(\u7_mem[0] [0]),
    .A2(n_49129),
    .B1(\u7_mem[2] [0]),
    .B2(n_63785),
    .Y(n_51051));
 AND2x4_ASAP7_75t_SL g200851_dup (.A(n_63785),
    .B(n_53365),
    .Y(n_53370));
 AOI22xp33_ASAP7_75t_SL g200852 (.A1(\u7_mem[0] [17]),
    .A2(n_49129),
    .B1(n_63785),
    .B2(\u7_mem[2] [17]),
    .Y(n_51053));
 BUFx3_ASAP7_75t_SL g200936 (.A(n_42248),
    .Y(n_51158));
 NAND2xp5_ASAP7_75t_SL g200938 (.A(n_51158),
    .B(out_slt8[13]),
    .Y(n_51159));
 HB1xp67_ASAP7_75t_L g201204 (.A(n_79178),
    .Y(n_51478));
 AOI22xp5_ASAP7_75t_SL g201208 (.A1(n_79178),
    .A2(\u8_mem[2] [0]),
    .B1(n_78273),
    .B2(\u8_mem[3] [0]),
    .Y(n_51481));
 AOI22xp33_ASAP7_75t_SL g201209 (.A1(n_79178),
    .A2(\u8_mem[2] [2]),
    .B1(n_78273),
    .B2(\u8_mem[3] [2]),
    .Y(n_51482));
 AOI22xp5_ASAP7_75t_SL g201210 (.A1(n_79178),
    .A2(\u8_mem[2] [15]),
    .B1(\u8_mem[3] [15]),
    .B2(n_78273),
    .Y(n_51483));
 AOI22xp5_ASAP7_75t_SL g201211 (.A1(n_79178),
    .A2(\u8_mem[2] [1]),
    .B1(n_78273),
    .B2(\u8_mem[3] [1]),
    .Y(n_51484));
 AOI22xp33_ASAP7_75t_SL g201213 (.A1(n_70885),
    .A2(\u8_mem[0] [16]),
    .B1(n_79178),
    .B2(\u8_mem[2] [16]),
    .Y(n_51486));
 AOI22xp5_ASAP7_75t_SL g201214 (.A1(n_79178),
    .A2(\u8_mem[2] [18]),
    .B1(n_78273),
    .B2(\u8_mem[3] [18]),
    .Y(n_51487));
 AND2x4_ASAP7_75t_SL g201215 (.A(n_636),
    .B(n_79178),
    .Y(n_51488));
 AOI22xp5_ASAP7_75t_SL g201216 (.A1(n_79178),
    .A2(\u8_mem[2] [17]),
    .B1(n_78273),
    .B2(\u8_mem[3] [17]),
    .Y(n_51489));
 AOI22xp5_ASAP7_75t_SL g201217 (.A1(\u8_mem[0] [5]),
    .A2(n_70885),
    .B1(n_79178),
    .B2(\u8_mem[2] [5]),
    .Y(n_51490));
 AOI22xp5_ASAP7_75t_SL g201220 (.A1(n_70885),
    .A2(\u8_mem[0] [7]),
    .B1(n_79178),
    .B2(\u8_mem[2] [7]),
    .Y(n_51493));
 AOI22xp33_ASAP7_75t_SL g201222 (.A1(n_79178),
    .A2(\u8_mem[2] [3]),
    .B1(n_78273),
    .B2(\u8_mem[3] [3]),
    .Y(n_51495));
 AOI22xp5_ASAP7_75t_SL g201223 (.A1(\u8_mem[0] [19]),
    .A2(n_70885),
    .B1(n_79178),
    .B2(\u8_mem[2] [19]),
    .Y(n_51496));
 AOI22xp5_ASAP7_75t_SL g201225 (.A1(n_79178),
    .A2(\u8_mem[2] [8]),
    .B1(\u8_mem[0] [8]),
    .B2(n_59474),
    .Y(n_51498));
 AOI22xp5_ASAP7_75t_SL g201226 (.A1(n_79178),
    .A2(\u8_mem[2] [11]),
    .B1(\u8_mem[3] [11]),
    .B2(n_78273),
    .Y(n_51499));
 AOI22xp5_ASAP7_75t_SL g201227 (.A1(\u8_mem[2] [4]),
    .A2(n_79178),
    .B1(\u8_mem[0] [4]),
    .B2(n_70885),
    .Y(n_51500));
 NAND2x1_ASAP7_75t_SL g202202 (.A(n_52768),
    .B(n_52769),
    .Y(n_52770));
 AND3x2_ASAP7_75t_SL g202203 (.A(n_370),
    .B(n_624),
    .C(n_36068),
    .Y(n_52769));
 AOI22xp5_ASAP7_75t_SL g202272 (.A1(\u5_mem[0] [1]),
    .A2(n_53101),
    .B1(\u5_mem[2] [1]),
    .B2(n_65643),
    .Y(n_52880));
 AOI22xp5_ASAP7_75t_SL g202287 (.A1(n_52893),
    .A2(n_66856),
    .B1(\u3_mem[0] [3]),
    .B2(n_51296),
    .Y(n_52895));
 AOI22xp5_ASAP7_75t_SL g202288 (.A1(n_52893),
    .A2(n_10891),
    .B1(\u3_mem[0] [1]),
    .B2(n_51296),
    .Y(n_52896));
 AOI22xp5_ASAP7_75t_SL g202289 (.A1(n_52893),
    .A2(n_66016),
    .B1(\u3_mem[0] [21]),
    .B2(n_51296),
    .Y(n_52897));
 AOI22xp5_ASAP7_75t_SL g202290 (.A1(n_52898),
    .A2(n_66004),
    .B1(\u3_mem[0] [6]),
    .B2(n_51288),
    .Y(n_52899));
 AOI22xp5_ASAP7_75t_SL g202292 (.A1(n_52893),
    .A2(n_66842),
    .B1(\u3_mem[0] [11]),
    .B2(n_51296),
    .Y(n_52900));
 AOI22xp5_ASAP7_75t_SL g202293 (.A1(n_52893),
    .A2(n_65952),
    .B1(\u3_mem[0] [17]),
    .B2(n_51288),
    .Y(n_52901));
 AOI22xp5_ASAP7_75t_SL g202294 (.A1(n_52893),
    .A2(n_65969),
    .B1(\u3_mem[0] [7]),
    .B2(n_51296),
    .Y(n_52902));
 AOI22xp5_ASAP7_75t_SL g202295 (.A1(n_52893),
    .A2(n_65915),
    .B1(\u3_mem[0] [24]),
    .B2(n_51288),
    .Y(n_52903));
 AOI22xp5_ASAP7_75t_SL g202297 (.A1(n_52893),
    .A2(n_10247),
    .B1(\u3_mem[0] [20]),
    .B2(n_51288),
    .Y(n_52905));
 AOI22xp5_ASAP7_75t_SL g202298 (.A1(n_52893),
    .A2(n_65925),
    .B1(\u3_mem[0] [25]),
    .B2(n_51288),
    .Y(n_52906));
 AOI22xp5_ASAP7_75t_SL g202299 (.A1(n_52893),
    .A2(n_35041),
    .B1(\u3_mem[0] [13]),
    .B2(n_51288),
    .Y(n_52907));
 AOI22xp5_ASAP7_75t_SL g202300 (.A1(n_52893),
    .A2(n_10638),
    .B1(\u3_mem[0] [30]),
    .B2(n_51296),
    .Y(n_52908));
 AOI22xp5_ASAP7_75t_SL g202301 (.A1(n_52893),
    .A2(n_28240),
    .B1(\u3_mem[0] [8]),
    .B2(n_51296),
    .Y(n_52909));
 AOI22xp5_ASAP7_75t_SL g202302 (.A1(n_52893),
    .A2(n_62940),
    .B1(\u3_mem[0] [27]),
    .B2(n_51288),
    .Y(n_52910));
 AOI22xp5_ASAP7_75t_SL g202303 (.A1(n_52898),
    .A2(n_9942),
    .B1(\u3_mem[0] [9]),
    .B2(n_51288),
    .Y(n_52911));
 AOI22xp5_ASAP7_75t_SL g202304 (.A1(n_52898),
    .A2(n_35437),
    .B1(\u3_mem[0] [26]),
    .B2(n_51296),
    .Y(n_52912));
 AOI22xp5_ASAP7_75t_SL g202305 (.A1(n_52898),
    .A2(n_10924),
    .B1(\u3_mem[0] [0]),
    .B2(n_51296),
    .Y(n_52913));
 AOI22xp5_ASAP7_75t_SL g202306 (.A1(n_52898),
    .A2(n_65920),
    .B1(\u3_mem[0] [28]),
    .B2(n_51296),
    .Y(n_52914));
 AOI22xp5_ASAP7_75t_SL g202307 (.A1(n_52898),
    .A2(n_10194),
    .B1(\u3_mem[0] [18]),
    .B2(n_51296),
    .Y(n_52915));
 AOI22xp5_ASAP7_75t_SL g202308 (.A1(n_52898),
    .A2(n_15920),
    .B1(\u3_mem[0] [31]),
    .B2(n_51288),
    .Y(n_52916));
 AOI22xp5_ASAP7_75t_SL g202309 (.A1(n_52898),
    .A2(n_22715),
    .B1(\u3_mem[0] [29]),
    .B2(n_51296),
    .Y(n_52917));
 AOI22xp5_ASAP7_75t_SL g202310 (.A1(n_52898),
    .A2(n_10196),
    .B1(\u3_mem[0] [19]),
    .B2(n_51296),
    .Y(n_52918));
 AOI22xp5_ASAP7_75t_SL g202311 (.A1(n_52898),
    .A2(n_28276),
    .B1(\u3_mem[0] [16]),
    .B2(n_51288),
    .Y(n_52919));
 AOI22xp5_ASAP7_75t_SL g202312 (.A1(n_52898),
    .A2(n_28913),
    .B1(\u3_mem[0] [15]),
    .B2(n_51296),
    .Y(n_52920));
 AOI22xp5_ASAP7_75t_SL g202313 (.A1(n_52898),
    .A2(n_65930),
    .B1(\u3_mem[0] [23]),
    .B2(n_51288),
    .Y(n_52921));
 AOI22xp5_ASAP7_75t_SL g202314 (.A1(n_52898),
    .A2(n_28251),
    .B1(\u3_mem[0] [14]),
    .B2(n_51288),
    .Y(n_52922));
 AOI22xp5_ASAP7_75t_SL g202315 (.A1(n_52898),
    .A2(n_10058),
    .B1(\u3_mem[0] [5]),
    .B2(n_51288),
    .Y(n_52923));
 AOI22xp5_ASAP7_75t_SL g202316 (.A1(n_52898),
    .A2(n_28330),
    .B1(\u3_mem[0] [2]),
    .B2(n_51288),
    .Y(n_52924));
 AOI22xp5_ASAP7_75t_SL g202318 (.A1(n_52898),
    .A2(n_10026),
    .B1(\u3_mem[0] [12]),
    .B2(n_51288),
    .Y(n_52926));
 NAND2xp5_ASAP7_75t_SL g202323 (.A(n_56844),
    .B(n_53102),
    .Y(n_52932));
 AOI21xp5_ASAP7_75t_SL g202325 (.A1(n_38368),
    .A2(n_31078),
    .B(n_52939),
    .Y(n_52940));
 AOI31xp33_ASAP7_75t_SL g202326 (.A1(n_52935),
    .A2(n_52936),
    .A3(n_52937),
    .B(n_52938),
    .Y(n_52939));
 AOI22xp33_ASAP7_75t_SL g202327 (.A1(n_7672),
    .A2(n_7673),
    .B1(n_698),
    .B2(n_65645),
    .Y(n_52935));
 AOI22xp33_ASAP7_75t_SL g202328 (.A1(n_698),
    .A2(n_29495),
    .B1(n_7672),
    .B2(n_7676),
    .Y(n_52936));
 NAND2xp33_ASAP7_75t_SL g202329 (.A(n_18704),
    .B(n_37200),
    .Y(n_52937));
 INVxp33_ASAP7_75t_L g202330 (.A(n_79104),
    .Y(n_52938));
 NAND3xp33_ASAP7_75t_SL g202336 (.A(n_52948),
    .B(n_52949),
    .C(n_52950),
    .Y(n_52951));
 AOI22xp5_ASAP7_75t_SL g202337 (.A1(i6_dout[15]),
    .A2(n_14933),
    .B1(i3_dout[15]),
    .B2(n_8341),
    .Y(n_52948));
 AOI221xp5_ASAP7_75t_SL g202338 (.A1(n_7082),
    .A2(u13_intm_r[15]),
    .B1(i4_dout[15]),
    .B2(n_8174),
    .C(n_10877),
    .Y(n_52949));
 AOI21xp33_ASAP7_75t_SL g202339 (.A1(n_10626),
    .A2(u13_ints_r[15]),
    .B(n_11015),
    .Y(n_52950));
 AOI21xp33_ASAP7_75t_SL g202359 (.A1(n_53003),
    .A2(n_37200),
    .B(n_52978),
    .Y(n_52979));
 OAI22xp5_ASAP7_75t_SL g202360 (.A1(n_4),
    .A2(n_64993),
    .B1(n_70),
    .B2(n_64994),
    .Y(n_52978));
 NAND2x1_ASAP7_75t_SL g202383 (.A(n_56858),
    .B(n_53002),
    .Y(n_53003));
 AOI22xp5_ASAP7_75t_SL g202384 (.A1(n_65642),
    .A2(\u5_mem[0] [9]),
    .B1(\u5_mem[2] [9]),
    .B2(n_65643),
    .Y(n_53002));
 AOI22xp33_ASAP7_75t_SL g202447 (.A1(\u5_mem[0] [3]),
    .A2(n_53101),
    .B1(n_65643),
    .B2(\u5_mem[2] [3]),
    .Y(n_53102));
 INVx3_ASAP7_75t_SL g202448 (.A(n_7872),
    .Y(n_53101));
 AND2x4_ASAP7_75t_SL g202672 (.A(u7_rp[0]),
    .B(n_50287),
    .Y(n_53365));
 AOI22xp33_ASAP7_75t_R g202673 (.A1(\u7_mem[2] [29]),
    .A2(n_53366),
    .B1(\u7_mem[3] [29]),
    .B2(n_73175),
    .Y(n_53367));
 AND2x2_ASAP7_75t_SL g202674 (.A(n_63785),
    .B(n_53365),
    .Y(n_53366));
 AOI22xp33_ASAP7_75t_R g202675 (.A1(\u7_mem[2] [28]),
    .A2(n_53366),
    .B1(\u7_mem[3] [28]),
    .B2(n_73175),
    .Y(n_53368));
 AOI22xp33_ASAP7_75t_L g202676 (.A1(\u7_mem[2] [31]),
    .A2(n_53366),
    .B1(\u7_mem[3] [31]),
    .B2(n_73175),
    .Y(n_53369));
 AOI22xp33_ASAP7_75t_L g202677 (.A1(\u7_mem[2] [27]),
    .A2(n_53370),
    .B1(\u7_mem[3] [27]),
    .B2(n_73175),
    .Y(n_53371));
 AOI22xp33_ASAP7_75t_L g202678 (.A1(\u7_mem[2] [30]),
    .A2(n_53370),
    .B1(\u7_mem[3] [30]),
    .B2(n_73175),
    .Y(n_53372));
 AOI22xp33_ASAP7_75t_SL g204759 (.A1(n_64744),
    .A2(n_50293),
    .B1(n_1840),
    .B2(n_50290),
    .Y(n_56059));
 AOI22xp5_ASAP7_75t_SL g204761 (.A1(n_63785),
    .A2(\u7_mem[2] [13]),
    .B1(\u7_mem[3] [13]),
    .B2(n_49618),
    .Y(n_56056));
 AOI22xp5_ASAP7_75t_SL g204762 (.A1(n_49129),
    .A2(\u7_mem[0] [13]),
    .B1(\u7_mem[1] [13]),
    .B2(n_49617),
    .Y(n_56057));
 NAND2xp5_ASAP7_75t_L g204763 (.A(n_50293),
    .B(n_64744),
    .Y(n_56060));
 INVxp67_ASAP7_75t_SL g204765 (.A(n_64744),
    .Y(n_56062));
 AND2x6_ASAP7_75t_SL g205395 (.A(u5_rp[1]),
    .B(u5_rp[2]),
    .Y(n_56842));
 AOI22xp33_ASAP7_75t_SL g205396 (.A1(n_64833),
    .A2(\u5_mem[1] [3]),
    .B1(n_56842),
    .B2(\u5_mem[3] [3]),
    .Y(n_56844));
 AOI22xp5_ASAP7_75t_SL g205397 (.A1(n_64833),
    .A2(\u5_mem[1] [2]),
    .B1(\u5_mem[3] [2]),
    .B2(n_56842),
    .Y(n_56845));
 AOI22xp5_ASAP7_75t_SL g205398 (.A1(n_31895),
    .A2(\u5_mem[1] [0]),
    .B1(\u5_mem[3] [0]),
    .B2(n_56842),
    .Y(n_56846));
 AOI22xp5_ASAP7_75t_SL g205399 (.A1(n_64833),
    .A2(\u5_mem[1] [16]),
    .B1(\u5_mem[3] [16]),
    .B2(n_56842),
    .Y(n_56847));
 AOI22xp5_ASAP7_75t_SL g205400 (.A1(n_31895),
    .A2(\u5_mem[1] [1]),
    .B1(\u5_mem[3] [1]),
    .B2(n_56842),
    .Y(n_56848));
 AOI22xp33_ASAP7_75t_SL g205401 (.A1(\u5_mem[1] [12]),
    .A2(n_31895),
    .B1(n_56842),
    .B2(\u5_mem[3] [12]),
    .Y(n_56849));
 XOR2xp5_ASAP7_75t_L g205402 (.A(u5_rp[3]),
    .B(n_56842),
    .Y(n_56850));
 AOI22xp5_ASAP7_75t_SL g205403 (.A1(\u5_mem[2] [7]),
    .A2(n_65643),
    .B1(\u5_mem[3] [7]),
    .B2(n_56842),
    .Y(n_56851));
 AOI22xp33_ASAP7_75t_SL g205404 (.A1(n_65643),
    .A2(\u5_mem[2] [5]),
    .B1(n_56842),
    .B2(\u5_mem[3] [5]),
    .Y(n_56852));
 AOI22xp33_ASAP7_75t_SL g205405 (.A1(\u5_mem[2] [19]),
    .A2(n_65643),
    .B1(\u5_mem[3] [19]),
    .B2(n_56842),
    .Y(n_56853));
 AOI22xp33_ASAP7_75t_SL g205406 (.A1(\u5_mem[2] [15]),
    .A2(n_65643),
    .B1(\u5_mem[3] [15]),
    .B2(n_56842),
    .Y(n_56854));
 AOI22xp33_ASAP7_75t_SL g205407 (.A1(n_65643),
    .A2(\u5_mem[2] [11]),
    .B1(n_56842),
    .B2(\u5_mem[3] [11]),
    .Y(n_56855));
 AOI22xp5_ASAP7_75t_L g205408 (.A1(n_65643),
    .A2(\u5_mem[2] [10]),
    .B1(\u5_mem[3] [10]),
    .B2(n_56842),
    .Y(n_56856));
 NAND2x1_ASAP7_75t_SL g205409 (.A(u5_rp[0]),
    .B(n_56842),
    .Y(n_56857));
 AOI22xp5_ASAP7_75t_SL g205410 (.A1(\u5_mem[3] [9]),
    .A2(n_56842),
    .B1(n_64833),
    .B2(\u5_mem[1] [9]),
    .Y(n_56858));
 AOI22xp5_ASAP7_75t_SL g205411 (.A1(n_64833),
    .A2(\u5_mem[1] [17]),
    .B1(\u5_mem[3] [17]),
    .B2(n_56842),
    .Y(n_56859));
 AOI22xp33_ASAP7_75t_SL g205412 (.A1(\u5_mem[2] [6]),
    .A2(n_65643),
    .B1(n_56842),
    .B2(\u5_mem[3] [6]),
    .Y(n_56860));
 AOI22xp5_ASAP7_75t_L g205413 (.A1(n_65643),
    .A2(\u5_mem[2] [14]),
    .B1(n_56842),
    .B2(\u5_mem[3] [14]),
    .Y(n_56861));
 AOI22xp33_ASAP7_75t_L g205415 (.A1(\u5_mem[2] [13]),
    .A2(n_65643),
    .B1(\u5_mem[3] [13]),
    .B2(n_56842),
    .Y(n_56863));
 AOI22xp33_ASAP7_75t_SL g205416 (.A1(\u5_mem[2] [4]),
    .A2(n_65643),
    .B1(n_56842),
    .B2(\u5_mem[3] [4]),
    .Y(n_56864));
 AND2x4_ASAP7_75t_SL g205417 (.A(n_7668),
    .B(n_56842),
    .Y(n_56865));
 NAND2xp5_ASAP7_75t_SL g205419 (.A(n_56866),
    .B(n_56867),
    .Y(n_56868));
 AOI22xp33_ASAP7_75t_SL g205420 (.A1(n_49129),
    .A2(\u7_mem[0] [1]),
    .B1(\u7_mem[2] [1]),
    .B2(n_63785),
    .Y(n_56866));
 AOI22xp5_ASAP7_75t_SL g205421 (.A1(n_49617),
    .A2(\u7_mem[1] [1]),
    .B1(\u7_mem[3] [1]),
    .B2(n_49618),
    .Y(n_56867));
 NAND2xp5_ASAP7_75t_SL g205423 (.A(n_56868),
    .B(n_50290),
    .Y(n_56871));
 AND2x2_ASAP7_75t_L g205517 (.A(n_65292),
    .B(n_78002),
    .Y(n_57041));
 INVx2_ASAP7_75t_SL g205538 (.A(n_636),
    .Y(n_57084));
 NAND2x1_ASAP7_75t_SL g205710 (.A(n_51498),
    .B(n_64672),
    .Y(n_57289));
 A2O1A1Ixp33_ASAP7_75t_SL g206130 (.A1(n_6144),
    .A2(n_50290),
    .B(n_64716),
    .C(n_52769),
    .Y(n_57733));
 AOI21xp5_ASAP7_75t_SL g206149 (.A1(n_57758),
    .A2(n_57759),
    .B(n_2753),
    .Y(n_57760));
 NAND2xp33_ASAP7_75t_SL g206150 (.A(n_2752),
    .B(n_29361),
    .Y(n_57758));
 NAND2xp33_ASAP7_75t_L g206151 (.A(n_29362),
    .B(o8_we),
    .Y(n_57759));
 AOI221xp5_ASAP7_75t_SL g206337 (.A1(n_57963),
    .A2(n_57964),
    .B1(n_20673),
    .B2(n_50109),
    .C(n_57965),
    .Y(n_57966));
 INVx1_ASAP7_75t_SL g206338 (.A(n_20673),
    .Y(n_57963));
 INVx2_ASAP7_75t_SL g206339 (.A(oc3_cfg[0]),
    .Y(n_57965));
 NAND2xp5_ASAP7_75t_SL g206949 (.A(n_58646),
    .B(n_58649),
    .Y(n_58650));
 INVx1_ASAP7_75t_L g206950 (.A(n_21024),
    .Y(n_58646));
 NOR2x1_ASAP7_75t_SL g206951 (.A(n_58647),
    .B(n_58648),
    .Y(n_58649));
 NAND2xp5_ASAP7_75t_SL g206952 (.A(n_36068),
    .B(n_34473),
    .Y(n_58647));
 NAND2xp5_ASAP7_75t_SL g206953 (.A(n_78094),
    .B(n_34472),
    .Y(n_58648));
 A2O1A1Ixp33_ASAP7_75t_SL g207000 (.A1(n_7665),
    .A2(n_4318),
    .B(n_38364),
    .C(n_66668),
    .Y(n_58710));
 AOI22xp5_ASAP7_75t_SL g207116 (.A1(\u4_mem[0] [10]),
    .A2(n_58959),
    .B1(\u4_mem[2] [10]),
    .B2(n_35632),
    .Y(n_58960));
 INVx5_ASAP7_75t_SL g207117 (.A(n_415),
    .Y(n_58959));
 INVx1_ASAP7_75t_R g207382 (.A(\u7_mem[2] [20]),
    .Y(n_59252));
 INVx3_ASAP7_75t_SL g207385 (.A(n_73175),
    .Y(n_59256));
 OAI21xp5_ASAP7_75t_SL g207467 (.A1(n_59338),
    .A2(n_59339),
    .B(n_59340),
    .Y(n_59341));
 INVx1_ASAP7_75t_SL g207468 (.A(\u5_mem[2] [29]),
    .Y(n_59338));
 INVx2_ASAP7_75t_SL g207469 (.A(n_1459),
    .Y(n_59339));
 NAND2xp5_ASAP7_75t_L g207470 (.A(\u5_mem[3] [29]),
    .B(n_56865),
    .Y(n_59340));
 AND2x4_ASAP7_75t_SL g207595 (.A(n_72057),
    .B(n_53263),
    .Y(n_59474));
 NAND2xp5_ASAP7_75t_SL g207597 (.A(n_59476),
    .B(n_51484),
    .Y(n_59477));
 AOI22xp33_ASAP7_75t_SL g207598 (.A1(n_59474),
    .A2(\u8_mem[0] [1]),
    .B1(n_78274),
    .B2(\u8_mem[1] [1]),
    .Y(n_59476));
 INVx1_ASAP7_75t_SL g207748 (.A(n_52932),
    .Y(n_59640));
 NAND2xp5_ASAP7_75t_SL g207749 (.A(n_643),
    .B(n_21015),
    .Y(n_59641));
 NAND2xp5_ASAP7_75t_R g207750 (.A(n_698),
    .B(n_42031),
    .Y(n_59642));
 INVx1_ASAP7_75t_SL g207751 (.A(n_698),
    .Y(n_59644));
 AOI22xp33_ASAP7_75t_SL g207843 (.A1(\u3_mem[2] [29]),
    .A2(n_77398),
    .B1(\u3_mem[3] [29]),
    .B2(n_22062),
    .Y(n_59759));
 OAI22xp5_ASAP7_75t_SL g207848 (.A1(u2_res_cnt[0]),
    .A2(n_31535),
    .B1(n_59763),
    .B2(n_1920),
    .Y(n_59764));
 INVx2_ASAP7_75t_SL g207849 (.A(n_31535),
    .Y(n_59763));
 AOI22xp5_ASAP7_75t_SL g208465 (.A1(\u10_mem[1] [29]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4693),
    .Y(n_60456));
 AOI22xp5_ASAP7_75t_SL g208588 (.A1(\u6_mem[3] [14]),
    .A2(n_77233),
    .B1(n_66032),
    .B2(n_61228),
    .Y(n_60588));
 AOI22xp33_ASAP7_75t_SL g208862 (.A1(n_60873),
    .A2(\u9_mem[1] [1]),
    .B1(n_24734),
    .B2(n_12482),
    .Y(n_60874));
 OR2x6_ASAP7_75t_SL g208863 (.A(n_24736),
    .B(n_203),
    .Y(n_60873));
 AOI22xp5_ASAP7_75t_SL g209203 (.A1(\u6_mem[3] [7]),
    .A2(n_77233),
    .B1(n_65969),
    .B2(n_61228),
    .Y(n_61229));
 INVx8_ASAP7_75t_SL g209205 (.A(n_35215),
    .Y(n_61228));
 AOI22xp5_ASAP7_75t_SL g209218 (.A1(n_61242),
    .A2(n_61243),
    .B1(\u10_mem[3] [11]),
    .B2(n_61244),
    .Y(n_61245));
 AND2x6_ASAP7_75t_SL g209219 (.A(n_33604),
    .B(n_33603),
    .Y(n_61242));
 OR2x6_ASAP7_75t_SL g209220 (.A(n_24975),
    .B(n_534),
    .Y(n_61244));
 AOI22xp5_ASAP7_75t_SL g209708 (.A1(\u11_mem[2] [20]),
    .A2(n_61785),
    .B1(n_4899),
    .B2(n_45625),
    .Y(n_61773));
 AOI22xp5_ASAP7_75t_SL g209721 (.A1(\u11_mem[2] [0]),
    .A2(n_61785),
    .B1(n_66076),
    .B2(n_28520),
    .Y(n_61786));
 OR2x6_ASAP7_75t_SL g209722 (.A(n_23286),
    .B(n_23285),
    .Y(n_61785));
 AOI22xp5_ASAP7_75t_SL g209801 (.A1(\u10_mem[1] [10]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_46479),
    .Y(n_61883));
 AOI22xp5_ASAP7_75t_SL g209803 (.A1(\u10_mem[1] [3]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_35392),
    .Y(n_61885));
 AOI22xp5_ASAP7_75t_SL g209805 (.A1(\u10_mem[1] [1]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_48456),
    .Y(n_61887));
 AOI22xp5_ASAP7_75t_SL g209807 (.A1(\u10_mem[1] [0]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_40956),
    .Y(n_61889));
 AOI22xp5_ASAP7_75t_SL g209813 (.A1(\u10_mem[1] [20]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4675),
    .Y(n_61895));
 AOI22xp5_ASAP7_75t_SL g209819 (.A1(\u10_mem[1] [22]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4671),
    .Y(n_61901));
 AOI22xp5_ASAP7_75t_SL g209875 (.A1(\u10_mem[1] [28]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4695),
    .Y(n_61957));
 AOI22xp5_ASAP7_75t_SL g209881 (.A1(\u10_mem[1] [25]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4665),
    .Y(n_61963));
 INVx4_ASAP7_75t_SL g21 (.A(u10_wp[1]),
    .Y(n_25438));
 AOI22xp5_ASAP7_75t_SL g210032 (.A1(\u10_mem[1] [24]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_4667),
    .Y(n_62124));
 AOI22xp5_ASAP7_75t_SL g210417 (.A1(n_62614),
    .A2(n_36971),
    .B1(\u10_mem[2] [2]),
    .B2(n_48153),
    .Y(n_62615));
 NAND2x1_ASAP7_75t_SL g210418 (.A(n_62612),
    .B(n_62613),
    .Y(n_62614));
 AOI22xp5_ASAP7_75t_SL g210419 (.A1(in_slt4[4]),
    .A2(n_1666),
    .B1(u10_din_tmp1[2]),
    .B2(n_24336),
    .Y(n_62612));
 NAND2xp5_ASAP7_75t_SL g210420 (.A(in_slt4[2]),
    .B(n_1667),
    .Y(n_62613));
 AOI22xp5_ASAP7_75t_SL g210439 (.A1(crac_out[21]),
    .A2(n_56881),
    .B1(n_73996),
    .B2(n_17579),
    .Y(n_62634));
 AOI22xp5_ASAP7_75t_SL g210458 (.A1(\u10_mem[1] [2]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_62614),
    .Y(n_62657));
 O2A1O1Ixp5_ASAP7_75t_SL g210505 (.A1(n_64974),
    .A2(n_62717),
    .B(n_5077),
    .C(n_4471),
    .Y(n_62718));
 NAND2xp5_ASAP7_75t_L g210507 (.A(n_2401),
    .B(n_53367),
    .Y(n_62717));
 BUFx3_ASAP7_75t_R g210669 (.A(out_slt0[9]),
    .Y(n_62918));
 BUFx12f_ASAP7_75t_SL g210670 (.A(n_36068),
    .Y(n_62919));
 NAND2xp5_ASAP7_75t_SL g210671 (.A(n_62919),
    .B(n_62918),
    .Y(n_62920));
 INVx3_ASAP7_75t_SL g210690 (.A(n_10486),
    .Y(n_62940));
 AOI22xp5_ASAP7_75t_SL g211398 (.A1(\u6_mem[2] [13]),
    .A2(n_77853),
    .B1(\u6_mem[3] [13]),
    .B2(n_41152),
    .Y(n_63778));
 AOI22xp5_ASAP7_75t_SL g211406 (.A1(\u7_mem[2] [14]),
    .A2(n_63785),
    .B1(\u7_mem[3] [14]),
    .B2(n_49618),
    .Y(n_63786));
 AND2x6_ASAP7_75t_SL g211407 (.A(u7_rp[2]),
    .B(n_51030),
    .Y(n_63785));
 NAND2xp5_ASAP7_75t_SL g211605 (.A(n_2073),
    .B(n_63999),
    .Y(n_64000));
 AND2x4_ASAP7_75t_SL g211606 (.A(n_76054),
    .B(n_31535),
    .Y(n_63999));
 OA21x2_ASAP7_75t_SL g211697 (.A1(n_247),
    .A2(n_50293),
    .B(n_70324),
    .Y(n_64102));
 OAI21xp33_ASAP7_75t_SL g211698 (.A1(n_247),
    .A2(n_50293),
    .B(n_70324),
    .Y(n_64103));
 INVxp33_ASAP7_75t_R g211860 (.A(dma_ack_i[2]),
    .Y(n_64296));
 AOI22xp5_ASAP7_75t_SL g212080 (.A1(\u8_mem[1] [8]),
    .A2(n_78274),
    .B1(\u8_mem[3] [8]),
    .B2(n_78273),
    .Y(n_64672));
 NOR2xp33_ASAP7_75t_L g212105 (.A(n_64696),
    .B(n_330),
    .Y(n_64697));
 INVx1_ASAP7_75t_L g212106 (.A(in_slt4[7]),
    .Y(n_64696));
 INVxp33_ASAP7_75t_SL g212117 (.A(n_64710),
    .Y(n_64711));
 NAND2xp5_ASAP7_75t_SL g212118 (.A(n_64708),
    .B(n_64709),
    .Y(n_64710));
 AOI22xp5_ASAP7_75t_SL g212119 (.A1(n_65642),
    .A2(\u5_mem[0] [8]),
    .B1(\u5_mem[1] [8]),
    .B2(n_31895),
    .Y(n_64708));
 AOI22xp33_ASAP7_75t_SL g212120 (.A1(\u5_mem[2] [8]),
    .A2(n_65643),
    .B1(\u5_mem[3] [8]),
    .B2(n_56842),
    .Y(n_64709));
 NAND2xp5_ASAP7_75t_SL g212122 (.A(n_2188),
    .B(n_64710),
    .Y(n_64713));
 NOR2xp33_ASAP7_75t_SL g212123 (.A(n_64714),
    .B(n_64715),
    .Y(n_64716));
 INVx2_ASAP7_75t_SL g212124 (.A(n_51030),
    .Y(n_64714));
 INVx4_ASAP7_75t_SL g212125 (.A(n_53365),
    .Y(n_64715));
 AOI22xp33_ASAP7_75t_SL g212183 (.A1(\u5_mem[0] [22]),
    .A2(n_64793),
    .B1(\u5_mem[1] [22]),
    .B2(n_6071),
    .Y(n_64794));
 INVx2_ASAP7_75t_SL g212184 (.A(n_64994),
    .Y(n_64793));
 NAND3xp33_ASAP7_75t_SL g212201 (.A(n_64812),
    .B(n_2403),
    .C(n_53368),
    .Y(n_64813));
 AOI222xp33_ASAP7_75t_SL g212202 (.A1(n_35407),
    .A2(n_50290),
    .B1(n_65056),
    .B2(\u7_mem[1] [28]),
    .C1(n_65055),
    .C2(\u7_mem[0] [28]),
    .Y(n_64812));
 BUFx3_ASAP7_75t_SL g212204 (.A(u8_wp[1]),
    .Y(n_64814));
 INVx1_ASAP7_75t_SL g212205 (.A(u8_wp[1]),
    .Y(n_64816));
 AND2x4_ASAP7_75t_SL g212206 (.A(n_64817),
    .B(n_64191),
    .Y(n_64818));
 INVx2_ASAP7_75t_L g212207 (.A(n_64816),
    .Y(n_64817));
 AND2x4_ASAP7_75t_SL g212208 (.A(n_64817),
    .B(n_64191),
    .Y(n_64819));
 BUFx6f_ASAP7_75t_SL g212232_dup (.A(n_66658),
    .Y(n_66672));
 AOI21x1_ASAP7_75t_SL g212233 (.A1(n_58646),
    .A2(n_28691),
    .B(n_5748),
    .Y(n_64847));
 OAI21xp33_ASAP7_75t_SL g212234 (.A1(n_58650),
    .A2(n_27321),
    .B(n_66660),
    .Y(n_64851));
 NAND2xp5_ASAP7_75t_SL g212237 (.A(n_47706),
    .B(n_47707),
    .Y(n_64849));
 INVx5_ASAP7_75t_SL g212238 (.A(n_7772),
    .Y(n_64852));
 AOI21xp5_ASAP7_75t_SL g212239 (.A1(n_23131),
    .A2(n_32585),
    .B(n_64855),
    .Y(n_64856));
 OAI21xp33_ASAP7_75t_SL g212240 (.A1(n_64853),
    .A2(n_64852),
    .B(n_64854),
    .Y(n_64855));
 AOI21xp33_ASAP7_75t_SL g212241 (.A1(n_35461),
    .A2(n_23129),
    .B(n_20973),
    .Y(n_64853));
 NAND2xp33_ASAP7_75t_SL g212242 (.A(out_slt4[10]),
    .B(n_7781),
    .Y(n_64854));
 AOI22xp5_ASAP7_75t_SL g212247 (.A1(n_62940),
    .A2(n_64861),
    .B1(\u6_mem[3] [27]),
    .B2(n_72084),
    .Y(n_64862));
 INVx8_ASAP7_75t_SL g212248 (.A(n_67568),
    .Y(n_64861));
 AO21x1_ASAP7_75t_SL g212358 (.A1(n_64744),
    .A2(n_50290),
    .B(n_64745),
    .Y(n_64974));
 OR2x2_ASAP7_75t_SL g212377 (.A(n_7872),
    .B(n_589),
    .Y(n_64994));
 AOI21xp33_ASAP7_75t_SL g212378 (.A1(n_64710),
    .A2(n_37200),
    .B(n_64997),
    .Y(n_64998));
 OAI22xp5_ASAP7_75t_SL g212379 (.A1(n_64993),
    .A2(n_64995),
    .B1(n_64996),
    .B2(n_64994),
    .Y(n_64997));
 INVxp67_ASAP7_75t_R g212380 (.A(\u5_mem[1] [24]),
    .Y(n_64995));
 INVxp67_ASAP7_75t_R g212381 (.A(\u5_mem[0] [24]),
    .Y(n_64996));
 AND2x2_ASAP7_75t_SL g212383 (.A(n_36635),
    .B(n_56861),
    .Y(n_65000));
 NAND2xp33_ASAP7_75t_SL g212384 (.A(n_36635),
    .B(n_56861),
    .Y(n_65001));
 OAI22xp5_ASAP7_75t_SL g212411 (.A1(n_6),
    .A2(n_59256),
    .B1(n_65029),
    .B2(n_116),
    .Y(n_65030));
 INVx4_ASAP7_75t_SL g212412 (.A(n_53370),
    .Y(n_65029));
 NOR2xp67_ASAP7_75t_SL g212429 (.A(n_73177),
    .B(n_65053),
    .Y(n_65054));
 AO22x1_ASAP7_75t_SL g212430 (.A1(n_65055),
    .A2(\u7_mem[0] [20]),
    .B1(\u7_mem[1] [20]),
    .B2(n_65056),
    .Y(n_65053));
 AND2x4_ASAP7_75t_SL g212432 (.A(n_53365),
    .B(n_49617),
    .Y(n_65056));
 NOR2xp67_ASAP7_75t_SL g212433 (.A(n_1789),
    .B(n_65057),
    .Y(n_65058));
 AO22x1_ASAP7_75t_SL g212434 (.A1(n_65055),
    .A2(\u7_mem[0] [23]),
    .B1(\u7_mem[1] [23]),
    .B2(n_65056),
    .Y(n_65057));
 AOI22xp5_ASAP7_75t_SL g212588 (.A1(n_66010),
    .A2(n_48109),
    .B1(n_65763),
    .B2(\u4_mem[1] [26]),
    .Y(n_65238));
 AND2x4_ASAP7_75t_SL g212590 (.A(n_35904),
    .B(n_24628),
    .Y(n_65236));
 AOI22xp5_ASAP7_75t_SL g212591 (.A1(n_65908),
    .A2(n_48109),
    .B1(n_65239),
    .B2(\u4_mem[1] [27]),
    .Y(n_65240));
 AOI22xp5_ASAP7_75t_SL g212593 (.A1(n_15920),
    .A2(n_48107),
    .B1(n_65239),
    .B2(\u4_mem[1] [31]),
    .Y(n_65241));
 AOI22xp5_ASAP7_75t_SL g212594 (.A1(n_28424),
    .A2(n_48109),
    .B1(n_65239),
    .B2(\u4_mem[1] [24]),
    .Y(n_65242));
 AOI22xp5_ASAP7_75t_SL g212595 (.A1(n_65930),
    .A2(n_48107),
    .B1(n_65239),
    .B2(\u4_mem[1] [23]),
    .Y(n_65243));
 AOI22xp5_ASAP7_75t_SL g212596 (.A1(n_65955),
    .A2(n_48109),
    .B1(n_65239),
    .B2(\u4_mem[1] [13]),
    .Y(n_65244));
 AOI22xp5_ASAP7_75t_SL g212597 (.A1(n_15867),
    .A2(n_48107),
    .B1(\u4_mem[1] [3]),
    .B2(n_65239),
    .Y(n_65245));
 AOI22xp5_ASAP7_75t_SL g212598 (.A1(n_66000),
    .A2(n_48109),
    .B1(\u4_mem[1] [2]),
    .B2(n_65239),
    .Y(n_65246));
 AOI22xp5_ASAP7_75t_SL g212599 (.A1(n_66032),
    .A2(n_48109),
    .B1(\u4_mem[1] [14]),
    .B2(n_65239),
    .Y(n_65247));
 AOI22xp5_ASAP7_75t_SL g212600 (.A1(n_28316),
    .A2(n_48107),
    .B1(\u4_mem[1] [25]),
    .B2(n_65239),
    .Y(n_65248));
 AOI22xp5_ASAP7_75t_SL g212601 (.A1(n_32916),
    .A2(n_48107),
    .B1(\u4_mem[1] [21]),
    .B2(n_65239),
    .Y(n_65249));
 AOI22xp5_ASAP7_75t_SL g212602 (.A1(n_33024),
    .A2(n_48109),
    .B1(\u4_mem[1] [20]),
    .B2(n_65239),
    .Y(n_65250));
 AOI22xp5_ASAP7_75t_SL g212603 (.A1(n_75733),
    .A2(n_48109),
    .B1(\u4_mem[1] [0]),
    .B2(n_65239),
    .Y(n_65251));
 AOI22xp5_ASAP7_75t_SL g212604 (.A1(n_10171),
    .A2(n_48109),
    .B1(\u4_mem[1] [18]),
    .B2(n_65239),
    .Y(n_65252));
 AOI22xp5_ASAP7_75t_SL g212605 (.A1(n_48109),
    .A2(n_10640),
    .B1(n_65763),
    .B2(\u4_mem[1] [30]),
    .Y(n_65253));
 AOI22xp5_ASAP7_75t_SL g212606 (.A1(n_65980),
    .A2(n_48109),
    .B1(\u4_mem[1] [8]),
    .B2(n_65763),
    .Y(n_65254));
 AOI22xp5_ASAP7_75t_SL g212607 (.A1(n_10000),
    .A2(n_48107),
    .B1(\u4_mem[1] [11]),
    .B2(n_65763),
    .Y(n_65255));
 AOI22xp5_ASAP7_75t_SL g212608 (.A1(n_65949),
    .A2(n_48109),
    .B1(\u4_mem[1] [16]),
    .B2(n_65763),
    .Y(n_65256));
 AOI22xp5_ASAP7_75t_SL g212609 (.A1(n_10143),
    .A2(n_48109),
    .B1(\u4_mem[1] [17]),
    .B2(n_65763),
    .Y(n_65257));
 AOI22xp5_ASAP7_75t_SL g212610 (.A1(n_10198),
    .A2(n_48107),
    .B1(\u4_mem[1] [19]),
    .B2(n_65763),
    .Y(n_65258));
 AOI22xp5_ASAP7_75t_SL g212612 (.A1(n_65920),
    .A2(n_48107),
    .B1(\u4_mem[1] [28]),
    .B2(n_65763),
    .Y(n_65260));
 AOI22xp5_ASAP7_75t_SL g212613 (.A1(n_32644),
    .A2(n_48109),
    .B1(\u4_mem[1] [6]),
    .B2(n_65763),
    .Y(n_65261));
 AOI22xp5_ASAP7_75t_SL g212614 (.A1(n_17578),
    .A2(n_48107),
    .B1(\u4_mem[1] [7]),
    .B2(n_65763),
    .Y(n_65262));
 AOI22xp5_ASAP7_75t_SL g212615 (.A1(n_65997),
    .A2(n_48107),
    .B1(\u4_mem[1] [12]),
    .B2(n_65763),
    .Y(n_65263));
 AOI22xp5_ASAP7_75t_SL g212617 (.A1(n_66868),
    .A2(n_48107),
    .B1(\u4_mem[1] [5]),
    .B2(n_65763),
    .Y(n_65265));
 AOI22xp5_ASAP7_75t_SL g212618 (.A1(n_79972),
    .A2(n_48109),
    .B1(n_65763),
    .B2(\u4_mem[1] [9]),
    .Y(n_65266));
 AOI22xp5_ASAP7_75t_SL g212619 (.A1(n_65941),
    .A2(n_48107),
    .B1(n_65763),
    .B2(\u4_mem[1] [22]),
    .Y(n_65267));
 AOI22xp5_ASAP7_75t_SL g212620 (.A1(n_28913),
    .A2(n_48109),
    .B1(n_65763),
    .B2(\u4_mem[1] [15]),
    .Y(n_65268));
 AOI22xp5_ASAP7_75t_SL g212621 (.A1(\u4_mem[1] [1]),
    .A2(n_65763),
    .B1(n_3815),
    .B2(n_48107),
    .Y(n_65269));
 AOI22xp5_ASAP7_75t_SL g212622 (.A1(n_48109),
    .A2(n_15952),
    .B1(n_65763),
    .B2(\u4_mem[1] [29]),
    .Y(n_65270));
 AND3x1_ASAP7_75t_SL g212625 (.A(n_21141),
    .B(n_672),
    .C(n_65297),
    .Y(n_65298));
 AOI22xp5_ASAP7_75t_SL g212626 (.A1(\u7_mem[3] [4]),
    .A2(n_49618),
    .B1(\u7_mem[2] [4]),
    .B2(n_63785),
    .Y(n_65297));
 INVx2_ASAP7_75t_SL g212652 (.A(u4_rp[3]),
    .Y(n_65325));
 NAND3xp33_ASAP7_75t_SL g212653 (.A(n_71395),
    .B(n_65328),
    .C(n_64014),
    .Y(n_65329));
 XNOR2xp5_ASAP7_75t_R g212654 (.A(n_65326),
    .B(n_65327),
    .Y(n_65328));
 NAND2xp5_ASAP7_75t_L g212655 (.A(n_30078),
    .B(n_71392),
    .Y(n_65326));
 XOR2xp5_ASAP7_75t_R g212656 (.A(n_65325),
    .B(u4_wp[2]),
    .Y(n_65327));
 NAND2xp5_ASAP7_75t_SL g212713 (.A(n_78959),
    .B(n_76764),
    .Y(n_65395));
 NAND2x1_ASAP7_75t_SL g212888 (.A(n_65577),
    .B(n_13983),
    .Y(n_65578));
 AOI22xp33_ASAP7_75t_SL g212889 (.A1(n_70885),
    .A2(\u8_mem[0] [9]),
    .B1(n_79178),
    .B2(\u8_mem[2] [9]),
    .Y(n_65577));
 AND2x4_ASAP7_75t_SL g212933 (.A(u5_rp[2]),
    .B(n_7869),
    .Y(n_65643));
 INVx1_ASAP7_75t_SL g212934 (.A(n_65644),
    .Y(n_65645));
 AOI22xp5_ASAP7_75t_SL g212935 (.A1(n_65642),
    .A2(\u5_mem[0] [16]),
    .B1(\u5_mem[2] [16]),
    .B2(n_65643),
    .Y(n_65644));
 AO21x1_ASAP7_75t_SL g212936 (.A1(n_56847),
    .A2(n_65644),
    .B(n_21026),
    .Y(n_65646));
 AOI22xp5_ASAP7_75t_SL g213021 (.A1(\u4_mem[1] [10]),
    .A2(n_65763),
    .B1(n_65975),
    .B2(n_48107),
    .Y(n_65764));
 INVx6_ASAP7_75t_SL g213022 (.A(n_65236),
    .Y(n_65763));
 NAND2xp5_ASAP7_75t_SL g213136 (.A(n_36478),
    .B(n_24337),
    .Y(n_65879));
 INVxp67_ASAP7_75t_R g213145 (.A(i3_dout[16]),
    .Y(n_65897));
 BUFx2_ASAP7_75t_R g213146 (.A(n_65899),
    .Y(n_65900));
 INVx3_ASAP7_75t_SL g213149 (.A(n_10330),
    .Y(n_65902));
 HB1xp67_ASAP7_75t_L g213155 (.A(n_65906),
    .Y(n_65910));
 INVxp67_ASAP7_75t_R g213156 (.A(n_10408),
    .Y(n_65914));
 INVx2_ASAP7_75t_SL g213157 (.A(n_65912),
    .Y(n_10408));
 INVx2_ASAP7_75t_SL g213160 (.A(n_10408),
    .Y(n_65915));
 BUFx2_ASAP7_75t_R g213162 (.A(n_65912),
    .Y(n_65917));
 BUFx3_ASAP7_75t_SL g213163 (.A(n_65919),
    .Y(n_65920));
 INVx1_ASAP7_75t_R g213166 (.A(n_10434),
    .Y(n_65924));
 INVx2_ASAP7_75t_SL g213167 (.A(n_65922),
    .Y(n_10434));
 INVxp33_ASAP7_75t_R g213170 (.A(wb_data_i[25]),
    .Y(n_65921));
 INVx2_ASAP7_75t_SL g213171 (.A(n_10434),
    .Y(n_65925));
 BUFx2_ASAP7_75t_R g213173 (.A(n_65922),
    .Y(n_65927));
 BUFx3_ASAP7_75t_SL g213174 (.A(n_65929),
    .Y(n_65930));
 INVxp33_ASAP7_75t_R g213177 (.A(wb_data_i[23]),
    .Y(n_65928));
 INVxp33_ASAP7_75t_R g213180 (.A(wb_data_i[19]),
    .Y(n_65931));
 BUFx3_ASAP7_75t_SL g213181 (.A(n_65934),
    .Y(n_10194));
 INVx2_ASAP7_75t_SL g213185 (.A(n_65937),
    .Y(n_10276));
 INVxp33_ASAP7_75t_R g213188 (.A(wb_data_i[22]),
    .Y(n_65936));
 INVx2_ASAP7_75t_SL g213193 (.A(n_10276),
    .Y(n_65941));
 BUFx4f_ASAP7_75t_SL g213196 (.A(n_65948),
    .Y(n_65949));
 BUFx4f_ASAP7_75t_SL g213199 (.A(n_65951),
    .Y(n_65952));
 INVxp33_ASAP7_75t_R g213204 (.A(wb_data_i[13]),
    .Y(n_65953));
 INVxp33_ASAP7_75t_R g213210 (.A(wb_data_i[5]),
    .Y(n_65958));
 INVxp33_ASAP7_75t_R g213214 (.A(wb_data_i[3]),
    .Y(n_65961));
 BUFx3_ASAP7_75t_SL g213218 (.A(n_65968),
    .Y(n_65969));
 INVxp33_ASAP7_75t_R g213223 (.A(wb_data_i[10]),
    .Y(n_65970));
 INVx2_ASAP7_75t_SL g213225 (.A(n_65971),
    .Y(n_9909));
 INVx2_ASAP7_75t_SL g213226 (.A(n_9909),
    .Y(n_65975));
 INVx3_ASAP7_75t_SL g213231 (.A(n_9880),
    .Y(n_65980));
 INVx2_ASAP7_75t_SL g213234 (.A(n_65984),
    .Y(n_9967));
 INVxp33_ASAP7_75t_R g213237 (.A(wb_data_i[4]),
    .Y(n_65983));
 BUFx3_ASAP7_75t_SL g213246 (.A(n_65996),
    .Y(n_65997));
 BUFx3_ASAP7_75t_SL g213249 (.A(n_65999),
    .Y(n_66000));
 INVxp33_ASAP7_75t_R g213254 (.A(wb_data_i[6]),
    .Y(n_66001));
 INVx2_ASAP7_75t_SL g213255 (.A(n_66003),
    .Y(n_66004));
 INVx1_ASAP7_75t_SL g213256 (.A(n_66002),
    .Y(n_66003));
 INVx2_ASAP7_75t_SL g213259 (.A(n_66008),
    .Y(n_10460));
 BUFx2_ASAP7_75t_R g213262 (.A(n_66008),
    .Y(n_66011));
 INVx3_ASAP7_75t_SL g213263 (.A(n_10460),
    .Y(n_66010));
 BUFx2_ASAP7_75t_L g213267 (.A(n_66015),
    .Y(n_66016));
 INVxp33_ASAP7_75t_R g213275 (.A(wb_data_i[20]),
    .Y(n_66023));
 INVx3_ASAP7_75t_SL g213276 (.A(n_66025),
    .Y(n_66026));
 INVx2_ASAP7_75t_L g213277 (.A(n_66024),
    .Y(n_66025));
 BUFx2_ASAP7_75t_L g213278 (.A(n_66024),
    .Y(n_10247));
 BUFx3_ASAP7_75t_SL g213281 (.A(n_66031),
    .Y(n_66032));
 XOR2xp5_ASAP7_75t_SL g213305 (.A(u9_wp[3]),
    .B(u9_rp[2]),
    .Y(n_66054));
 AO222x2_ASAP7_75t_SL g213327 (.A1(in_slt6[0]),
    .A2(n_46192),
    .B1(n_13236),
    .B2(u11_din_tmp1[0]),
    .C1(in_slt6[2]),
    .C2(n_1523),
    .Y(n_66076));
 AND2x2_ASAP7_75t_SL g213424 (.A(n_43395),
    .B(n_33792),
    .Y(n_66198));
 NAND2xp5_ASAP7_75t_SL g213425 (.A(n_43395),
    .B(n_33792),
    .Y(n_66199));
 AOI22xp33_ASAP7_75t_SL g213700 (.A1(n_66659),
    .A2(n_64848),
    .B1(n_64847),
    .B2(n_64849),
    .Y(n_66660));
 BUFx6f_ASAP7_75t_SL g213701 (.A(n_66658),
    .Y(n_66659));
 AOI21x1_ASAP7_75t_SL g213702 (.A1(n_34472),
    .A2(n_5789),
    .B(n_43100),
    .Y(n_66658));
 AND2x2_ASAP7_75t_R g213704 (.A(out_slt6[5]),
    .B(n_66659),
    .Y(n_66662));
 NAND2xp5_ASAP7_75t_R g213706 (.A(out_slt6[17]),
    .B(n_66659),
    .Y(n_66664));
 AOI222xp33_ASAP7_75t_SL g213707 (.A1(n_38363),
    .A2(n_18704),
    .B1(n_36224),
    .B2(n_22163),
    .C1(n_66659),
    .C2(out_slt6[2]),
    .Y(n_66665));
 NAND2xp5_ASAP7_75t_L g213708 (.A(n_66659),
    .B(out_slt6[14]),
    .Y(n_66666));
 NAND2xp5_ASAP7_75t_L g213709 (.A(out_slt6[11]),
    .B(n_66659),
    .Y(n_66667));
 NAND2xp5_ASAP7_75t_SL g213710 (.A(n_66659),
    .B(out_slt6[6]),
    .Y(n_66668));
 NAND2xp5_ASAP7_75t_R g213711 (.A(out_slt6[18]),
    .B(n_66659),
    .Y(n_66669));
 INVx2_ASAP7_75t_SL g213712 (.A(n_66659),
    .Y(n_66670));
 AND2x2_ASAP7_75t_R g213713 (.A(out_slt6[12]),
    .B(n_66659),
    .Y(n_66671));
 NAND2xp5_ASAP7_75t_R g213714 (.A(out_slt6[9]),
    .B(n_66672),
    .Y(n_66673));
 NAND2xp5_ASAP7_75t_R g213715 (.A(out_slt6[8]),
    .B(n_66672),
    .Y(n_66674));
 NOR2xp33_ASAP7_75t_SL g213716 (.A(n_66672),
    .B(n_64847),
    .Y(n_66675));
 AND2x2_ASAP7_75t_R g213717 (.A(out_slt6[7]),
    .B(n_66672),
    .Y(n_66676));
 NAND2xp5_ASAP7_75t_R g213718 (.A(out_slt6[16]),
    .B(n_66672),
    .Y(n_66677));
 AND2x2_ASAP7_75t_R g213719 (.A(out_slt6[13]),
    .B(n_66672),
    .Y(n_66678));
 AOI222xp33_ASAP7_75t_SL g213720 (.A1(n_38363),
    .A2(n_26098),
    .B1(n_22163),
    .B2(n_52932),
    .C1(n_66672),
    .C2(out_slt6[3]),
    .Y(n_66679));
 NAND2xp5_ASAP7_75t_SL g213721 (.A(n_66672),
    .B(out_slt6[10]),
    .Y(n_66680));
 NAND2xp5_ASAP7_75t_SL g213723 (.A(n_66672),
    .B(out_slt6[4]),
    .Y(n_66682));
 AOI22xp5_ASAP7_75t_SL g213724 (.A1(out_slt6[0]),
    .A2(n_66672),
    .B1(n_18704),
    .B2(n_28690),
    .Y(n_66683));
 AOI22xp33_ASAP7_75t_SL g213833 (.A1(crac_out[22]),
    .A2(n_56881),
    .B1(n_67246),
    .B2(n_12219),
    .Y(n_66799));
 AOI22xp5_ASAP7_75t_SL g213836 (.A1(n_3188),
    .A2(n_66801),
    .B1(\u7_mem[2] [22]),
    .B2(n_13325),
    .Y(n_66802));
 AOI22xp5_ASAP7_75t_SL g213837 (.A1(n_3420),
    .A2(n_67246),
    .B1(\u6_mem[0] [22]),
    .B2(n_3415),
    .Y(n_66803));
 AOI22xp5_ASAP7_75t_SL g213838 (.A1(n_67246),
    .A2(n_16797),
    .B1(n_16798),
    .B2(n_40824),
    .Y(n_66804));
 AOI22xp5_ASAP7_75t_SL g213839 (.A1(n_52898),
    .A2(n_67246),
    .B1(\u3_mem[0] [22]),
    .B2(n_51296),
    .Y(n_66805));
 AOI22xp5_ASAP7_75t_SL g213840 (.A1(n_67246),
    .A2(n_3461),
    .B1(\u8_mem[0] [22]),
    .B2(n_3453),
    .Y(n_66806));
 AOI22xp5_ASAP7_75t_SL g213841 (.A1(n_67246),
    .A2(n_32163),
    .B1(\u5_mem[1] [22]),
    .B2(n_13500),
    .Y(n_66807));
 AOI22xp5_ASAP7_75t_SL g213842 (.A1(n_3320),
    .A2(n_67246),
    .B1(\u8_mem[2] [22]),
    .B2(n_16900),
    .Y(n_66808));
 AOI22xp5_ASAP7_75t_SL g213843 (.A1(n_67246),
    .A2(n_43537),
    .B1(\u7_mem[1] [22]),
    .B2(n_50220),
    .Y(n_66809));
 AOI22xp5_ASAP7_75t_SL g213844 (.A1(n_24633),
    .A2(n_67246),
    .B1(\u4_mem[2] [22]),
    .B2(n_13304),
    .Y(n_66810));
 AOI22xp5_ASAP7_75t_SL g213846 (.A1(n_24806),
    .A2(n_67246),
    .B1(\u3_mem[2] [22]),
    .B2(n_15954),
    .Y(n_66812));
 AOI22xp5_ASAP7_75t_SL g213847 (.A1(n_12403),
    .A2(n_67246),
    .B1(\u7_mem[0] [22]),
    .B2(n_3365),
    .Y(n_66813));
 AOI22xp5_ASAP7_75t_SL g213848 (.A1(n_67246),
    .A2(n_6748),
    .B1(u13_intm_r[22]),
    .B2(n_32319),
    .Y(n_66814));
 AOI22xp5_ASAP7_75t_SL g213849 (.A1(n_29790),
    .A2(n_67246),
    .B1(\u4_mem[0] [22]),
    .B2(n_33655),
    .Y(n_66815));
 AOI22xp5_ASAP7_75t_SL g213850 (.A1(n_22577),
    .A2(\u3_mem[1] [22]),
    .B1(n_66801),
    .B2(n_15143),
    .Y(n_66816));
 AOI22xp5_ASAP7_75t_SL g213851 (.A1(n_66817),
    .A2(n_3454),
    .B1(\u8_mem[0] [10]),
    .B2(n_3453),
    .Y(n_66818));
 INVx5_ASAP7_75t_SL g213852 (.A(n_9909),
    .Y(n_66817));
 AOI22xp5_ASAP7_75t_SL g213853 (.A1(n_66817),
    .A2(n_32164),
    .B1(\u5_mem[1] [10]),
    .B2(n_13508),
    .Y(n_66819));
 AOI22xp5_ASAP7_75t_SL g213854 (.A1(crac_out[10]),
    .A2(n_28367),
    .B1(n_66817),
    .B2(n_17579),
    .Y(n_66820));
 AOI22xp5_ASAP7_75t_SL g213855 (.A1(\u6_mem[3] [10]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_66817),
    .Y(n_66821));
 AOI22xp5_ASAP7_75t_SL g213856 (.A1(n_66817),
    .A2(n_75734),
    .B1(n_31464),
    .B2(\u8_mem[1] [10]),
    .Y(n_66822));
 AOI22xp33_ASAP7_75t_SL g213858 (.A1(n_22577),
    .A2(\u3_mem[1] [10]),
    .B1(n_66824),
    .B2(n_16009),
    .Y(n_66825));
 AOI22xp5_ASAP7_75t_SL g213860 (.A1(n_3285),
    .A2(n_66817),
    .B1(\u5_mem[2] [10]),
    .B2(n_43028),
    .Y(n_66826));
 AOI22xp5_ASAP7_75t_SL g213861 (.A1(n_24633),
    .A2(n_66817),
    .B1(\u4_mem[2] [10]),
    .B2(n_13304),
    .Y(n_66827));
 AOI22xp5_ASAP7_75t_SL g213862 (.A1(n_3420),
    .A2(n_66817),
    .B1(\u6_mem[0] [10]),
    .B2(n_3415),
    .Y(n_66828));
 AOI22xp5_ASAP7_75t_SL g213863 (.A1(n_66817),
    .A2(n_12403),
    .B1(\u7_mem[0] [10]),
    .B2(n_3386),
    .Y(n_66829));
 AOI22xp5_ASAP7_75t_SL g213864 (.A1(n_477),
    .A2(n_26541),
    .B1(n_66817),
    .B2(n_15272),
    .Y(n_66830));
 AOI22xp5_ASAP7_75t_SL g213865 (.A1(n_66817),
    .A2(n_6732),
    .B1(n_211),
    .B2(n_32335),
    .Y(n_66831));
 AOI22xp5_ASAP7_75t_SL g213866 (.A1(n_29790),
    .A2(n_66817),
    .B1(\u4_mem[0] [10]),
    .B2(n_33657),
    .Y(n_66832));
 AOI22xp5_ASAP7_75t_SL g213867 (.A1(n_66817),
    .A2(n_43537),
    .B1(\u7_mem[1] [10]),
    .B2(n_50220),
    .Y(n_66833));
 AOI22xp5_ASAP7_75t_SL g213868 (.A1(n_66824),
    .A2(n_67247),
    .B1(n_396),
    .B2(n_29621),
    .Y(n_66834));
 AOI22xp5_ASAP7_75t_SL g213869 (.A1(n_52893),
    .A2(n_66817),
    .B1(\u3_mem[0] [10]),
    .B2(n_51288),
    .Y(n_66835));
 AOI22xp33_ASAP7_75t_SL g214227 (.A1(n_67246),
    .A2(n_67247),
    .B1(oc2_cfg[6]),
    .B2(n_67248),
    .Y(n_67249));
 INVx3_ASAP7_75t_SL g214228 (.A(n_10276),
    .Y(n_67246));
 INVx5_ASAP7_75t_SL g214229 (.A(n_9555),
    .Y(n_67247));
 BUFx6f_ASAP7_75t_SL g214230 (.A(n_29619),
    .Y(n_67248));
 NAND2xp5_ASAP7_75t_SL g214470 (.A(n_13995),
    .B(n_67546),
    .Y(n_67490));
 AOI22xp5_ASAP7_75t_SL g214503 (.A1(n_79178),
    .A2(\u8_mem[2] [13]),
    .B1(\u8_mem[0] [13]),
    .B2(n_70885),
    .Y(n_67546));
 INVx4_ASAP7_75t_SL g214942 (.A(n_9967),
    .Y(n_68207));
 AOI22xp5_ASAP7_75t_SL g214943 (.A1(n_68207),
    .A2(n_78410),
    .B1(n_31741),
    .B2(\u6_mem[1] [4]),
    .Y(n_68211));
 AOI22xp5_ASAP7_75t_SL g214944 (.A1(n_68207),
    .A2(n_64818),
    .B1(\u8_mem[3] [4]),
    .B2(n_70622),
    .Y(n_68212));
 AOI22xp5_ASAP7_75t_SL g214946 (.A1(n_68207),
    .A2(n_12403),
    .B1(\u7_mem[0] [4]),
    .B2(n_3386),
    .Y(n_68215));
 AOI22xp5_ASAP7_75t_SL g214948 (.A1(\u8_mem[1] [4]),
    .A2(n_31464),
    .B1(n_68207),
    .B2(n_75734),
    .Y(n_68217));
 AOI22xp5_ASAP7_75t_SL g214950 (.A1(n_24806),
    .A2(n_68207),
    .B1(\u3_mem[2] [4]),
    .B2(n_13295),
    .Y(n_68219));
 AOI22xp5_ASAP7_75t_SL g214952 (.A1(n_68207),
    .A2(n_43535),
    .B1(\u7_mem[1] [4]),
    .B2(n_50220),
    .Y(n_68221));
 AOI22xp5_ASAP7_75t_SL g214954 (.A1(n_68207),
    .A2(n_6732),
    .B1(n_307),
    .B2(n_32335),
    .Y(n_68223));
 AOI21xp5_ASAP7_75t_SL g214958 (.A1(n_16797),
    .A2(n_68207),
    .B(n_2644),
    .Y(n_68227));
 AOI22xp5_ASAP7_75t_SL g214960 (.A1(n_11128),
    .A2(n_68207),
    .B1(\u5_mem[3] [4]),
    .B2(n_9476),
    .Y(n_68229));
 AOI22xp5_ASAP7_75t_SL g214962 (.A1(n_52893),
    .A2(n_68207),
    .B1(\u3_mem[0] [4]),
    .B2(n_51296),
    .Y(n_68231));
 AOI22xp5_ASAP7_75t_SL g215495 (.A1(n_69010),
    .A2(n_3461),
    .B1(\u8_mem[0] [4]),
    .B2(n_3460),
    .Y(n_69011));
 AOI22xp5_ASAP7_75t_SL g215497 (.A1(crac_out[4]),
    .A2(n_28367),
    .B1(n_69010),
    .B2(n_17579),
    .Y(n_69012));
 AOI22xp5_ASAP7_75t_SL g215498 (.A1(\u6_mem[3] [4]),
    .A2(n_77233),
    .B1(n_69010),
    .B2(n_61228),
    .Y(n_69013));
 AOI22xp5_ASAP7_75t_SL g215499 (.A1(n_3320),
    .A2(n_69010),
    .B1(\u8_mem[2] [4]),
    .B2(n_16900),
    .Y(n_69014));
 AOI22xp5_ASAP7_75t_SL g215500 (.A1(n_29790),
    .A2(n_69010),
    .B1(\u4_mem[0] [4]),
    .B2(n_33655),
    .Y(n_69015));
 AOI22xp5_ASAP7_75t_SL g215501 (.A1(n_3188),
    .A2(n_69010),
    .B1(\u7_mem[2] [4]),
    .B2(n_13325),
    .Y(n_69016));
 AOI22xp5_ASAP7_75t_SL g215502 (.A1(n_69010),
    .A2(n_21311),
    .B1(n_230),
    .B2(n_26541),
    .Y(n_69017));
 AOI22xp5_ASAP7_75t_SL g215503 (.A1(n_3420),
    .A2(n_69010),
    .B1(\u6_mem[0] [4]),
    .B2(n_3425),
    .Y(n_69018));
 AOI22xp5_ASAP7_75t_SL g215504 (.A1(n_26385),
    .A2(n_69010),
    .B1(\u5_mem[0] [4]),
    .B2(n_26389),
    .Y(n_69019));
 AOI22xp5_ASAP7_75t_SL g215505 (.A1(n_69010),
    .A2(n_32164),
    .B1(\u5_mem[1] [4]),
    .B2(n_13500),
    .Y(n_69020));
 AOI22xp5_ASAP7_75t_SL g215506 (.A1(n_3285),
    .A2(n_69010),
    .B1(\u5_mem[2] [4]),
    .B2(n_43020),
    .Y(n_69021));
 AOI22xp5_ASAP7_75t_SL g215507 (.A1(n_69010),
    .A2(n_30253),
    .B1(\u4_mem[3] [4]),
    .B2(n_35908),
    .Y(n_69022));
 AOI22xp5_ASAP7_75t_SL g215508 (.A1(n_24633),
    .A2(n_69010),
    .B1(\u4_mem[2] [4]),
    .B2(n_13312),
    .Y(n_69023));
 AOI22xp5_ASAP7_75t_SL g215509 (.A1(n_69010),
    .A2(n_48107),
    .B1(\u4_mem[1] [4]),
    .B2(n_65763),
    .Y(n_69024));
 AOI22xp33_ASAP7_75t_SL g215510 (.A1(n_69025),
    .A2(n_14570),
    .B1(\u7_mem[3] [4]),
    .B2(n_33772),
    .Y(n_69026));
 AOI22xp33_ASAP7_75t_SL g215511 (.A1(n_69025),
    .A2(n_21527),
    .B1(\u3_mem[3] [4]),
    .B2(n_21550),
    .Y(n_69027));
 AOI22xp33_ASAP7_75t_SL g215512 (.A1(n_22577),
    .A2(\u3_mem[1] [4]),
    .B1(n_69025),
    .B2(n_16009),
    .Y(n_69028));
 AOI22xp5_ASAP7_75t_SL g215513 (.A1(n_69010),
    .A2(n_67247),
    .B1(n_18899),
    .B2(n_67248),
    .Y(n_69029));
 INVx3_ASAP7_75t_SL g216235 (.A(n_24750),
    .Y(n_69795));
 NAND2x1p5_ASAP7_75t_SL g216236 (.A(u6_wp[0]),
    .B(o7_we),
    .Y(n_69796));
 AOI22xp5_ASAP7_75t_SL g216448 (.A1(\u6_mem[2] [4]),
    .A2(n_70039),
    .B1(n_68207),
    .B2(n_78043),
    .Y(n_70040));
 INVx4_ASAP7_75t_SL g216449 (.A(n_70038),
    .Y(n_70039));
 AND3x4_ASAP7_75t_SL g216450 (.A(n_24750),
    .B(n_20669),
    .C(o7_we),
    .Y(n_70038));
 AOI22xp5_ASAP7_75t_SL g216451 (.A1(\u6_mem[2] [18]),
    .A2(n_78042),
    .B1(n_10194),
    .B2(n_78043),
    .Y(n_70042));
 AOI22xp5_ASAP7_75t_SL g216453 (.A1(\u6_mem[2] [14]),
    .A2(n_78042),
    .B1(n_28251),
    .B2(n_78043),
    .Y(n_70043));
 AOI22xp5_ASAP7_75t_SL g216454 (.A1(\u6_mem[2] [23]),
    .A2(n_78042),
    .B1(n_65930),
    .B2(n_78043),
    .Y(n_70044));
 AOI22xp5_ASAP7_75t_SL g216455 (.A1(\u6_mem[2] [28]),
    .A2(n_78042),
    .B1(n_65920),
    .B2(n_78043),
    .Y(n_70045));
 AOI22xp5_ASAP7_75t_SL g216456 (.A1(\u6_mem[2] [5]),
    .A2(n_78042),
    .B1(n_66869),
    .B2(n_78043),
    .Y(n_70046));
 AOI22xp5_ASAP7_75t_SL g216457 (.A1(n_78043),
    .A2(n_65908),
    .B1(\u6_mem[2] [27]),
    .B2(n_78042),
    .Y(n_70047));
 AOI22xp5_ASAP7_75t_SL g216458 (.A1(n_78043),
    .A2(n_65925),
    .B1(\u6_mem[2] [25]),
    .B2(n_78042),
    .Y(n_70048));
 AOI22xp5_ASAP7_75t_SL g216460 (.A1(n_78043),
    .A2(n_10638),
    .B1(\u6_mem[2] [30]),
    .B2(n_78042),
    .Y(n_70050));
 AOI22xp5_ASAP7_75t_SL g216461 (.A1(\u6_mem[2] [21]),
    .A2(n_78042),
    .B1(n_32916),
    .B2(n_78043),
    .Y(n_70051));
 AOI22xp5_ASAP7_75t_SL g216462 (.A1(\u6_mem[2] [24]),
    .A2(n_78042),
    .B1(n_65914),
    .B2(n_78043),
    .Y(n_70052));
 AOI22xp5_ASAP7_75t_SL g216463 (.A1(\u6_mem[2] [20]),
    .A2(n_78042),
    .B1(n_33024),
    .B2(n_78043),
    .Y(n_70053));
 AOI22xp5_ASAP7_75t_SL g216464 (.A1(\u6_mem[2] [15]),
    .A2(n_78042),
    .B1(n_28913),
    .B2(n_78043),
    .Y(n_70054));
 AOI22xp5_ASAP7_75t_SL g216465 (.A1(\u6_mem[2] [19]),
    .A2(n_78042),
    .B1(n_10196),
    .B2(n_78043),
    .Y(n_70055));
 AOI22xp5_ASAP7_75t_SL g216466 (.A1(\u6_mem[2] [0]),
    .A2(n_78042),
    .B1(n_10924),
    .B2(n_78043),
    .Y(n_70056));
 AOI22xp5_ASAP7_75t_SL g216467 (.A1(\u6_mem[2] [10]),
    .A2(n_70039),
    .B1(n_66817),
    .B2(n_78043),
    .Y(n_70057));
 AOI22xp5_ASAP7_75t_SL g216468 (.A1(\u6_mem[2] [2]),
    .A2(n_70039),
    .B1(n_66000),
    .B2(n_78043),
    .Y(n_70058));
 AOI22xp5_ASAP7_75t_SL g216469 (.A1(\u6_mem[2] [8]),
    .A2(n_70039),
    .B1(n_65980),
    .B2(n_78043),
    .Y(n_70059));
 AOI22xp5_ASAP7_75t_SL g216470 (.A1(\u6_mem[2] [16]),
    .A2(n_70039),
    .B1(n_28276),
    .B2(n_78043),
    .Y(n_70060));
 AOI22xp5_ASAP7_75t_SL g216471 (.A1(\u6_mem[2] [9]),
    .A2(n_70039),
    .B1(n_79972),
    .B2(n_78043),
    .Y(n_70061));
 AOI22xp5_ASAP7_75t_SL g216472 (.A1(\u6_mem[2] [3]),
    .A2(n_70039),
    .B1(n_15867),
    .B2(n_78043),
    .Y(n_70062));
 AOI22xp5_ASAP7_75t_SL g216473 (.A1(\u6_mem[2] [29]),
    .A2(n_70039),
    .B1(n_15952),
    .B2(n_78043),
    .Y(n_70063));
 AOI22xp5_ASAP7_75t_SL g216474 (.A1(\u6_mem[2] [26]),
    .A2(n_70039),
    .B1(n_35437),
    .B2(n_78043),
    .Y(n_70064));
 AOI22xp5_ASAP7_75t_SL g216475 (.A1(\u6_mem[2] [6]),
    .A2(n_70039),
    .B1(n_66004),
    .B2(n_78043),
    .Y(n_70065));
 AOI22xp5_ASAP7_75t_SL g216476 (.A1(n_78043),
    .A2(n_10026),
    .B1(\u6_mem[2] [12]),
    .B2(n_70039),
    .Y(n_70066));
 AOI22xp5_ASAP7_75t_SL g216477 (.A1(n_78043),
    .A2(n_15920),
    .B1(\u6_mem[2] [31]),
    .B2(n_70039),
    .Y(n_70067));
 AOI22xp5_ASAP7_75t_SL g216478 (.A1(\u6_mem[2] [13]),
    .A2(n_70039),
    .B1(n_35041),
    .B2(n_78043),
    .Y(n_70068));
 AOI22xp5_ASAP7_75t_SL g216479 (.A1(\u6_mem[2] [7]),
    .A2(n_70039),
    .B1(n_17578),
    .B2(n_78043),
    .Y(n_70069));
 AOI22xp5_ASAP7_75t_SL g216480 (.A1(\u6_mem[2] [11]),
    .A2(n_70039),
    .B1(n_66843),
    .B2(n_78043),
    .Y(n_70070));
 AOI22xp5_ASAP7_75t_SL g216481 (.A1(\u6_mem[2] [17]),
    .A2(n_70039),
    .B1(n_65952),
    .B2(n_78043),
    .Y(n_70071));
 AOI22xp5_ASAP7_75t_SL g216482 (.A1(\u6_mem[2] [22]),
    .A2(n_70039),
    .B1(n_67246),
    .B2(n_78043),
    .Y(n_70072));
 NAND2xp5_ASAP7_75t_SL g216619 (.A(n_70240),
    .B(n_56854),
    .Y(n_70241));
 AOI22xp5_ASAP7_75t_SL g216620 (.A1(\u5_mem[1] [15]),
    .A2(n_64833),
    .B1(\u5_mem[0] [15]),
    .B2(n_65642),
    .Y(n_70240));
 NOR2x1_ASAP7_75t_SL g216674 (.A(n_70323),
    .B(n_70322),
    .Y(n_70324));
 INVx4_ASAP7_75t_SL g216675 (.A(n_36068),
    .Y(n_70322));
 NAND3xp33_ASAP7_75t_L g216676 (.A(n_33644),
    .B(out_slt0[7]),
    .C(oc4_cfg[0]),
    .Y(n_70323));
 NAND2xp5_ASAP7_75t_SL g216677 (.A(out_slt0[7]),
    .B(n_33644),
    .Y(n_70325));
 INVx2_ASAP7_75t_SL g216678 (.A(oc4_cfg[0]),
    .Y(n_70326));
 NAND2xp5_ASAP7_75t_SL g216707 (.A(n_78041),
    .B(n_70413),
    .Y(n_70414));
 NAND2xp5_ASAP7_75t_SL g216708 (.A(n_70411),
    .B(n_78942),
    .Y(n_70413));
 AOI22xp33_ASAP7_75t_SL g216709 (.A1(n_77853),
    .A2(\u6_mem[2] [17]),
    .B1(n_41152),
    .B2(\u6_mem[3] [17]),
    .Y(n_70411));
 INVx1_ASAP7_75t_SL g216711 (.A(n_70413),
    .Y(n_70415));
 OR2x6_ASAP7_75t_SL g216872 (.A(n_64192),
    .B(n_70621),
    .Y(n_70622));
 INVx2_ASAP7_75t_SL g216873 (.A(n_64814),
    .Y(n_70621));
 AND2x2_ASAP7_75t_SL g216898 (.A(n_4028),
    .B(n_70648),
    .Y(n_70649));
 NOR3x1_ASAP7_75t_SL g216899 (.A(n_34538),
    .B(n_43082),
    .C(n_19133),
    .Y(n_70648));
 NAND2x1_ASAP7_75t_SL g217132 (.A(n_70886),
    .B(n_13982),
    .Y(n_70887));
 AOI22xp5_ASAP7_75t_SL g217133 (.A1(n_79178),
    .A2(\u8_mem[2] [12]),
    .B1(n_70885),
    .B2(\u8_mem[0] [12]),
    .Y(n_70886));
 NAND2xp5_ASAP7_75t_SL g217531 (.A(n_71350),
    .B(n_71351),
    .Y(n_71352));
 INVx2_ASAP7_75t_SL g217560 (.A(u4_rp[0]),
    .Y(n_71390));
 XOR2xp5_ASAP7_75t_SL g217561 (.A(n_50810),
    .B(n_12275),
    .Y(n_71391));
 BUFx2_ASAP7_75t_L g217562 (.A(u4_rp[0]),
    .Y(n_71392));
 INVx1_ASAP7_75t_SL g217563 (.A(n_71391),
    .Y(n_71393));
 AOI21xp33_ASAP7_75t_SL g217564 (.A1(n_36008),
    .A2(n_7766),
    .B(n_71394),
    .Y(n_71395));
 AOI22xp33_ASAP7_75t_SL g217565 (.A1(n_71390),
    .A2(n_71391),
    .B1(n_71393),
    .B2(n_71392),
    .Y(n_71394));
 AND2x2_ASAP7_75t_SL g218106 (.A(u3_rp[1]),
    .B(n_33784),
    .Y(n_71971));
 AND2x6_ASAP7_75t_SL g218107 (.A(u3_rp[1]),
    .B(u3_rp[2]),
    .Y(n_71972));
 NAND2xp5_ASAP7_75t_SL g218108 (.A(n_20756),
    .B(n_71973),
    .Y(n_71974));
 AOI22xp33_ASAP7_75t_SL g218109 (.A1(n_71971),
    .A2(\u3_mem[1] [19]),
    .B1(n_71972),
    .B2(\u3_mem[3] [19]),
    .Y(n_71973));
 INVx2_ASAP7_75t_SL g218176 (.A(u8_rp[2]),
    .Y(n_72057));
 HB1xp67_ASAP7_75t_SL g218178 (.A(n_72058),
    .Y(n_72059));
 XOR2xp5_ASAP7_75t_L g218180 (.A(n_78135),
    .B(n_72058),
    .Y(n_72060));
 AO21x1_ASAP7_75t_L g218181 (.A1(n_16853),
    .A2(n_21190),
    .B(n_72059),
    .Y(n_72062));
 NAND3xp33_ASAP7_75t_L g218182 (.A(n_16853),
    .B(n_72059),
    .C(n_21190),
    .Y(n_72063));
 OA21x2_ASAP7_75t_SL g218183 (.A1(n_72058),
    .A2(n_14765),
    .B(n_72064),
    .Y(n_72065));
 NAND2x1_ASAP7_75t_SL g218184 (.A(n_64817),
    .B(n_72058),
    .Y(n_72064));
 AOI21xp33_ASAP7_75t_SL g218198 (.A1(n_72083),
    .A2(n_72084),
    .B(n_78167),
    .Y(n_72087));
 AOI221xp5_ASAP7_75t_SL g218313 (.A1(n_72307),
    .A2(n_5028),
    .B1(n_4988),
    .B2(out_slt9[19]),
    .C(n_4340),
    .Y(n_72308));
 NAND4xp25_ASAP7_75t_SL g218314 (.A(n_79197),
    .B(n_43667),
    .C(n_43666),
    .D(n_43665),
    .Y(n_72307));
 AOI31xp33_ASAP7_75t_SL g218860 (.A1(n_72908),
    .A2(n_556),
    .A3(u8_wp[2]),
    .B(n_2744),
    .Y(n_72909));
 OR2x2_ASAP7_75t_SL g218861 (.A(n_70621),
    .B(n_64192),
    .Y(n_72908));
 NAND2x1_ASAP7_75t_SL g219093 (.A(n_78954),
    .B(n_12106),
    .Y(n_73154));
 NAND2xp5_ASAP7_75t_SL g219102 (.A(n_49203),
    .B(n_643),
    .Y(n_73169));
 AOI21xp5_ASAP7_75t_SL g219103 (.A1(n_73173),
    .A2(n_79104),
    .B(n_38382),
    .Y(n_73174));
 NAND4xp25_ASAP7_75t_SL g219104 (.A(n_73170),
    .B(n_73169),
    .C(n_73171),
    .D(n_73172),
    .Y(n_73173));
 AOI22xp33_ASAP7_75t_SL g219105 (.A1(\u5_mem[0] [30]),
    .A2(n_64793),
    .B1(\u5_mem[1] [30]),
    .B2(n_6071),
    .Y(n_73170));
 NAND2xp33_ASAP7_75t_L g219106 (.A(n_65001),
    .B(n_37200),
    .Y(n_73171));
 AOI22xp33_ASAP7_75t_R g219107 (.A1(\u5_mem[2] [30]),
    .A2(n_1459),
    .B1(\u5_mem[3] [30]),
    .B2(n_56865),
    .Y(n_73172));
 AND2x4_ASAP7_75t_SL g219108 (.A(n_49618),
    .B(n_53365),
    .Y(n_73175));
 OAI21xp5_ASAP7_75t_SL g219109 (.A1(n_59252),
    .A2(n_65029),
    .B(n_73176),
    .Y(n_73177));
 NAND2xp5_ASAP7_75t_SL g219110 (.A(n_73175),
    .B(\u7_mem[3] [20]),
    .Y(n_73176));
 OA21x2_ASAP7_75t_SL g219218 (.A1(n_70322),
    .A2(n_21341),
    .B(n_47740),
    .Y(n_73300));
 BUFx6f_ASAP7_75t_SL g219220 (.A(n_73300),
    .Y(n_73301));
 NAND2xp5_ASAP7_75t_SL g219222 (.A(n_73301),
    .B(out_slt9[8]),
    .Y(n_73304));
 AND2x2_ASAP7_75t_R g219224 (.A(out_slt9[17]),
    .B(n_73301),
    .Y(n_73306));
 HB1xp67_ASAP7_75t_SL g219226 (.A(n_73301),
    .Y(n_73307));
 AND2x2_ASAP7_75t_R g219230 (.A(out_slt9[16]),
    .B(n_73301),
    .Y(n_73312));
 HB1xp67_ASAP7_75t_R g219231 (.A(n_73301),
    .Y(n_73313));
 AOI22xp5_ASAP7_75t_SL g219293 (.A1(n_79971),
    .A2(n_75734),
    .B1(\u8_mem[1] [9]),
    .B2(n_75735),
    .Y(n_73388));
 AOI22xp5_ASAP7_75t_SL g219306 (.A1(\u8_mem[1] [18]),
    .A2(n_73399),
    .B1(n_10171),
    .B2(n_73997),
    .Y(n_73400));
 INVx4_ASAP7_75t_SL g219307 (.A(n_26501),
    .Y(n_73399));
 AOI22xp5_ASAP7_75t_SL g219876 (.A1(n_73996),
    .A2(n_73997),
    .B1(\u8_mem[1] [21]),
    .B2(n_75735),
    .Y(n_73999));
 INVx3_ASAP7_75t_SL g219877 (.A(n_66017),
    .Y(n_73996));
 AND2x4_ASAP7_75t_SL g219878 (.A(n_14763),
    .B(n_40978),
    .Y(n_73997));
 AND2x6_ASAP7_75t_SL g22 (.A(n_24801),
    .B(n_33604),
    .Y(n_24803));
 AOI22xp5_ASAP7_75t_SL g221581 (.A1(n_75733),
    .A2(n_75734),
    .B1(\u8_mem[1] [0]),
    .B2(n_75735),
    .Y(n_75736));
 BUFx6f_ASAP7_75t_SL g221582 (.A(wb_din[0]),
    .Y(n_75733));
 AND2x4_ASAP7_75t_SL g221583 (.A(n_14763),
    .B(n_40978),
    .Y(n_75734));
 INVx4_ASAP7_75t_SL g221584 (.A(n_26501),
    .Y(n_75735));
 NAND3xp33_ASAP7_75t_SL g221642 (.A(n_75792),
    .B(n_75793),
    .C(n_75794),
    .Y(n_75795));
 XNOR2xp5_ASAP7_75t_SL g221643 (.A(u3_wp[2]),
    .B(n_21793),
    .Y(n_75792));
 AOI21xp33_ASAP7_75t_L g221644 (.A1(n_20317),
    .A2(n_2454),
    .B(n_20319),
    .Y(n_75793));
 INVxp67_ASAP7_75t_SL g221645 (.A(n_2162),
    .Y(n_75794));
 NAND2xp5_ASAP7_75t_SL g221872 (.A(n_76054),
    .B(n_76055),
    .Y(n_76056));
 INVx2_ASAP7_75t_SL g221873 (.A(ac97_rst_force),
    .Y(n_76054));
 INVx1_ASAP7_75t_SL g221874 (.A(n_42613),
    .Y(n_76055));
 AOI22xp5_ASAP7_75t_SL g222523 (.A1(\u6_mem[1] [4]),
    .A2(n_76763),
    .B1(\u6_mem[3] [4]),
    .B2(n_41152),
    .Y(n_76764));
 AND2x6_ASAP7_75t_SL g222524 (.A(u6_rp[1]),
    .B(n_78938),
    .Y(n_76763));
 AOI22xp5_ASAP7_75t_SL g222537 (.A1(\u6_mem[3] [2]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_66000),
    .Y(n_76778));
 AOI22xp5_ASAP7_75t_SL g222740 (.A1(\u6_mem[3] [6]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_32644),
    .Y(n_76986));
 AOI22xp5_ASAP7_75t_SL g222985 (.A1(\u6_mem[3] [12]),
    .A2(n_77233),
    .B1(n_61228),
    .B2(n_65997),
    .Y(n_77234));
 OR2x6_ASAP7_75t_SL g222986 (.A(n_69796),
    .B(n_69795),
    .Y(n_77233));
 AOI22xp5_ASAP7_75t_SL g223 (.A1(n_49625),
    .A2(n_24735),
    .B1(\u9_mem[3] [18]),
    .B2(n_45330),
    .Y(n_49626));
 AOI22xp5_ASAP7_75t_SL g223141 (.A1(\u3_mem[2] [30]),
    .A2(n_77396),
    .B1(\u3_mem[3] [30]),
    .B2(n_22062),
    .Y(n_77397));
 INVxp33_ASAP7_75t_SL g223142 (.A(n_1783),
    .Y(n_77396));
 INVx2_ASAP7_75t_SL g223143 (.A(n_1783),
    .Y(n_77398));
 OAI22xp5_ASAP7_75t_SL g223449 (.A1(n_18964),
    .A2(n_18739),
    .B1(u6_wp[0]),
    .B2(n_77796),
    .Y(n_77797));
 INVx3_ASAP7_75t_SL g223450 (.A(n_18739),
    .Y(n_77796));
 AND2x6_ASAP7_75t_SL g223484 (.A(u6_rp[2]),
    .B(n_78937),
    .Y(n_77853));
 AND2x2_ASAP7_75t_SL g223485 (.A(n_48404),
    .B(n_78941),
    .Y(n_77855));
 AO21x1_ASAP7_75t_SL g223535 (.A1(n_48404),
    .A2(n_78941),
    .B(n_21076),
    .Y(n_77964));
 AOI22xp5_ASAP7_75t_SL g223555 (.A1(\u8_mem[1] [6]),
    .A2(n_78274),
    .B1(\u8_mem[3] [6]),
    .B2(n_78273),
    .Y(n_78002));
 AO21x1_ASAP7_75t_SL g223595 (.A1(n_48423),
    .A2(n_78946),
    .B(n_21076),
    .Y(n_78040));
 INVx6_ASAP7_75t_SL g223596 (.A(n_21076),
    .Y(n_78041));
 AOI22xp33_ASAP7_75t_SL g223597 (.A1(\u6_mem[2] [1]),
    .A2(n_78042),
    .B1(n_78043),
    .B2(n_78044),
    .Y(n_78045));
 INVx4_ASAP7_75t_SL g223598 (.A(n_70038),
    .Y(n_78042));
 AND3x4_ASAP7_75t_SL g223599 (.A(n_20671),
    .B(n_24750),
    .C(o7_we),
    .Y(n_78043));
 INVx2_ASAP7_75t_SL g223600 (.A(n_10890),
    .Y(n_78044));
 BUFx3_ASAP7_75t_SL g223648 (.A(oc2_cfg[0]),
    .Y(n_78094));
 NOR2xp33_ASAP7_75t_R g223681 (.A(n_78931),
    .B(n_78932),
    .Y(n_78134));
 AND2x2_ASAP7_75t_SL g223683 (.A(n_78932),
    .B(u8_rp[0]),
    .Y(n_78135));
 A2O1A1Ixp33_ASAP7_75t_SL g223687 (.A1(n_36528),
    .A2(n_78137),
    .B(n_78138),
    .C(n_15007),
    .Y(n_78139));
 NOR2xp33_ASAP7_75t_L g223688 (.A(n_78932),
    .B(n_57084),
    .Y(n_78138));
 NAND2xp33_ASAP7_75t_R g223689 (.A(n_73300),
    .B(n_78137),
    .Y(n_78140));
 NOR4xp25_ASAP7_75t_SL g223712 (.A(n_245),
    .B(n_78166),
    .C(n_20673),
    .D(n_24741),
    .Y(n_78167));
 NAND2xp5_ASAP7_75t_SL g223713 (.A(n_78164),
    .B(n_57964),
    .Y(n_78166));
 INVx1_ASAP7_75t_SL g223714 (.A(u6_wp[2]),
    .Y(n_78164));
 INVx1_ASAP7_75t_SL g223715 (.A(n_50109),
    .Y(n_57964));
 AND2x6_ASAP7_75t_SL g223809 (.A(u8_rp[2]),
    .B(u8_rp[1]),
    .Y(n_78273));
 AND2x6_ASAP7_75t_SL g223810 (.A(u8_rp[1]),
    .B(n_7888),
    .Y(n_78274));
 NAND2xp5_ASAP7_75t_SL g223811 (.A(n_79179),
    .B(n_78275),
    .Y(n_78276));
 AOI22xp5_ASAP7_75t_SL g223812 (.A1(\u8_mem[3] [14]),
    .A2(n_78273),
    .B1(n_78274),
    .B2(\u8_mem[1] [14]),
    .Y(n_78275));
 AOI22xp5_ASAP7_75t_SL g223942 (.A1(n_65925),
    .A2(n_78410),
    .B1(n_22396),
    .B2(\u6_mem[1] [25]),
    .Y(n_78411));
 AND3x4_ASAP7_75t_SL g223943 (.A(n_18966),
    .B(n_29352),
    .C(o7_we),
    .Y(n_78410));
 OAI22xp5_ASAP7_75t_SL g224 (.A1(n_50458),
    .A2(n_1678),
    .B1(n_48056),
    .B2(n_48648),
    .Y(n_49625));
 AOI22xp5_ASAP7_75t_SL g224146 (.A1(\u10_mem[1] [5]),
    .A2(n_78621),
    .B1(n_24803),
    .B2(n_50553),
    .Y(n_78622));
 OR2x6_ASAP7_75t_SL g224147 (.A(n_32299),
    .B(n_32300),
    .Y(n_78621));
 AOI22xp33_ASAP7_75t_SL g224208 (.A1(\u6_mem[0] [25]),
    .A2(n_79305),
    .B1(\u6_mem[2] [25]),
    .B2(n_79306),
    .Y(n_78683));
 NAND2xp5_ASAP7_75t_L g224209 (.A(n_73154),
    .B(n_78810),
    .Y(n_78684));
 NAND2xp5_ASAP7_75t_SL g224210 (.A(n_31107),
    .B(n_78041),
    .Y(n_78685));
 AOI22xp33_ASAP7_75t_L g224211 (.A1(\u6_mem[1] [25]),
    .A2(n_48415),
    .B1(\u6_mem[3] [25]),
    .B2(n_17704),
    .Y(n_78686));
 AND2x4_ASAP7_75t_SL g224333 (.A(n_678),
    .B(n_21076),
    .Y(n_78810));
 NAND4xp25_ASAP7_75t_SL g224335 (.A(n_2113),
    .B(n_79327),
    .C(n_1430),
    .D(n_1406),
    .Y(n_78813));
 INVx4_ASAP7_75t_SL g224453 (.A(u8_wp[0]),
    .Y(n_78931));
 AOI31xp33_ASAP7_75t_SL g224455 (.A1(n_72065),
    .A2(n_78933),
    .A3(n_43075),
    .B(oc5_int_set[2]),
    .Y(n_78934));
 AOI22xp5_ASAP7_75t_SL g224456 (.A1(u8_wp[0]),
    .A2(n_78930),
    .B1(n_78932),
    .B2(n_78931),
    .Y(n_78933));
 OAI22xp33_ASAP7_75t_L g224457 (.A1(n_78935),
    .A2(u8_rp[0]),
    .B1(n_497),
    .B2(n_78933),
    .Y(n_78936));
 INVx1_ASAP7_75t_SL g224458 (.A(n_78933),
    .Y(n_78935));
 AOI22xp5_ASAP7_75t_SL g224461 (.A1(n_78939),
    .A2(\u6_mem[0] [8]),
    .B1(n_76763),
    .B2(\u6_mem[1] [8]),
    .Y(n_78940));
 AND2x6_ASAP7_75t_SL g224462 (.A(n_78938),
    .B(n_78937),
    .Y(n_78939));
 AOI22xp5_ASAP7_75t_SL g224463 (.A1(\u6_mem[0] [18]),
    .A2(n_78939),
    .B1(n_77853),
    .B2(\u6_mem[2] [18]),
    .Y(n_78941));
 AOI22xp5_ASAP7_75t_SL g224464 (.A1(n_78939),
    .A2(\u6_mem[0] [17]),
    .B1(\u6_mem[1] [17]),
    .B2(n_76763),
    .Y(n_78942));
 AOI22xp5_ASAP7_75t_SL g224465 (.A1(n_78939),
    .A2(\u6_mem[0] [10]),
    .B1(\u6_mem[1] [10]),
    .B2(n_76763),
    .Y(n_78943));
 AOI22xp5_ASAP7_75t_SL g224466 (.A1(\u6_mem[0] [5]),
    .A2(n_78939),
    .B1(n_77853),
    .B2(\u6_mem[2] [5]),
    .Y(n_78944));
 AOI22xp5_ASAP7_75t_SL g224467 (.A1(n_78939),
    .A2(\u6_mem[0] [12]),
    .B1(\u6_mem[2] [12]),
    .B2(n_77853),
    .Y(n_78945));
 AOI22xp5_ASAP7_75t_SL g224468 (.A1(\u6_mem[0] [19]),
    .A2(n_78939),
    .B1(n_77853),
    .B2(\u6_mem[2] [19]),
    .Y(n_78946));
 AOI22xp5_ASAP7_75t_SL g224469 (.A1(\u6_mem[0] [6]),
    .A2(n_78939),
    .B1(n_77853),
    .B2(\u6_mem[2] [6]),
    .Y(n_78947));
 AOI22xp5_ASAP7_75t_SL g224470 (.A1(\u6_mem[0] [7]),
    .A2(n_78939),
    .B1(\u6_mem[2] [7]),
    .B2(n_77853),
    .Y(n_78948));
 AOI22xp5_ASAP7_75t_SL g224471 (.A1(n_78939),
    .A2(\u6_mem[0] [11]),
    .B1(n_76763),
    .B2(\u6_mem[1] [11]),
    .Y(n_78949));
 AOI22xp5_ASAP7_75t_SL g224472 (.A1(n_78939),
    .A2(\u6_mem[0] [15]),
    .B1(n_76763),
    .B2(\u6_mem[1] [15]),
    .Y(n_78950));
 AOI22xp5_ASAP7_75t_SL g224473 (.A1(\u6_mem[0] [2]),
    .A2(n_78939),
    .B1(\u6_mem[1] [2]),
    .B2(n_76763),
    .Y(n_78951));
 AOI22xp5_ASAP7_75t_SL g224474 (.A1(n_78939),
    .A2(\u6_mem[0] [1]),
    .B1(\u6_mem[1] [1]),
    .B2(n_76763),
    .Y(n_78952));
 AOI22xp5_ASAP7_75t_SL g224475 (.A1(n_78939),
    .A2(\u6_mem[0] [0]),
    .B1(n_76763),
    .B2(\u6_mem[1] [0]),
    .Y(n_78953));
 AOI22xp5_ASAP7_75t_SL g224476 (.A1(n_76763),
    .A2(\u6_mem[1] [9]),
    .B1(n_78939),
    .B2(\u6_mem[0] [9]),
    .Y(n_78954));
 AOI22xp5_ASAP7_75t_SL g224477 (.A1(n_78939),
    .A2(\u6_mem[0] [14]),
    .B1(\u6_mem[1] [14]),
    .B2(n_76763),
    .Y(n_78955));
 AOI22xp5_ASAP7_75t_SL g224478 (.A1(\u6_mem[0] [13]),
    .A2(n_78939),
    .B1(n_76763),
    .B2(\u6_mem[1] [13]),
    .Y(n_78956));
 AOI22xp5_ASAP7_75t_SL g224479 (.A1(\u6_mem[0] [3]),
    .A2(n_78939),
    .B1(n_76763),
    .B2(\u6_mem[1] [3]),
    .Y(n_78957));
 AOI22xp33_ASAP7_75t_SL g224480 (.A1(n_78939),
    .A2(\u6_mem[0] [16]),
    .B1(n_76763),
    .B2(\u6_mem[1] [16]),
    .Y(n_78958));
 AOI22xp33_ASAP7_75t_SL g224481 (.A1(n_78939),
    .A2(\u6_mem[0] [4]),
    .B1(n_77853),
    .B2(\u6_mem[2] [4]),
    .Y(n_78959));
 NAND2xp5_ASAP7_75t_SL g224522 (.A(n_36068),
    .B(n_78094),
    .Y(n_79016));
 INVx1_ASAP7_75t_SL g224523 (.A(n_34472),
    .Y(n_79017));
 NAND3xp33_ASAP7_75t_SL g224524 (.A(n_34472),
    .B(n_78094),
    .C(n_36068),
    .Y(n_79019));
 AND2x4_ASAP7_75t_SL g224572 (.A(n_34473),
    .B(n_79103),
    .Y(n_79104));
 NOR2x1_ASAP7_75t_SL g224573 (.A(n_79017),
    .B(n_79016),
    .Y(n_79103));
 AOI221xp5_ASAP7_75t_SL g224630 (.A1(n_79167),
    .A2(n_25956),
    .B1(n_5062),
    .B2(out_slt7[13]),
    .C(n_4425),
    .Y(n_79168));
 NAND4xp25_ASAP7_75t_SL g224631 (.A(n_78684),
    .B(n_78683),
    .C(n_78686),
    .D(n_78685),
    .Y(n_79167));
 XOR2xp5_ASAP7_75t_SL g224638 (.A(n_79175),
    .B(n_13990),
    .Y(n_79176));
 XOR2xp5_ASAP7_75t_L g224639 (.A(u8_wp[2]),
    .B(u8_rp[3]),
    .Y(n_79175));
 XNOR2xp5_ASAP7_75t_SL g224640 (.A(u8_rp[3]),
    .B(n_13990),
    .Y(n_79177));
 AOI22xp33_ASAP7_75t_SL g224641 (.A1(n_79178),
    .A2(\u8_mem[2] [14]),
    .B1(\u8_mem[0] [14]),
    .B2(n_59474),
    .Y(n_79179));
 AND2x6_ASAP7_75t_SL g224642 (.A(u8_rp[2]),
    .B(n_53264),
    .Y(n_79178));
 INVx2_ASAP7_75t_SL g224651 (.A(n_79192),
    .Y(n_79193));
 BUFx2_ASAP7_75t_SL g224652 (.A(n_253),
    .Y(n_79192));
 NOR3xp33_ASAP7_75t_SL g224653 (.A(n_477),
    .B(n_79194),
    .C(n_4119),
    .Y(n_79195));
 BUFx2_ASAP7_75t_SL g224654 (.A(n_79192),
    .Y(n_79194));
 NOR2xp33_ASAP7_75t_SL g224655 (.A(n_79194),
    .B(n_4119),
    .Y(n_79196));
 AO21x1_ASAP7_75t_SL g224656 (.A1(n_51496),
    .A2(n_13988),
    .B(n_79194),
    .Y(n_79197));
 INVx2_ASAP7_75t_SL g224658 (.A(n_79193),
    .Y(n_79198));
 INVx2_ASAP7_75t_SL g224662 (.A(n_79194),
    .Y(n_79203));
 NAND2xp5_ASAP7_75t_SL g224663 (.A(n_79198),
    .B(n_15007),
    .Y(n_79204));
 AND2x2_ASAP7_75t_SL g224664 (.A(n_79198),
    .B(n_15007),
    .Y(n_79205));
 INVxp67_ASAP7_75t_R g224665 (.A(n_79198),
    .Y(n_79206));
 OAI211xp5_ASAP7_75t_SL g224666 (.A1(n_79198),
    .A2(n_4341),
    .B(n_1435),
    .C(n_2236),
    .Y(n_79207));
 OAI222xp33_ASAP7_75t_SL g224667 (.A1(n_2440),
    .A2(n_23655),
    .B1(n_17617),
    .B2(n_79198),
    .C1(n_25928),
    .C2(n_57084),
    .Y(n_79208));
 AND3x2_ASAP7_75t_SL g224740 (.A(n_7712),
    .B(n_18739),
    .C(n_37337),
    .Y(n_79305));
 AND2x4_ASAP7_75t_SL g224741 (.A(n_37337),
    .B(n_77853),
    .Y(n_79306));
 NAND4xp25_ASAP7_75t_SL g224742 (.A(n_16749),
    .B(n_16751),
    .C(n_79307),
    .D(n_16750),
    .Y(n_79308));
 AOI22xp33_ASAP7_75t_SL g224743 (.A1(\u6_mem[0] [24]),
    .A2(n_79305),
    .B1(n_79306),
    .B2(\u6_mem[2] [24]),
    .Y(n_79307));
 NAND2x1_ASAP7_75t_SL g224755 (.A(n_48413),
    .B(n_78948),
    .Y(n_79326));
 HB1xp67_ASAP7_75t_SL g23 (.A(n_78938),
    .Y(n_7712));
 AOI31xp33_ASAP7_75t_SL g233 (.A1(n_58734),
    .A2(n_71391),
    .A3(n_2696),
    .B(oc1_int_set[2]),
    .Y(n_58735));
 OAI22xp5_ASAP7_75t_SL g234 (.A1(n_48110),
    .A2(n_42779),
    .B1(n_23526),
    .B2(n_48106),
    .Y(n_58734));
 AOI22xp5_ASAP7_75t_SL g2349 (.A1(n_7486),
    .A2(n_38758),
    .B1(n_25405),
    .B2(n_14792),
    .Y(n_7491));
 NAND3xp33_ASAP7_75t_SL g2351 (.A(n_4381),
    .B(n_16672),
    .C(n_13955),
    .Y(n_7486));
 INVx4_ASAP7_75t_SL g24 (.A(wb_addr_i[4]),
    .Y(n_8296));
 AOI21xp5_ASAP7_75t_SL g244 (.A1(n_26710),
    .A2(n_26712),
    .B(n_26713),
    .Y(n_26714));
 NOR2xp33_ASAP7_75t_R g245 (.A(n_26711),
    .B(n_18857),
    .Y(n_26712));
 INVxp67_ASAP7_75t_SL g248 (.A(n_4280),
    .Y(n_26710));
 NAND2x1p5_ASAP7_75t_SL g25 (.A(n_8262),
    .B(n_21331),
    .Y(n_21332));
 NAND4xp25_ASAP7_75t_SL g253 (.A(n_1401),
    .B(n_1421),
    .C(n_2092),
    .D(n_77964),
    .Y(n_14448));
 INVxp33_ASAP7_75t_R g26 (.A(n_31534),
    .Y(n_31396));
 AOI22xp33_ASAP7_75t_SL g263 (.A1(n_29006),
    .A2(n_26553),
    .B1(n_20594),
    .B2(\u11_mem[3] [7]),
    .Y(n_7500));
 AOI22xp33_ASAP7_75t_SL g264 (.A1(n_26553),
    .A2(n_28953),
    .B1(n_20593),
    .B2(\u11_mem[1] [7]),
    .Y(n_7501));
 NOR2xp33_ASAP7_75t_SL g265 (.A(n_34524),
    .B(n_34525),
    .Y(n_34526));
 O2A1O1Ixp33_ASAP7_75t_SL g266 (.A1(i4_status[0]),
    .A2(ic1_cfg[4]),
    .B(i4_status[1]),
    .C(ic1_cfg[5]),
    .Y(n_34525));
 OAI31xp33_ASAP7_75t_SL g267 (.A1(ic1_cfg[4]),
    .A2(i4_status[1]),
    .A3(i4_status[0]),
    .B(n_2228),
    .Y(n_34524));
 INVx2_ASAP7_75t_SL g27 (.A(n_50293),
    .Y(n_52768));
 OAI21xp5_ASAP7_75t_SL g273 (.A1(n_59639),
    .A2(n_4320),
    .B(n_65646),
    .Y(n_7641));
 NOR2xp33_ASAP7_75t_SL g275 (.A(n_72081),
    .B(n_72082),
    .Y(n_72083));
 OR2x2_ASAP7_75t_SL g276 (.A(n_69796),
    .B(n_69795),
    .Y(n_72084));
 INVxp33_ASAP7_75t_SL g278 (.A(n_179),
    .Y(n_72082));
 INVxp33_ASAP7_75t_SL g279 (.A(u6_wp[2]),
    .Y(n_72081));
 INVxp33_ASAP7_75t_R g28 (.A(n_8334),
    .Y(n_8336));
 NOR2xp67_ASAP7_75t_SL g291 (.A(n_31795),
    .B(n_31747),
    .Y(n_29874));
 NOR2xp33_ASAP7_75t_R g3 (.A(n_14763),
    .B(n_40978),
    .Y(n_17545));
 NOR2xp33_ASAP7_75t_R g30 (.A(n_33100),
    .B(n_503),
    .Y(n_23504));
 INVx2_ASAP7_75t_SL g300 (.A(u14_u2_en_out_l2),
    .Y(n_31581));
 AND2x2_ASAP7_75t_L g309 (.A(out_slt4[5]),
    .B(n_43087),
    .Y(n_51464));
 INVx1_ASAP7_75t_R g31 (.A(n_8234),
    .Y(n_8236));
 AOI222xp33_ASAP7_75t_SL g310 (.A1(n_78810),
    .A2(n_34190),
    .B1(n_79305),
    .B2(\u6_mem[0] [28]),
    .C1(n_79306),
    .C2(\u6_mem[2] [28]),
    .Y(n_7569));
 AO22x1_ASAP7_75t_SL g311 (.A1(\u7_mem[1] [29]),
    .A2(n_65056),
    .B1(\u7_mem[0] [29]),
    .B2(n_65055),
    .Y(n_64745));
 NAND2x1_ASAP7_75t_SL g312 (.A(n_56056),
    .B(n_56057),
    .Y(n_64744));
 NAND2xp5_ASAP7_75t_SL g32 (.A(n_37200),
    .B(n_70241),
    .Y(n_31870));
 XNOR2xp5_ASAP7_75t_SL g329 (.A(n_78134),
    .B(n_72065),
    .Y(n_58150));
 NAND2xp5_ASAP7_75t_SL g33 (.A(n_70241),
    .B(n_643),
    .Y(n_31871));
 INVxp67_ASAP7_75t_SL g34 (.A(n_27004),
    .Y(n_13594));
 INVx1_ASAP7_75t_R g35 (.A(n_66003),
    .Y(n_66005));
 INVxp33_ASAP7_75t_R g36 (.A(\u3_mem[1] [21]),
    .Y(n_24509));
 AOI22xp5_ASAP7_75t_SL g37 (.A1(\u3_mem[3] [0]),
    .A2(n_71972),
    .B1(n_50388),
    .B2(\u3_mem[2] [0]),
    .Y(n_21231));
 INVx1_ASAP7_75t_SL g38 (.A(in_slt3[6]),
    .Y(n_48056));
 NOR3xp33_ASAP7_75t_R g39 (.A(n_117),
    .B(u14_u8_full_empty_r),
    .C(n_4075),
    .Y(n_13599));
 HB1xp67_ASAP7_75t_L g4 (.A(n_65971),
    .Y(n_65972));
 NAND3xp33_ASAP7_75t_SL g40 (.A(n_43720),
    .B(n_65058),
    .C(n_2503),
    .Y(n_43721));
 AOI22xp33_ASAP7_75t_SL g41 (.A1(n_60873),
    .A2(\u9_mem[1] [11]),
    .B1(n_24734),
    .B2(n_15693),
    .Y(n_22694));
 INVx1_ASAP7_75t_SL g42 (.A(n_21225),
    .Y(n_13598));
 NAND3xp33_ASAP7_75t_SL g426 (.A(n_8252),
    .B(n_28674),
    .C(n_10620),
    .Y(n_8255));
 AOI22xp5_ASAP7_75t_R g429 (.A1(n_8235),
    .A2(i3_dout[5]),
    .B1(n_14933),
    .B2(i6_dout[5]),
    .Y(n_8252));
 NAND3xp33_ASAP7_75t_SL g43 (.A(n_7691),
    .B(n_7692),
    .C(n_7693),
    .Y(n_7694));
 NAND3xp33_ASAP7_75t_SL g433 (.A(n_43169),
    .B(n_43170),
    .C(n_43171),
    .Y(n_43172));
 AOI222xp33_ASAP7_75t_SL g434 (.A1(n_8173),
    .A2(i4_dout[19]),
    .B1(i3_dout[19]),
    .B2(n_8235),
    .C1(i6_dout[19]),
    .C2(n_8338),
    .Y(n_43171));
 AOI21xp33_ASAP7_75t_SL g435 (.A1(u13_ints_r[19]),
    .A2(n_10614),
    .B(n_10869),
    .Y(n_43170));
 AOI22xp5_ASAP7_75t_SL g436 (.A1(n_7083),
    .A2(n_291),
    .B1(n_6961),
    .B2(n_512),
    .Y(n_43169));
 AOI211xp5_ASAP7_75t_SL g439 (.A1(n_28103),
    .A2(n_25405),
    .B(n_7524),
    .C(n_4383),
    .Y(n_14418));
 NOR2x1_ASAP7_75t_L g44 (.A(n_1701),
    .B(n_10937),
    .Y(n_30483));
 NAND3xp33_ASAP7_75t_SL g448 (.A(n_8248),
    .B(n_22928),
    .C(n_10627),
    .Y(n_8251));
 INVx1_ASAP7_75t_SL g45 (.A(ic2_cfg[3]),
    .Y(n_7693));
 AOI22xp5_ASAP7_75t_R g451 (.A1(n_8235),
    .A2(i3_dout[13]),
    .B1(n_8338),
    .B2(i6_dout[13]),
    .Y(n_8248));
 AOI211xp5_ASAP7_75t_SL g455 (.A1(n_52933),
    .A2(n_32582),
    .B(n_4546),
    .C(n_51464),
    .Y(n_52934));
 OAI222xp33_ASAP7_75t_SL g456 (.A1(n_23671),
    .A2(n_26801),
    .B1(n_17712),
    .B2(n_36007),
    .C1(n_17711),
    .C2(n_8113),
    .Y(n_52933));
 INVx1_ASAP7_75t_SL g46 (.A(u14_u8_en_out_l2),
    .Y(n_7695));
 AND2x2_ASAP7_75t_L g463 (.A(out_slt4[6]),
    .B(n_43087),
    .Y(n_7426));
 INVx1_ASAP7_75t_SL g47 (.A(ic2_cfg[2]),
    .Y(n_7692));
 AOI211x1_ASAP7_75t_SL g471 (.A1(n_54564),
    .A2(n_79104),
    .B(n_66662),
    .C(n_38379),
    .Y(n_54566));
 OAI222xp33_ASAP7_75t_SL g472 (.A1(n_16781),
    .A2(n_59644),
    .B1(n_59639),
    .B2(n_31733),
    .C1(n_43206),
    .C2(n_27013),
    .Y(n_54564));
 INVxp67_ASAP7_75t_R g48 (.A(u11_wp[0]),
    .Y(n_7691));
 NAND4xp25_ASAP7_75t_SL g486 (.A(n_22025),
    .B(n_28692),
    .C(n_22027),
    .D(n_22028),
    .Y(n_22029));
 AOI222xp33_ASAP7_75t_SL g487 (.A1(n_8173),
    .A2(i4_dout[18]),
    .B1(i6_dout[18]),
    .B2(n_8338),
    .C1(i3_dout[18]),
    .C2(n_8235),
    .Y(n_22028));
 NAND2xp5_ASAP7_75t_L g489 (.A(n_10614),
    .B(n_2048),
    .Y(n_22027));
 AOI22xp5_ASAP7_75t_SL g49 (.A1(n_71972),
    .A2(\u3_mem[3] [14]),
    .B1(n_50342),
    .B2(\u3_mem[2] [14]),
    .Y(n_31849));
 NAND3xp33_ASAP7_75t_SL g490 (.A(n_16741),
    .B(n_35469),
    .C(n_16742),
    .Y(n_16743));
 AOI22xp33_ASAP7_75t_L g492 (.A1(\u4_mem[1] [23]),
    .A2(n_1765),
    .B1(\u4_mem[0] [23]),
    .B2(n_1766),
    .Y(n_16741));
 AOI22xp33_ASAP7_75t_R g493 (.A1(\u4_mem[3] [23]),
    .A2(n_23531),
    .B1(n_17624),
    .B2(\u4_mem[2] [23]),
    .Y(n_16742));
 INVx2_ASAP7_75t_SL g5 (.A(n_8339),
    .Y(n_8340));
 AOI22xp33_ASAP7_75t_SL g50 (.A1(\u5_mem[1] [18]),
    .A2(n_64833),
    .B1(\u5_mem[3] [18]),
    .B2(n_56842),
    .Y(n_64834));
 OAI21xp5_ASAP7_75t_SL g501 (.A1(n_70198),
    .A2(n_70199),
    .B(n_70200),
    .Y(n_70201));
 O2A1O1Ixp33_ASAP7_75t_SL g502 (.A1(o9_status[0]),
    .A2(oc5_cfg[4]),
    .B(o9_status[1]),
    .C(oc5_cfg[5]),
    .Y(n_70199));
 OAI31xp33_ASAP7_75t_SL g503 (.A1(oc5_cfg[4]),
    .A2(o9_status[1]),
    .A3(o9_status[0]),
    .B(n_2964),
    .Y(n_70198));
 NOR3xp33_ASAP7_75t_SL g504 (.A(n_47739),
    .B(n_1381),
    .C(dma_ack_i[5]),
    .Y(n_70200));
 INVx2_ASAP7_75t_SL g51 (.A(n_66015),
    .Y(n_66017));
 AOI221xp5_ASAP7_75t_SL g519 (.A1(n_36361),
    .A2(out_slt7[6]),
    .B1(n_37344),
    .B2(n_25954),
    .C(n_4413),
    .Y(n_29970));
 NAND2x1p5_ASAP7_75t_SL g52 (.A(u3_rp[1]),
    .B(n_33784),
    .Y(n_7567));
 AOI22xp33_ASAP7_75t_SL g53 (.A1(n_30253),
    .A2(n_10683),
    .B1(n_35911),
    .B2(\u4_mem[3] [29]),
    .Y(n_30247));
 INVx8_ASAP7_75t_SL g54 (.A(n_35910),
    .Y(n_30253));
 NOR5xp2_ASAP7_75t_R g549 (.A(n_19009),
    .B(n_24725),
    .C(n_47541),
    .D(n_50088),
    .E(n_303),
    .Y(n_14947));
 NAND2x1_ASAP7_75t_SL g55 (.A(wb_addr_i[3]),
    .B(wb_addr_i[2]),
    .Y(n_8183));
 NAND2x1_ASAP7_75t_SL g56 (.A(wb_addr_i[3]),
    .B(wb_addr_i[2]),
    .Y(n_8189));
 NAND4xp25_ASAP7_75t_SL g57 (.A(n_445),
    .B(n_47794),
    .C(n_363),
    .D(n_452),
    .Y(n_14226));
 NOR2xp33_ASAP7_75t_SL g58 (.A(n_1760),
    .B(n_1972),
    .Y(n_49319));
 OAI211xp5_ASAP7_75t_SL g583 (.A1(n_65000),
    .A2(n_2596),
    .B(n_1452),
    .C(n_16739),
    .Y(n_7941));
 INVxp33_ASAP7_75t_R g586 (.A(out_slt6[15]),
    .Y(n_7270));
 INVx2_ASAP7_75t_L g59 (.A(n_8186),
    .Y(n_375));
 AND2x2_ASAP7_75t_SL g6 (.A(n_8315),
    .B(n_8232),
    .Y(n_8339));
 INVx2_ASAP7_75t_SL g60 (.A(ic0_cfg[0]),
    .Y(n_8186));
 AOI221xp5_ASAP7_75t_SL g606 (.A1(u13_intm_r[13]),
    .A2(n_7082),
    .B1(n_8174),
    .B2(i4_dout[13]),
    .C(n_22927),
    .Y(n_22928));
 OAI22xp5_ASAP7_75t_SL g607 (.A1(n_18903),
    .A2(n_28669),
    .B1(n_14909),
    .B2(n_47),
    .Y(n_22927));
 XNOR2xp5_ASAP7_75t_SL g61 (.A(u6_rp[3]),
    .B(n_12067),
    .Y(n_13898));
 NAND4xp25_ASAP7_75t_SL g62 (.A(n_2191),
    .B(n_8123),
    .C(n_1801),
    .D(n_1751),
    .Y(n_8124));
 NAND2xp5_ASAP7_75t_L g63 (.A(n_425),
    .B(n_31850),
    .Y(n_8123));
 NAND2xp5_ASAP7_75t_SL g64 (.A(n_47551),
    .B(n_31850),
    .Y(n_8128));
 XNOR2x1_ASAP7_75t_SL g66 (.B(n_56857),
    .Y(n_37311),
    .A(u5_rp[3]));
 INVxp67_ASAP7_75t_SL g67 (.A(n_41378),
    .Y(n_64014));
 INVx1_ASAP7_75t_R g676 (.A(n_78810),
    .Y(n_7442));
 NAND2xp5_ASAP7_75t_SL g678 (.A(out_slt4[15]),
    .B(n_7781),
    .Y(n_14924));
 AND2x4_ASAP7_75t_SL g69 (.A(n_24316),
    .B(n_33774),
    .Y(n_14570));
 OAI211xp5_ASAP7_75t_SL g692 (.A1(n_4324),
    .A2(n_842),
    .B(n_1955),
    .C(n_66667),
    .Y(n_7597));
 AND2x2_ASAP7_75t_SL g7 (.A(n_8232),
    .B(n_8315),
    .Y(n_8341));
 INVx1_ASAP7_75t_SL g70 (.A(n_31272),
    .Y(n_31273));
 INVx3_ASAP7_75t_SL g71 (.A(n_10486),
    .Y(n_65908));
 INVx2_ASAP7_75t_SL g72 (.A(n_65906),
    .Y(n_10486));
 AOI211xp5_ASAP7_75t_SL g73 (.A1(n_59643),
    .A2(n_79104),
    .B(n_38378),
    .C(n_66676),
    .Y(n_7308));
 NAND4xp25_ASAP7_75t_SL g75 (.A(n_15080),
    .B(n_36256),
    .C(n_1802),
    .D(n_46485),
    .Y(n_46486));
 OAI211xp5_ASAP7_75t_SL g756 (.A1(n_5706),
    .A2(n_842),
    .B(n_64711),
    .C(n_66680),
    .Y(n_7430));
 AOI21xp5_ASAP7_75t_SL g76 (.A1(n_7994),
    .A2(n_28696),
    .B(n_38381),
    .Y(n_7995));
 OAI211xp5_ASAP7_75t_SL g77 (.A1(n_59639),
    .A2(n_27013),
    .B(n_2486),
    .C(n_2149),
    .Y(n_7994));
 NOR2x1_ASAP7_75t_SL g78 (.A(wb_addr_i[6]),
    .B(wb_addr_i[5]),
    .Y(n_8220));
 AO21x1_ASAP7_75t_L g79 (.A1(n_1863),
    .A2(n_7414),
    .B(n_2523),
    .Y(n_14791));
 AND2x4_ASAP7_75t_SL g8 (.A(n_35632),
    .B(n_36008),
    .Y(n_17624));
 NAND2xp33_ASAP7_75t_SL g80 (.A(n_425),
    .B(n_47552),
    .Y(n_14789));
 NAND2xp5_ASAP7_75t_SL g81 (.A(n_47551),
    .B(n_43320),
    .Y(n_14788));
 AOI22xp5_ASAP7_75t_SL g82 (.A1(crac_out[12]),
    .A2(n_28367),
    .B1(n_65997),
    .B2(n_17579),
    .Y(n_17525));
 AOI22xp5_ASAP7_75t_SL g83 (.A1(\u3_mem[2] [13]),
    .A2(n_7562),
    .B1(\u3_mem[0] [13]),
    .B2(n_50341),
    .Y(n_7563));
 INVxp67_ASAP7_75t_SL g84 (.A(n_43320),
    .Y(n_14794));
 AOI22xp5_ASAP7_75t_SL g85 (.A1(crac_out[6]),
    .A2(n_28367),
    .B1(n_66004),
    .B2(n_17579),
    .Y(n_17528));
 OAI22xp33_ASAP7_75t_SL g86 (.A1(n_12098),
    .A2(n_12062),
    .B1(n_2693),
    .B2(n_3999),
    .Y(n_28110));
 AOI22xp5_ASAP7_75t_SL g87 (.A1(\u5_mem[1] [19]),
    .A2(n_64833),
    .B1(\u5_mem[0] [19]),
    .B2(n_65642),
    .Y(n_42030));
 AOI22xp5_ASAP7_75t_SL g88 (.A1(n_65920),
    .A2(n_64819),
    .B1(\u8_mem[3] [28]),
    .B2(n_72908),
    .Y(n_47157));
 AOI22xp5_ASAP7_75t_SL g89 (.A1(n_28424),
    .A2(n_73997),
    .B1(\u8_mem[1] [24]),
    .B2(n_31460),
    .Y(n_15927));
 AND2x4_ASAP7_75t_SL g8_dup217131 (.A(n_72057),
    .B(n_78930),
    .Y(n_70885));
 INVx1_ASAP7_75t_SL g9 (.A(u14_u0_en_out_l2),
    .Y(n_19132));
 AOI22xp5_ASAP7_75t_SL g90 (.A1(n_45625),
    .A2(n_45624),
    .B1(\u11_mem[2] [19]),
    .B2(n_61785),
    .Y(n_45627));
 OAI21xp5_ASAP7_75t_SL g91 (.A1(n_35474),
    .A2(n_31535),
    .B(n_36662),
    .Y(n_35476));
 AOI221xp5_ASAP7_75t_SL g92 (.A1(oc4_cfg[1]),
    .A2(n_11006),
    .B1(i6_dout[1]),
    .B2(n_8338),
    .C(n_2118),
    .Y(n_8242));
 O2A1O1Ixp5_ASAP7_75t_SL g93 (.A1(n_8012),
    .A2(n_26904),
    .B(n_4976),
    .C(n_38380),
    .Y(n_8013));
 OAI21xp33_ASAP7_75t_SL g94 (.A1(n_7665),
    .A2(n_59639),
    .B(n_64713),
    .Y(n_8012));
 OAI22xp33_ASAP7_75t_SL g95 (.A1(n_273),
    .A2(n_27320),
    .B1(n_27315),
    .B2(n_26428),
    .Y(n_27321));
 NOR2x1p5_ASAP7_75t_SL g96 (.A(wb_addr_i[4]),
    .B(wb_addr_i[2]),
    .Y(n_8238));
 AOI21xp5_ASAP7_75t_SL g97 (.A1(n_31464),
    .A2(\u8_mem[1] [3]),
    .B(n_19378),
    .Y(n_15869));
 INVxp67_ASAP7_75t_L g98 (.A(n_7672),
    .Y(n_43206));
 AOI21xp5_ASAP7_75t_SL g99 (.A1(\u3_mem[1] [0]),
    .A2(n_22505),
    .B(n_15495),
    .Y(n_15496));
 DFFHQNx1_ASAP7_75t_R \in_valid_s1_reg[0]  (.CLK(clk_i),
    .D(n_2442),
    .QN(in_valid_s1[0]));
 DFFHQNx1_ASAP7_75t_R \in_valid_s1_reg[1]  (.CLK(clk_i),
    .D(n_2222),
    .QN(in_valid_s1[1]));
 DFFHQNx1_ASAP7_75t_R \in_valid_s1_reg[2]  (.CLK(clk_i),
    .D(n_2271),
    .QN(in_valid_s1[2]));
 DFFHQNx1_ASAP7_75t_SL \in_valid_s_reg[0]  (.CLK(clk_i),
    .D(n_20821),
    .QN(in_valid_s[0]));
 DFFHQNx1_ASAP7_75t_SL \in_valid_s_reg[1]  (.CLK(clk_i),
    .D(n_2557),
    .QN(in_valid_s[1]));
 DFFHQNx1_ASAP7_75t_SL \in_valid_s_reg[2]  (.CLK(clk_i),
    .D(n_18928),
    .QN(in_valid_s[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5517),
    .QN(u0_slt0_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5528),
    .QN(u0_slt0_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5530),
    .QN(u0_slt0_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5533),
    .QN(u0_slt0_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5534),
    .QN(u0_slt0_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5536),
    .QN(u0_slt0_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5537),
    .QN(u0_slt0_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5518),
    .QN(u0_slt0_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5519),
    .QN(u0_slt0_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5520),
    .QN(u0_slt0_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5521),
    .QN(u0_slt0_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5523),
    .QN(u0_slt0_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5524),
    .QN(u0_slt0_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5525),
    .QN(u0_slt0_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5526),
    .QN(u0_slt0_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt0_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5527),
    .QN(u0_slt0_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5497),
    .QN(u0_slt1_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5507),
    .QN(u0_slt1_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5508),
    .QN(u0_slt1_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5509),
    .QN(u0_slt1_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5510),
    .QN(u0_slt1_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5511),
    .QN(u0_slt1_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5512),
    .QN(u0_slt1_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5513),
    .QN(u0_slt1_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5514),
    .QN(u0_slt1_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5515),
    .QN(u0_slt1_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5516),
    .QN(u0_slt1_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5498),
    .QN(u0_slt1_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5499),
    .QN(u0_slt1_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5500),
    .QN(u0_slt1_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5501),
    .QN(u0_slt1_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5502),
    .QN(u0_slt1_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5503),
    .QN(u0_slt1_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5504),
    .QN(u0_slt1_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5505),
    .QN(u0_slt1_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt1_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5506),
    .QN(u0_slt1_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5477),
    .QN(u0_slt2_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5487),
    .QN(u0_slt2_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5488),
    .QN(u0_slt2_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5489),
    .QN(u0_slt2_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5490),
    .QN(u0_slt2_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5491),
    .QN(u0_slt2_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5492),
    .QN(u0_slt2_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5493),
    .QN(u0_slt2_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5494),
    .QN(u0_slt2_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5495),
    .QN(u0_slt2_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5496),
    .QN(u0_slt2_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5478),
    .QN(u0_slt2_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5479),
    .QN(u0_slt2_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5480),
    .QN(u0_slt2_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5481),
    .QN(u0_slt2_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5482),
    .QN(u0_slt2_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5483),
    .QN(u0_slt2_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5484),
    .QN(u0_slt2_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5485),
    .QN(u0_slt2_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt2_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5486),
    .QN(u0_slt2_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5457),
    .QN(u0_slt3_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5467),
    .QN(u0_slt3_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5468),
    .QN(u0_slt3_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5469),
    .QN(u0_slt3_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5470),
    .QN(u0_slt3_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5471),
    .QN(u0_slt3_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5472),
    .QN(u0_slt3_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5473),
    .QN(u0_slt3_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5474),
    .QN(u0_slt3_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5475),
    .QN(u0_slt3_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5476),
    .QN(u0_slt3_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5458),
    .QN(u0_slt3_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5459),
    .QN(u0_slt3_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5460),
    .QN(u0_slt3_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5461),
    .QN(u0_slt3_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5462),
    .QN(u0_slt3_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5463),
    .QN(u0_slt3_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5464),
    .QN(u0_slt3_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5465),
    .QN(u0_slt3_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt3_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5466),
    .QN(u0_slt3_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5437),
    .QN(u0_slt4_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5447),
    .QN(u0_slt4_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5448),
    .QN(u0_slt4_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5449),
    .QN(u0_slt4_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5450),
    .QN(u0_slt4_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5451),
    .QN(u0_slt4_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5452),
    .QN(u0_slt4_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5453),
    .QN(u0_slt4_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5454),
    .QN(u0_slt4_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5455),
    .QN(u0_slt4_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5456),
    .QN(u0_slt4_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5438),
    .QN(u0_slt4_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5439),
    .QN(u0_slt4_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5440),
    .QN(u0_slt4_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5441),
    .QN(u0_slt4_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5442),
    .QN(u0_slt4_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5443),
    .QN(u0_slt4_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5444),
    .QN(u0_slt4_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5445),
    .QN(u0_slt4_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt4_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5446),
    .QN(u0_slt4_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5417),
    .QN(u0_slt5_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5427),
    .QN(u0_slt5_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5428),
    .QN(u0_slt5_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5429),
    .QN(u0_slt5_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5430),
    .QN(u0_slt5_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5431),
    .QN(u0_slt5_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5432),
    .QN(u0_slt5_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5433),
    .QN(u0_slt5_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5434),
    .QN(u0_slt5_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5435),
    .QN(u0_slt5_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5436),
    .QN(u0_slt5_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5418),
    .QN(u0_slt5_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5419),
    .QN(u0_slt5_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5420),
    .QN(u0_slt5_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5421),
    .QN(u0_slt5_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5422),
    .QN(u0_slt5_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5423),
    .QN(u0_slt5_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5424),
    .QN(u0_slt5_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5425),
    .QN(u0_slt5_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt5_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5426),
    .QN(u0_slt5_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5397),
    .QN(u0_slt6_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5407),
    .QN(u0_slt6_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5408),
    .QN(u0_slt6_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5409),
    .QN(u0_slt6_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5410),
    .QN(u0_slt6_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5411),
    .QN(u0_slt6_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5412),
    .QN(u0_slt6_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5413),
    .QN(u0_slt6_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5414),
    .QN(u0_slt6_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5415),
    .QN(u0_slt6_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5416),
    .QN(u0_slt6_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5398),
    .QN(u0_slt6_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5399),
    .QN(u0_slt6_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5400),
    .QN(u0_slt6_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5401),
    .QN(u0_slt6_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5402),
    .QN(u0_slt6_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5403),
    .QN(u0_slt6_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5404),
    .QN(u0_slt6_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5405),
    .QN(u0_slt6_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt6_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5406),
    .QN(u0_slt6_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5377),
    .QN(u0_slt7_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5387),
    .QN(u0_slt7_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5388),
    .QN(u0_slt7_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5389),
    .QN(u0_slt7_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5390),
    .QN(u0_slt7_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5391),
    .QN(u0_slt7_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5392),
    .QN(u0_slt7_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5393),
    .QN(u0_slt7_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5394),
    .QN(u0_slt7_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5395),
    .QN(u0_slt7_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5396),
    .QN(u0_slt7_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5378),
    .QN(u0_slt7_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5379),
    .QN(u0_slt7_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5380),
    .QN(u0_slt7_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5381),
    .QN(u0_slt7_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5382),
    .QN(u0_slt7_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5383),
    .QN(u0_slt7_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5384),
    .QN(u0_slt7_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5385),
    .QN(u0_slt7_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt7_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5386),
    .QN(u0_slt7_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_5357),
    .QN(u0_slt8_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5367),
    .QN(u0_slt8_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5368),
    .QN(u0_slt8_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5369),
    .QN(u0_slt8_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5370),
    .QN(u0_slt8_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5371),
    .QN(u0_slt8_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5372),
    .QN(u0_slt8_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5373),
    .QN(u0_slt8_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5374),
    .QN(u0_slt8_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5375),
    .QN(u0_slt8_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5376),
    .QN(u0_slt8_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_5358),
    .QN(u0_slt8_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_5359),
    .QN(u0_slt8_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_5360),
    .QN(u0_slt8_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5361),
    .QN(u0_slt8_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5362),
    .QN(u0_slt8_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5363),
    .QN(u0_slt8_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5364),
    .QN(u0_slt8_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5365),
    .QN(u0_slt8_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt8_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5366),
    .QN(u0_slt8_r[9]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2277),
    .QN(u0_slt9_r[0]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5332),
    .QN(u0_slt9_r[10]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5348),
    .QN(u0_slt9_r[11]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5349),
    .QN(u0_slt9_r[12]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5350),
    .QN(u0_slt9_r[13]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5351),
    .QN(u0_slt9_r[14]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5352),
    .QN(u0_slt9_r[15]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5353),
    .QN(u0_slt9_r[16]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5354),
    .QN(u0_slt9_r[17]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5355),
    .QN(u0_slt9_r[18]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5356),
    .QN(u0_slt9_r[19]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_2741),
    .QN(u0_slt9_r[1]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_3985),
    .QN(u0_slt9_r[2]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_4487),
    .QN(u0_slt9_r[3]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_5266),
    .QN(u0_slt9_r[4]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_5279),
    .QN(u0_slt9_r[5]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_5293),
    .QN(u0_slt9_r[6]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5303),
    .QN(u0_slt9_r[7]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5314),
    .QN(u0_slt9_r[8]));
 DFFHQNx1_ASAP7_75t_R \u0_slt9_r_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5325),
    .QN(u0_slt9_r[9]));
 DFFHQNx1_ASAP7_75t_SL \u10_din_tmp1_reg[0]  (.CLK(clk_i),
    .D(n_34614),
    .QN(u10_din_tmp1[0]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[10]  (.CLK(clk_i),
    .D(n_29885),
    .QN(u10_din_tmp1[10]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[11]  (.CLK(clk_i),
    .D(n_34413),
    .QN(u10_din_tmp1[11]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[12]  (.CLK(clk_i),
    .D(n_34378),
    .QN(u10_din_tmp1[12]));
 DFFHQNx1_ASAP7_75t_SL \u10_din_tmp1_reg[13]  (.CLK(clk_i),
    .D(n_29899),
    .QN(u10_din_tmp1[13]));
 DFFHQNx1_ASAP7_75t_SL \u10_din_tmp1_reg[14]  (.CLK(clk_i),
    .D(n_29909),
    .QN(u10_din_tmp1[14]));
 DFFHQNx1_ASAP7_75t_SL \u10_din_tmp1_reg[15]  (.CLK(clk_i),
    .D(n_29907),
    .QN(u10_din_tmp1[15]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[1]  (.CLK(clk_i),
    .D(n_29889),
    .QN(u10_din_tmp1[1]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[2]  (.CLK(clk_i),
    .D(n_29905),
    .QN(u10_din_tmp1[2]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[3]  (.CLK(clk_i),
    .D(n_29915),
    .QN(u10_din_tmp1[3]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[4]  (.CLK(clk_i),
    .D(n_29891),
    .QN(u10_din_tmp1[4]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[5]  (.CLK(clk_i),
    .D(n_29897),
    .QN(u10_din_tmp1[5]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[6]  (.CLK(clk_i),
    .D(n_34422),
    .QN(u10_din_tmp1[6]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[7]  (.CLK(clk_i),
    .D(n_29911),
    .QN(u10_din_tmp1[7]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[8]  (.CLK(clk_i),
    .D(n_34363),
    .QN(u10_din_tmp1[8]));
 DFFHQNx2_ASAP7_75t_SL \u10_din_tmp1_reg[9]  (.CLK(clk_i),
    .D(n_29903),
    .QN(u10_din_tmp1[9]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[0]  (.CLK(clk_i),
    .D(n_1598),
    .Q(i4_dout[0]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[10]  (.CLK(clk_i),
    .D(n_1552),
    .Q(i4_dout[10]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[11]  (.CLK(clk_i),
    .D(n_1597),
    .Q(i4_dout[11]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[12]  (.CLK(clk_i),
    .D(n_1596),
    .Q(i4_dout[12]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[13]  (.CLK(clk_i),
    .D(n_1545),
    .Q(i4_dout[13]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[14]  (.CLK(clk_i),
    .D(n_1595),
    .Q(i4_dout[14]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[15]  (.CLK(clk_i),
    .D(n_1590),
    .Q(i4_dout[15]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[16]  (.CLK(clk_i),
    .D(n_1588),
    .Q(i4_dout[16]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[17]  (.CLK(clk_i),
    .D(n_1519),
    .Q(i4_dout[17]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[18]  (.CLK(clk_i),
    .D(n_1637),
    .Q(i4_dout[18]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[19]  (.CLK(clk_i),
    .D(n_1546),
    .Q(i4_dout[19]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[1]  (.CLK(clk_i),
    .D(n_1599),
    .Q(i4_dout[1]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[20]  (.CLK(clk_i),
    .D(n_1560),
    .Q(i4_dout[20]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[21]  (.CLK(clk_i),
    .D(n_1549),
    .Q(i4_dout[21]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[22]  (.CLK(clk_i),
    .D(n_1573),
    .Q(i4_dout[22]));
 DFFHQNx2_ASAP7_75t_SL \u10_dout_reg[23]  (.CLK(clk_i),
    .D(n_29874),
    .QN(i4_dout[23]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[24]  (.CLK(clk_i),
    .D(n_1587),
    .Q(i4_dout[24]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[25]  (.CLK(clk_i),
    .D(n_1593),
    .Q(i4_dout[25]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[26]  (.CLK(clk_i),
    .D(n_1631),
    .Q(i4_dout[26]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[27]  (.CLK(clk_i),
    .D(n_1592),
    .Q(i4_dout[27]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[28]  (.CLK(clk_i),
    .D(n_1591),
    .Q(i4_dout[28]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[29]  (.CLK(clk_i),
    .D(n_1586),
    .Q(i4_dout[29]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[2]  (.CLK(clk_i),
    .D(n_1610),
    .Q(i4_dout[2]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[30]  (.CLK(clk_i),
    .D(n_1630),
    .Q(i4_dout[30]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[31]  (.CLK(clk_i),
    .D(n_1544),
    .Q(i4_dout[31]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[3]  (.CLK(clk_i),
    .D(n_1632),
    .Q(i4_dout[3]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[4]  (.CLK(clk_i),
    .D(n_1554),
    .Q(i4_dout[4]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[5]  (.CLK(clk_i),
    .D(n_1633),
    .Q(i4_dout[5]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[6]  (.CLK(clk_i),
    .D(n_1551),
    .Q(i4_dout[6]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[7]  (.CLK(clk_i),
    .D(n_1635),
    .Q(i4_dout[7]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[8]  (.CLK(clk_i),
    .D(n_1540),
    .Q(i4_dout[8]));
 DFFHQx4_ASAP7_75t_SL \u10_dout_reg[9]  (.CLK(clk_i),
    .D(n_1594),
    .Q(i4_dout[9]));
 DFFHQNx2_ASAP7_75t_SL u10_empty_reg (.CLK(clk_i),
    .D(n_20245),
    .QN(i4_empty));
 DFFHQNx1_ASAP7_75t_SL u10_full_reg (.CLK(clk_i),
    .D(n_20246),
    .QN(i4_full));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_4489),
    .QN(\u10_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_46480),
    .QN(\u10_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_18591),
    .QN(\u10_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_28235),
    .QN(\u10_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_4475),
    .QN(\u10_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_4474),
    .QN(\u10_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_4473),
    .QN(\u10_mem[0] [15]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_4472),
    .QN(\u10_mem[0] [16]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_4470),
    .QN(\u10_mem[0] [17]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_11697),
    .QN(\u10_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_16664),
    .QN(\u10_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_4502),
    .QN(\u10_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_4588),
    .QN(\u10_mem[0] [20]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_4604),
    .QN(\u10_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_4603),
    .QN(\u10_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_4600),
    .QN(\u10_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_4599),
    .QN(\u10_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_4598),
    .QN(\u10_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_4597),
    .QN(\u10_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_4596),
    .QN(\u10_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_4595),
    .QN(\u10_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_4594),
    .QN(\u10_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_4488),
    .QN(\u10_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_4593),
    .QN(\u10_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_4592),
    .QN(\u10_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_4498),
    .QN(\u10_mem[0] [3]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_4500),
    .QN(\u10_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_4483),
    .QN(\u10_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_21938),
    .QN(\u10_mem[0] [6]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_4481),
    .QN(\u10_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_21947),
    .QN(\u10_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_18068),
    .QN(\u10_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_61889),
    .QN(\u10_mem[1] [0]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_61883),
    .QN(\u10_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_4656),
    .QN(\u10_mem[1] [11]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_4721),
    .QN(\u10_mem[1] [12]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_4719),
    .QN(\u10_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_4717),
    .QN(\u10_mem[1] [14]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_4715),
    .QN(\u10_mem[1] [15]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_4713),
    .QN(\u10_mem[1] [16]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_4711),
    .QN(\u10_mem[1] [17]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_11699),
    .QN(\u10_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_4707),
    .QN(\u10_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_61887),
    .QN(\u10_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_61895),
    .QN(\u10_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_4674),
    .QN(\u10_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_61901),
    .QN(\u10_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_4670),
    .QN(\u10_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_62124),
    .QN(\u10_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_61963),
    .QN(\u10_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_4664),
    .QN(\u10_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_4662),
    .QN(\u10_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_61957),
    .QN(\u10_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_60456),
    .QN(\u10_mem[1] [29]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_62657),
    .QN(\u10_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_4658),
    .QN(\u10_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_4657),
    .QN(\u10_mem[1] [31]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_61885),
    .QN(\u10_mem[1] [3]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_50660),
    .QN(\u10_mem[1] [4]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_78622),
    .QN(\u10_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_44556),
    .QN(\u10_mem[1] [6]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_42801),
    .QN(\u10_mem[1] [7]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_4807),
    .QN(\u10_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_46750),
    .QN(\u10_mem[1] [9]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_48177),
    .QN(\u10_mem[2] [0]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_48171),
    .QN(\u10_mem[2] [10]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_48163),
    .QN(\u10_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_48158),
    .QN(\u10_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_48172),
    .QN(\u10_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_48161),
    .QN(\u10_mem[2] [14]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_48173),
    .QN(\u10_mem[2] [15]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_48156),
    .QN(\u10_mem[2] [16]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_48157),
    .QN(\u10_mem[2] [17]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_48170),
    .QN(\u10_mem[2] [18]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_48162),
    .QN(\u10_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_48159),
    .QN(\u10_mem[2] [1]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_48148),
    .QN(\u10_mem[2] [20]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_48152),
    .QN(\u10_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_48150),
    .QN(\u10_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_48149),
    .QN(\u10_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_47772),
    .QN(\u10_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_48165),
    .QN(\u10_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_48166),
    .QN(\u10_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_48168),
    .QN(\u10_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_48169),
    .QN(\u10_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_48147),
    .QN(\u10_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_62615),
    .QN(\u10_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_48151),
    .QN(\u10_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_48167),
    .QN(\u10_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_48164),
    .QN(\u10_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_48175),
    .QN(\u10_mem[2] [4]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_48176),
    .QN(\u10_mem[2] [5]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_48174),
    .QN(\u10_mem[2] [6]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_48160),
    .QN(\u10_mem[2] [7]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_48154),
    .QN(\u10_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_48155),
    .QN(\u10_mem[2] [9]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_25004),
    .QN(\u10_mem[3] [0]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_24992),
    .QN(\u10_mem[3] [10]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_61245),
    .QN(\u10_mem[3] [11]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_24991),
    .QN(\u10_mem[3] [12]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_24990),
    .QN(\u10_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_24989),
    .QN(\u10_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_24988),
    .QN(\u10_mem[3] [15]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_24987),
    .QN(\u10_mem[3] [16]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_24986),
    .QN(\u10_mem[3] [17]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_24985),
    .QN(\u10_mem[3] [18]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_24978),
    .QN(\u10_mem[3] [19]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_25002),
    .QN(\u10_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_24984),
    .QN(\u10_mem[3] [20]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_25008),
    .QN(\u10_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_25005),
    .QN(\u10_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_35122),
    .QN(\u10_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_24981),
    .QN(\u10_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_25007),
    .QN(\u10_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_25006),
    .QN(\u10_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_24982),
    .QN(\u10_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_25010),
    .QN(\u10_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_24979),
    .QN(\u10_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_25001),
    .QN(\u10_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_25009),
    .QN(\u10_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_24980),
    .QN(\u10_mem[3] [31]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_35393),
    .QN(\u10_mem[3] [3]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_24999),
    .QN(\u10_mem[3] [4]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_24998),
    .QN(\u10_mem[3] [5]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_24997),
    .QN(\u10_mem[3] [6]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_36405),
    .QN(\u10_mem[3] [7]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_24995),
    .QN(\u10_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u10_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_24993),
    .QN(\u10_mem[3] [9]));
 DFFHQx4_ASAP7_75t_SL \u10_rp_reg[0]  (.CLK(clk_i),
    .D(n_21148),
    .Q(u10_rp[0]));
 DFFHQNx2_ASAP7_75t_SL \u10_rp_reg[1]  (.CLK(clk_i),
    .D(n_29940),
    .QN(u10_rp[1]));
 DFFHQNx1_ASAP7_75t_SL \u10_rp_reg[2]  (.CLK(clk_i),
    .D(n_47500),
    .QN(u10_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u10_status_reg[0]  (.CLK(clk_i),
    .D(n_20247),
    .QN(i4_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u10_status_reg[1]  (.CLK(clk_i),
    .D(n_21695),
    .QN(i4_status[1]));
 DFFHQNx1_ASAP7_75t_SL \u10_wp_reg[0]  (.CLK(clk_i),
    .D(n_4578),
    .QN(u10_wp[0]));
 DFFHQx4_ASAP7_75t_SL \u10_wp_reg[1]  (.CLK(clk_i),
    .D(n_19047),
    .Q(u10_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u10_wp_reg[2]  (.CLK(clk_i),
    .D(n_26646),
    .QN(u10_wp[2]));
 DFFHQx4_ASAP7_75t_SL \u10_wp_reg[3]  (.CLK(clk_i),
    .D(n_4579),
    .Q(u10_wp[3]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[0]  (.CLK(clk_i),
    .D(n_29089),
    .QN(u11_din_tmp1[0]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[10]  (.CLK(clk_i),
    .D(n_29083),
    .QN(u11_din_tmp1[10]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[11]  (.CLK(clk_i),
    .D(n_29105),
    .QN(u11_din_tmp1[11]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[12]  (.CLK(clk_i),
    .D(n_29095),
    .QN(u11_din_tmp1[12]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[13]  (.CLK(clk_i),
    .D(n_29103),
    .QN(u11_din_tmp1[13]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[14]  (.CLK(clk_i),
    .D(n_29093),
    .QN(u11_din_tmp1[14]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[15]  (.CLK(clk_i),
    .D(n_29077),
    .QN(u11_din_tmp1[15]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[1]  (.CLK(clk_i),
    .D(n_34483),
    .QN(u11_din_tmp1[1]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[2]  (.CLK(clk_i),
    .D(n_29079),
    .QN(u11_din_tmp1[2]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[3]  (.CLK(clk_i),
    .D(n_34487),
    .QN(u11_din_tmp1[3]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[4]  (.CLK(clk_i),
    .D(n_29107),
    .QN(u11_din_tmp1[4]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[5]  (.CLK(clk_i),
    .D(n_29097),
    .QN(u11_din_tmp1[5]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[6]  (.CLK(clk_i),
    .D(n_29099),
    .QN(u11_din_tmp1[6]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[7]  (.CLK(clk_i),
    .D(n_36291),
    .QN(u11_din_tmp1[7]));
 DFFHQNx2_ASAP7_75t_SL \u11_din_tmp1_reg[8]  (.CLK(clk_i),
    .D(n_29101),
    .QN(u11_din_tmp1[8]));
 DFFHQNx1_ASAP7_75t_SL \u11_din_tmp1_reg[9]  (.CLK(clk_i),
    .D(n_29081),
    .QN(u11_din_tmp1[9]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[0]  (.CLK(clk_i),
    .D(n_1585),
    .Q(i6_dout[0]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[10]  (.CLK(clk_i),
    .D(n_1576),
    .Q(i6_dout[10]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[11]  (.CLK(clk_i),
    .D(n_1634),
    .Q(i6_dout[11]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[12]  (.CLK(clk_i),
    .D(n_1575),
    .Q(i6_dout[12]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[13]  (.CLK(clk_i),
    .D(n_1574),
    .Q(i6_dout[13]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[14]  (.CLK(clk_i),
    .D(n_1572),
    .Q(i6_dout[14]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[15]  (.CLK(clk_i),
    .D(n_1571),
    .Q(i6_dout[15]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[16]  (.CLK(clk_i),
    .D(n_1570),
    .Q(i6_dout[16]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[17]  (.CLK(clk_i),
    .D(n_1569),
    .Q(i6_dout[17]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[18]  (.CLK(clk_i),
    .D(n_1568),
    .Q(i6_dout[18]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[19]  (.CLK(clk_i),
    .D(n_1553),
    .Q(i6_dout[19]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[1]  (.CLK(clk_i),
    .D(n_1584),
    .Q(i6_dout[1]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[20]  (.CLK(clk_i),
    .D(n_1567),
    .Q(i6_dout[20]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[21]  (.CLK(clk_i),
    .D(n_1566),
    .Q(i6_dout[21]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[22]  (.CLK(clk_i),
    .D(n_1565),
    .Q(i6_dout[22]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[23]  (.CLK(clk_i),
    .D(n_1555),
    .Q(i6_dout[23]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[24]  (.CLK(clk_i),
    .D(n_1516),
    .Q(i6_dout[24]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[25]  (.CLK(clk_i),
    .D(n_1564),
    .Q(i6_dout[25]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[26]  (.CLK(clk_i),
    .D(n_1563),
    .Q(i6_dout[26]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[27]  (.CLK(clk_i),
    .D(n_1660),
    .Q(i6_dout[27]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[28]  (.CLK(clk_i),
    .D(n_1548),
    .Q(i6_dout[28]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[29]  (.CLK(clk_i),
    .D(n_1561),
    .Q(i6_dout[29]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[2]  (.CLK(clk_i),
    .D(n_1583),
    .Q(i6_dout[2]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[30]  (.CLK(clk_i),
    .D(n_1589),
    .Q(i6_dout[30]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[31]  (.CLK(clk_i),
    .D(n_1559),
    .Q(i6_dout[31]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[3]  (.CLK(clk_i),
    .D(n_1582),
    .Q(i6_dout[3]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[4]  (.CLK(clk_i),
    .D(n_1581),
    .Q(i6_dout[4]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[5]  (.CLK(clk_i),
    .D(n_1550),
    .Q(i6_dout[5]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[6]  (.CLK(clk_i),
    .D(n_1580),
    .Q(i6_dout[6]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[7]  (.CLK(clk_i),
    .D(n_1579),
    .Q(i6_dout[7]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[8]  (.CLK(clk_i),
    .D(n_1578),
    .Q(i6_dout[8]));
 DFFHQx4_ASAP7_75t_SL \u11_dout_reg[9]  (.CLK(clk_i),
    .D(n_1577),
    .Q(i6_dout[9]));
 DFFHQNx1_ASAP7_75t_SL u11_empty_reg (.CLK(clk_i),
    .D(n_10936),
    .QN(i6_empty));
 DFFHQNx1_ASAP7_75t_SL u11_full_reg (.CLK(clk_i),
    .D(n_1558),
    .QN(i6_full));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_29019),
    .QN(\u11_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_29009),
    .QN(\u11_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_29041),
    .QN(\u11_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_29022),
    .QN(\u11_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_29013),
    .QN(\u11_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_29020),
    .QN(\u11_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_29016),
    .QN(\u11_mem[0] [15]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_29018),
    .QN(\u11_mem[0] [16]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_29036),
    .QN(\u11_mem[0] [17]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_29015),
    .QN(\u11_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_29028),
    .QN(\u11_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_29012),
    .QN(\u11_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_29030),
    .QN(\u11_mem[0] [20]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_29037),
    .QN(\u11_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_29038),
    .QN(\u11_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_29027),
    .QN(\u11_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_29035),
    .QN(\u11_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_29032),
    .QN(\u11_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_29029),
    .QN(\u11_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_29040),
    .QN(\u11_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_29031),
    .QN(\u11_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_29026),
    .QN(\u11_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_29017),
    .QN(\u11_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_29039),
    .QN(\u11_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_29034),
    .QN(\u11_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_29014),
    .QN(\u11_mem[0] [3]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_29023),
    .QN(\u11_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_29033),
    .QN(\u11_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_29025),
    .QN(\u11_mem[0] [6]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_29024),
    .QN(\u11_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_29021),
    .QN(\u11_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_29010),
    .QN(\u11_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_4840),
    .QN(\u11_mem[1] [0]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_4860),
    .QN(\u11_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_4863),
    .QN(\u11_mem[1] [11]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_18483),
    .QN(\u11_mem[1] [12]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_4870),
    .QN(\u11_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_4875),
    .QN(\u11_mem[1] [14]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_4878),
    .QN(\u11_mem[1] [15]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_21554),
    .QN(\u11_mem[1] [16]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_4882),
    .QN(\u11_mem[1] [17]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_4884),
    .QN(\u11_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_4886),
    .QN(\u11_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_4842),
    .QN(\u11_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_4928),
    .QN(\u11_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_4929),
    .QN(\u11_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_4932),
    .QN(\u11_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_4936),
    .QN(\u11_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_4937),
    .QN(\u11_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_4938),
    .QN(\u11_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_4939),
    .QN(\u11_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_4940),
    .QN(\u11_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_4942),
    .QN(\u11_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_4945),
    .QN(\u11_mem[1] [29]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_4844),
    .QN(\u11_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_4950),
    .QN(\u11_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_4952),
    .QN(\u11_mem[1] [31]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_4846),
    .QN(\u11_mem[1] [3]));
 DFFHQNx1_ASAP7_75t_SL \u11_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_4848),
    .QN(\u11_mem[1] [4]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_4850),
    .QN(\u11_mem[1] [5]));
 DFFHQNx1_ASAP7_75t_SL \u11_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_4852),
    .QN(\u11_mem[1] [6]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_7501),
    .QN(\u11_mem[1] [7]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_4856),
    .QN(\u11_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_16439),
    .QN(\u11_mem[1] [9]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_61786),
    .QN(\u11_mem[2] [0]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_21320),
    .QN(\u11_mem[2] [10]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_12837),
    .QN(\u11_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_12859),
    .QN(\u11_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_12858),
    .QN(\u11_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_28521),
    .QN(\u11_mem[2] [14]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_12854),
    .QN(\u11_mem[2] [15]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_12856),
    .QN(\u11_mem[2] [16]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_12855),
    .QN(\u11_mem[2] [17]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_12857),
    .QN(\u11_mem[2] [18]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_45627),
    .QN(\u11_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_12867),
    .QN(\u11_mem[2] [1]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_61773),
    .QN(\u11_mem[2] [20]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_12846),
    .QN(\u11_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_12842),
    .QN(\u11_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_12839),
    .QN(\u11_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_12838),
    .QN(\u11_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_45569),
    .QN(\u11_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_12848),
    .QN(\u11_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_12843),
    .QN(\u11_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_12847),
    .QN(\u11_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_12845),
    .QN(\u11_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_12865),
    .QN(\u11_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_12849),
    .QN(\u11_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_45607),
    .QN(\u11_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_27880),
    .QN(\u11_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_21328),
    .QN(\u11_mem[2] [4]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_12851),
    .QN(\u11_mem[2] [5]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_12863),
    .QN(\u11_mem[2] [6]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_26556),
    .QN(\u11_mem[2] [7]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_21324),
    .QN(\u11_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_12861),
    .QN(\u11_mem[2] [9]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_4824),
    .QN(\u11_mem[3] [0]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_5098),
    .QN(\u11_mem[3] [10]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_5097),
    .QN(\u11_mem[3] [11]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_5094),
    .QN(\u11_mem[3] [12]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_4829),
    .QN(\u11_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_18092),
    .QN(\u11_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_4831),
    .QN(\u11_mem[3] [15]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_4832),
    .QN(\u11_mem[3] [16]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_4833),
    .QN(\u11_mem[3] [17]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_4834),
    .QN(\u11_mem[3] [18]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_4835),
    .QN(\u11_mem[3] [19]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_4823),
    .QN(\u11_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_4900),
    .QN(\u11_mem[3] [20]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_4902),
    .QN(\u11_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_4904),
    .QN(\u11_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_4906),
    .QN(\u11_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_4908),
    .QN(\u11_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_4910),
    .QN(\u11_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_4912),
    .QN(\u11_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_4914),
    .QN(\u11_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_4916),
    .QN(\u11_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_4918),
    .QN(\u11_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_15137),
    .QN(\u11_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_4920),
    .QN(\u11_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_4922),
    .QN(\u11_mem[3] [31]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_15141),
    .QN(\u11_mem[3] [3]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_4819),
    .QN(\u11_mem[3] [4]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_4817),
    .QN(\u11_mem[3] [5]));
 DFFHQNx1_ASAP7_75t_SL \u11_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_4818),
    .QN(\u11_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u11_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_7500),
    .QN(\u11_mem[3] [7]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_4825),
    .QN(\u11_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u11_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_4992),
    .QN(\u11_mem[3] [9]));
 DFFHQx4_ASAP7_75t_SL \u11_rp_reg[0]  (.CLK(clk_i),
    .D(n_2706),
    .Q(u11_rp[0]));
 DFFHQNx2_ASAP7_75t_SL \u11_rp_reg[1]  (.CLK(clk_i),
    .D(n_11478),
    .QN(u11_rp[1]));
 DFFHQNx1_ASAP7_75t_SL \u11_rp_reg[2]  (.CLK(clk_i),
    .D(n_2957),
    .QN(u11_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u11_status_reg[0]  (.CLK(clk_i),
    .D(n_707),
    .QN(i6_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u11_status_reg[1]  (.CLK(clk_i),
    .D(n_21541),
    .QN(i6_status[1]));
 DFFHQNx1_ASAP7_75t_SL \u11_wp_reg[0]  (.CLK(clk_i),
    .D(n_18655),
    .QN(u11_wp[0]));
 DFFHQx4_ASAP7_75t_SL \u11_wp_reg[1]  (.CLK(clk_i),
    .D(n_28951),
    .Q(u11_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u11_wp_reg[2]  (.CLK(clk_i),
    .D(n_20597),
    .QN(u11_wp[2]));
 DFFHQx4_ASAP7_75t_SL \u11_wp_reg[3]  (.CLK(clk_i),
    .D(n_4641),
    .Q(u11_wp[3]));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[0]  (.CLK(clk_i),
    .D(n_128),
    .QN(wb_din[0]));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[10]  (.CLK(clk_i),
    .D(n_65970),
    .QN(n_65971));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[11]  (.CLK(clk_i),
    .D(n_65964),
    .QN(n_65965));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[12]  (.CLK(clk_i),
    .D(n_65995),
    .QN(n_65996));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[13]  (.CLK(clk_i),
    .D(n_65953),
    .QN(n_65954));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[14]  (.CLK(clk_i),
    .D(n_66030),
    .QN(n_66031));
 DFFHQNx2_ASAP7_75t_SL \u12_dout_reg[15]  (.CLK(clk_i),
    .D(n_65989),
    .QN(n_65990));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[16]  (.CLK(clk_i),
    .D(n_65947),
    .QN(n_65948));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[17]  (.CLK(clk_i),
    .D(n_65950),
    .QN(n_65951));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[18]  (.CLK(clk_i),
    .D(n_65933),
    .QN(n_65934));
 DFFHQNx2_ASAP7_75t_SL \u12_dout_reg[19]  (.CLK(clk_i),
    .D(n_65931),
    .QN(n_65932));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[1]  (.CLK(clk_i),
    .D(n_64),
    .QN(wb_din[1]));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[20]  (.CLK(clk_i),
    .D(n_66023),
    .QN(n_66024));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[21]  (.CLK(clk_i),
    .D(n_66014),
    .QN(n_66015));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[22]  (.CLK(clk_i),
    .D(n_65936),
    .QN(n_65937));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[23]  (.CLK(clk_i),
    .D(n_65928),
    .QN(n_65929));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[24]  (.CLK(clk_i),
    .D(n_65911),
    .QN(n_65912));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[25]  (.CLK(clk_i),
    .D(n_65921),
    .QN(n_65922));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[26]  (.CLK(clk_i),
    .D(n_66007),
    .QN(n_66008));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[27]  (.CLK(clk_i),
    .D(n_65905),
    .QN(n_65906));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[28]  (.CLK(clk_i),
    .D(n_65918),
    .QN(n_65919));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[29]  (.CLK(clk_i),
    .D(n_44),
    .QN(wb_din[29]));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[2]  (.CLK(clk_i),
    .D(n_65998),
    .QN(n_65999));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[30]  (.CLK(clk_i),
    .D(n_140),
    .QN(wb_din[30]));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[31]  (.CLK(clk_i),
    .D(n_65898),
    .QN(n_65899));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[3]  (.CLK(clk_i),
    .D(n_65961),
    .QN(n_65962));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[4]  (.CLK(clk_i),
    .D(n_65983),
    .QN(n_65984));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[5]  (.CLK(clk_i),
    .D(n_65958),
    .QN(n_65959));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[6]  (.CLK(clk_i),
    .D(n_66001),
    .QN(n_66002));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[7]  (.CLK(clk_i),
    .D(n_65967),
    .QN(n_65968));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[8]  (.CLK(clk_i),
    .D(n_65977),
    .QN(n_65978));
 DFFHQNx1_ASAP7_75t_SL \u12_dout_reg[9]  (.CLK(clk_i),
    .D(n_65992),
    .QN(n_65993));
 DFFHQNx2_ASAP7_75t_SL u12_i3_re_reg (.CLK(clk_i),
    .D(n_7221),
    .QN(i3_re));
 DFFHQNx2_ASAP7_75t_SL u12_i4_re_reg (.CLK(clk_i),
    .D(n_1857),
    .QN(i4_re));
 DFFHQNx2_ASAP7_75t_SL u12_i6_re_reg (.CLK(clk_i),
    .D(n_14935),
    .QN(i6_re));
 DFFHQx4_ASAP7_75t_SL u12_o3_we_reg (.CLK(clk_i),
    .D(n_2155),
    .Q(o3_we));
 DFFHQx4_ASAP7_75t_SL u12_o4_we_reg (.CLK(clk_i),
    .D(n_24627),
    .Q(o4_we));
 DFFHQx4_ASAP7_75t_SL u12_o6_we_reg (.CLK(clk_i),
    .D(n_13792),
    .Q(o6_we));
 DFFHQx4_ASAP7_75t_SL u12_o7_we_reg (.CLK(clk_i),
    .D(n_47778),
    .Q(o7_we));
 DFFHQx4_ASAP7_75t_SL u12_o8_we_reg (.CLK(clk_i),
    .D(n_13796),
    .Q(o8_we));
 DFFHQx4_ASAP7_75t_SL u12_o9_we_reg (.CLK(clk_i),
    .D(n_13794),
    .Q(o9_we));
 DFFHQNx1_ASAP7_75t_SL u12_re1_reg (.CLK(clk_i),
    .D(n_35638),
    .QN(u12_re1));
 DFFHQNx1_ASAP7_75t_SL u12_re2_reg (.CLK(clk_i),
    .D(n_35634),
    .QN(u12_re2));
 DFFHQx4_ASAP7_75t_SL u12_rf_we_reg (.CLK(clk_i),
    .D(n_1869),
    .Q(rf_we));
 DFFHQNx2_ASAP7_75t_SL u12_wb_ack_o_reg (.CLK(clk_i),
    .D(n_2216),
    .QN(u12_wb_ack_o_745));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[0]  (.CLK(clk_i),
    .D(n_16725),
    .Q(\u12_wb_data_o[0]_713 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[10]  (.CLK(clk_i),
    .D(n_14985),
    .Q(\u12_wb_data_o[10]_723 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[11]  (.CLK(clk_i),
    .D(n_22846),
    .Q(\u12_wb_data_o[11]_724 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[12]  (.CLK(clk_i),
    .D(n_2721),
    .Q(\u12_wb_data_o[12]_725 ));
 DFFHQx4_ASAP7_75t_L \u12_wb_data_o_reg[13]  (.CLK(clk_i),
    .D(n_8251),
    .Q(\u12_wb_data_o[13]_726 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[14]  (.CLK(clk_i),
    .D(n_2712),
    .Q(\u12_wb_data_o[14]_727 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[15]  (.CLK(clk_i),
    .D(n_52951),
    .Q(\u12_wb_data_o[15]_728 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[16]  (.CLK(clk_i),
    .D(n_49175),
    .QN(\u12_wb_data_o[16]_729 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[17]  (.CLK(clk_i),
    .D(n_2724),
    .Q(\u12_wb_data_o[17]_730 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[18]  (.CLK(clk_i),
    .D(n_22029),
    .Q(\u12_wb_data_o[18]_731 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[19]  (.CLK(clk_i),
    .D(n_43172),
    .Q(\u12_wb_data_o[19]_732 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[1]  (.CLK(clk_i),
    .D(n_2683),
    .Q(\u12_wb_data_o[1]_714 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[20]  (.CLK(clk_i),
    .D(n_2931),
    .QN(\u12_wb_data_o[20]_733 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[21]  (.CLK(clk_i),
    .D(n_2932),
    .QN(\u12_wb_data_o[21]_734 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[22]  (.CLK(clk_i),
    .D(n_2933),
    .QN(\u12_wb_data_o[22]_735 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[23]  (.CLK(clk_i),
    .D(n_2977),
    .Q(\u12_wb_data_o[23]_736 ));
 DFFHQx4_ASAP7_75t_L \u12_wb_data_o_reg[24]  (.CLK(clk_i),
    .D(n_2727),
    .Q(\u12_wb_data_o[24]_737 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[25]  (.CLK(clk_i),
    .D(n_2934),
    .QN(\u12_wb_data_o[25]_738 ));
 DFFHQNx1_ASAP7_75t_SL \u12_wb_data_o_reg[26]  (.CLK(clk_i),
    .D(n_2935),
    .QN(\u12_wb_data_o[26]_739 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[27]  (.CLK(clk_i),
    .D(n_8280),
    .QN(\u12_wb_data_o[27]_740 ));
 DFFHQNx1_ASAP7_75t_SL \u12_wb_data_o_reg[28]  (.CLK(clk_i),
    .D(n_8333),
    .QN(\u12_wb_data_o[28]_741 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[29]  (.CLK(clk_i),
    .D(n_7227),
    .QN(\u12_wb_data_o[29]_742 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[2]  (.CLK(clk_i),
    .D(n_2715),
    .Q(\u12_wb_data_o[2]_715 ));
 DFFHQNx2_ASAP7_75t_SL \u12_wb_data_o_reg[30]  (.CLK(clk_i),
    .D(n_7226),
    .QN(\u12_wb_data_o[30]_743 ));
 DFFHQx4_ASAP7_75t_L \u12_wb_data_o_reg[31]  (.CLK(clk_i),
    .D(n_2653),
    .Q(\u12_wb_data_o[31]_744 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[3]  (.CLK(clk_i),
    .D(n_16733),
    .Q(\u12_wb_data_o[3]_716 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[4]  (.CLK(clk_i),
    .D(n_2716),
    .Q(\u12_wb_data_o[4]_717 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[5]  (.CLK(clk_i),
    .D(n_8255),
    .Q(\u12_wb_data_o[5]_718 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[6]  (.CLK(clk_i),
    .D(n_16728),
    .Q(\u12_wb_data_o[6]_719 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[7]  (.CLK(clk_i),
    .D(n_2713),
    .Q(\u12_wb_data_o[7]_720 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[8]  (.CLK(clk_i),
    .D(n_16723),
    .Q(\u12_wb_data_o[8]_721 ));
 DFFHQx4_ASAP7_75t_SL \u12_wb_data_o_reg[9]  (.CLK(clk_i),
    .D(n_2719),
    .Q(\u12_wb_data_o[9]_722 ));
 DFFHQNx1_ASAP7_75t_SL u12_we1_reg (.CLK(clk_i),
    .D(n_18889),
    .QN(u12_we1));
 DFFHQNx1_ASAP7_75t_SL u12_we2_reg (.CLK(clk_i),
    .D(n_13413),
    .QN(u12_we2));
 DFFHQNx2_ASAP7_75t_SL u13_ac97_rst_force_reg (.CLK(clk_i),
    .D(n_10916),
    .QN(ac97_rst_force));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[0]  (.CLK(clk_i),
    .D(n_22919),
    .QN(crac_out[0]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[10]  (.CLK(clk_i),
    .D(n_66820),
    .QN(crac_out[10]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[11]  (.CLK(clk_i),
    .D(n_17577),
    .QN(crac_out[11]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[12]  (.CLK(clk_i),
    .D(n_17525),
    .QN(crac_out[12]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[13]  (.CLK(clk_i),
    .D(n_17583),
    .QN(crac_out[13]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[14]  (.CLK(clk_i),
    .D(n_17534),
    .QN(crac_out[14]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[15]  (.CLK(clk_i),
    .D(n_17542),
    .QN(crac_out[15]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[1]  (.CLK(clk_i),
    .D(n_17513),
    .QN(crac_out[1]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[2]  (.CLK(clk_i),
    .D(n_17532),
    .QN(crac_out[2]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[3]  (.CLK(clk_i),
    .D(n_17563),
    .QN(crac_out[3]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[4]  (.CLK(clk_i),
    .D(n_69012),
    .QN(crac_out[4]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[5]  (.CLK(clk_i),
    .D(n_17567),
    .QN(crac_out[5]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[6]  (.CLK(clk_i),
    .D(n_17528),
    .QN(crac_out[6]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[7]  (.CLK(clk_i),
    .D(n_28368),
    .QN(crac_out[7]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[8]  (.CLK(clk_i),
    .D(n_17530),
    .QN(crac_out[8]));
 DFFHQNx2_ASAP7_75t_SL \u13_crac_dout_r_reg[9]  (.CLK(clk_i),
    .D(n_17565),
    .QN(crac_out[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[0]  (.CLK(clk_i),
    .D(n_16819),
    .QN(crac_out[16]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[1]  (.CLK(clk_i),
    .D(n_16807),
    .QN(crac_out[17]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[2]  (.CLK(clk_i),
    .D(n_46163),
    .QN(crac_out[18]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[3]  (.CLK(clk_i),
    .D(n_16828),
    .QN(crac_out[19]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[4]  (.CLK(clk_i),
    .D(n_16788),
    .QN(crac_out[20]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[5]  (.CLK(clk_i),
    .D(n_62634),
    .QN(crac_out[21]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[6]  (.CLK(clk_i),
    .D(n_66799),
    .QN(crac_out[22]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_crac_r_reg[7]  (.CLK(clk_i),
    .D(n_16816),
    .QN(crac_out[31]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[0]  (.CLK(clk_i),
    .D(n_8192),
    .QN(ic0_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[10]  (.CLK(clk_i),
    .D(n_9936),
    .QN(ic1_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[11]  (.CLK(clk_i),
    .D(n_10022),
    .QN(ic1_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[12]  (.CLK(clk_i),
    .D(n_10050),
    .QN(ic1_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[13]  (.CLK(clk_i),
    .D(n_10107),
    .QN(ic1_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[14]  (.CLK(clk_i),
    .D(n_9760),
    .QN(ic1_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[15]  (.CLK(clk_i),
    .D(n_9790),
    .QN(u13_icc_r[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[16]  (.CLK(clk_i),
    .D(n_10138),
    .QN(ic2_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[17]  (.CLK(clk_i),
    .D(n_10165),
    .QN(ic2_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[18]  (.CLK(clk_i),
    .D(n_10192),
    .QN(ic2_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[19]  (.CLK(clk_i),
    .D(n_10218),
    .QN(ic2_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[1]  (.CLK(clk_i),
    .D(n_14099),
    .QN(ic0_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[20]  (.CLK(clk_i),
    .D(n_10244),
    .QN(ic2_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[21]  (.CLK(clk_i),
    .D(n_10272),
    .QN(ic2_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[22]  (.CLK(clk_i),
    .D(n_66804),
    .QN(ic2_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[23]  (.CLK(clk_i),
    .D(n_10327),
    .QN(u13_icc_r[23]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[2]  (.CLK(clk_i),
    .D(n_9849),
    .QN(ic0_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[3]  (.CLK(clk_i),
    .D(n_9877),
    .QN(ic0_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[4]  (.CLK(clk_i),
    .D(n_68227),
    .QN(ic0_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[5]  (.CLK(clk_i),
    .D(n_10079),
    .QN(ic0_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[6]  (.CLK(clk_i),
    .D(n_9731),
    .QN(ic0_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[7]  (.CLK(clk_i),
    .D(n_9817),
    .QN(u13_icc_r[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[8]  (.CLK(clk_i),
    .D(n_9907),
    .QN(ic1_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_icc_r_reg[9]  (.CLK(clk_i),
    .D(n_9963),
    .QN(ic1_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx2_ASAP7_75t_SL u13_int_reg (.CLK(clk_i),
    .D(n_14227),
    .QN(u13_int_1643));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[0]  (.CLK(clk_i),
    .D(n_32321),
    .QN(u13_intm_r[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[10]  (.CLK(clk_i),
    .D(n_66831),
    .QN(u13_intm_r[10]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[11]  (.CLK(clk_i),
    .D(n_32320),
    .QN(u13_intm_r[11]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[12]  (.CLK(clk_i),
    .D(n_32339),
    .QN(u13_intm_r[12]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[13]  (.CLK(clk_i),
    .D(n_32337),
    .QN(u13_intm_r[13]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[14]  (.CLK(clk_i),
    .D(n_47792),
    .QN(u13_intm_r[14]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[15]  (.CLK(clk_i),
    .D(n_32346),
    .QN(u13_intm_r[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[16]  (.CLK(clk_i),
    .D(n_32336),
    .QN(u13_intm_r[16]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[17]  (.CLK(clk_i),
    .D(n_32334),
    .QN(u13_intm_r[17]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[18]  (.CLK(clk_i),
    .D(n_32333),
    .QN(u13_intm_r[18]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[19]  (.CLK(clk_i),
    .D(n_32332),
    .QN(u13_intm_r[19]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[1]  (.CLK(clk_i),
    .D(n_32322),
    .QN(u13_intm_r[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[20]  (.CLK(clk_i),
    .D(n_32331),
    .QN(u13_intm_r[20]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[21]  (.CLK(clk_i),
    .D(n_32330),
    .QN(u13_intm_r[21]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[22]  (.CLK(clk_i),
    .D(n_66814),
    .QN(u13_intm_r[22]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[23]  (.CLK(clk_i),
    .D(n_32328),
    .QN(u13_intm_r[23]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[24]  (.CLK(clk_i),
    .D(n_32326),
    .QN(u13_intm_r[24]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[25]  (.CLK(clk_i),
    .D(n_32325),
    .QN(u13_intm_r[25]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[26]  (.CLK(clk_i),
    .D(n_32324),
    .QN(u13_intm_r[26]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[27]  (.CLK(clk_i),
    .D(n_32323),
    .QN(u13_intm_r[27]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[28]  (.CLK(clk_i),
    .D(n_32327),
    .QN(u13_intm_r[28]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[2]  (.CLK(clk_i),
    .D(n_32344),
    .QN(u13_intm_r[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[3]  (.CLK(clk_i),
    .D(n_32349),
    .QN(u13_intm_r[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[4]  (.CLK(clk_i),
    .D(n_68223),
    .QN(u13_intm_r[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[5]  (.CLK(clk_i),
    .D(n_32338),
    .QN(u13_intm_r[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[6]  (.CLK(clk_i),
    .D(n_32348),
    .QN(u13_intm_r[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[7]  (.CLK(clk_i),
    .D(n_32345),
    .QN(u13_intm_r[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[8]  (.CLK(clk_i),
    .D(n_32343),
    .QN(u13_intm_r[8]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_intm_r_reg[9]  (.CLK(clk_i),
    .D(n_32341),
    .QN(u13_intm_r[9]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[0]  (.CLK(clk_i),
    .D(n_22179),
    .QN(u13_ints_r[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[10]  (.CLK(clk_i),
    .D(n_22186),
    .QN(u13_ints_r[10]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[11]  (.CLK(clk_i),
    .D(n_22270),
    .QN(u13_ints_r[11]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[12]  (.CLK(clk_i),
    .D(n_22175),
    .QN(u13_ints_r[12]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[13]  (.CLK(clk_i),
    .D(n_22178),
    .QN(u13_ints_r[13]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[14]  (.CLK(clk_i),
    .D(n_22272),
    .QN(u13_ints_r[14]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[15]  (.CLK(clk_i),
    .D(n_22177),
    .QN(u13_ints_r[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[16]  (.CLK(clk_i),
    .D(n_22187),
    .QN(u13_ints_r[16]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[17]  (.CLK(clk_i),
    .D(n_22273),
    .QN(u13_ints_r[17]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[18]  (.CLK(clk_i),
    .D(n_22280),
    .QN(u13_ints_r[18]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[19]  (.CLK(clk_i),
    .D(n_22188),
    .QN(u13_ints_r[19]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[1]  (.CLK(clk_i),
    .D(n_22269),
    .QN(u13_ints_r[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[20]  (.CLK(clk_i),
    .D(n_22278),
    .QN(u13_ints_r[20]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[21]  (.CLK(clk_i),
    .D(n_22282),
    .QN(u13_ints_r[21]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[22]  (.CLK(clk_i),
    .D(n_22176),
    .QN(u13_ints_r[22]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[23]  (.CLK(clk_i),
    .D(n_22277),
    .QN(u13_ints_r[23]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[24]  (.CLK(clk_i),
    .D(n_22189),
    .QN(u13_ints_r[24]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[25]  (.CLK(clk_i),
    .D(n_22190),
    .QN(u13_ints_r[25]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[26]  (.CLK(clk_i),
    .D(n_22279),
    .QN(u13_ints_r[26]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[27]  (.CLK(clk_i),
    .D(n_22281),
    .QN(u13_ints_r[27]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[28]  (.CLK(clk_i),
    .D(n_22283),
    .QN(u13_ints_r[28]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[2]  (.CLK(clk_i),
    .D(n_22271),
    .QN(u13_ints_r[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[3]  (.CLK(clk_i),
    .D(n_22180),
    .QN(u13_ints_r[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[4]  (.CLK(clk_i),
    .D(n_22181),
    .QN(u13_ints_r[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[5]  (.CLK(clk_i),
    .D(n_22275),
    .QN(u13_ints_r[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[6]  (.CLK(clk_i),
    .D(n_22182),
    .QN(u13_ints_r[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[7]  (.CLK(clk_i),
    .D(n_22184),
    .QN(u13_ints_r[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[8]  (.CLK(clk_i),
    .D(n_22274),
    .QN(u13_ints_r[8]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_ints_r_reg[9]  (.CLK(clk_i),
    .D(n_22185),
    .QN(u13_ints_r[9]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[0]  (.CLK(clk_i),
    .D(n_12455),
    .QN(oc0_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[10]  (.CLK(clk_i),
    .D(n_66834),
    .QN(oc1_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[11]  (.CLK(clk_i),
    .D(n_35460),
    .QN(oc1_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[12]  (.CLK(clk_i),
    .D(n_12450),
    .QN(oc1_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[13]  (.CLK(clk_i),
    .D(n_12448),
    .QN(oc1_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[14]  (.CLK(clk_i),
    .D(n_12453),
    .QN(oc1_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[15]  (.CLK(clk_i),
    .D(n_12470),
    .QN(u13_occ0_r[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[16]  (.CLK(clk_i),
    .D(n_12463),
    .QN(oc2_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[17]  (.CLK(clk_i),
    .D(n_12447),
    .QN(oc2_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[18]  (.CLK(clk_i),
    .D(n_24753),
    .QN(oc2_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[19]  (.CLK(clk_i),
    .D(n_12445),
    .QN(oc2_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[1]  (.CLK(clk_i),
    .D(n_12456),
    .QN(oc0_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[20]  (.CLK(clk_i),
    .D(n_19005),
    .QN(oc2_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[21]  (.CLK(clk_i),
    .D(n_12461),
    .QN(oc2_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[22]  (.CLK(clk_i),
    .D(n_67249),
    .QN(oc2_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[23]  (.CLK(clk_i),
    .D(n_12459),
    .QN(u13_occ0_r[23]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[24]  (.CLK(clk_i),
    .D(n_12458),
    .QN(oc3_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[25]  (.CLK(clk_i),
    .D(n_12442),
    .QN(oc3_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[26]  (.CLK(clk_i),
    .D(n_12441),
    .QN(oc3_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[27]  (.CLK(clk_i),
    .D(n_12440),
    .QN(oc3_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[28]  (.CLK(clk_i),
    .D(n_24623),
    .QN(oc3_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[29]  (.CLK(clk_i),
    .D(n_12457),
    .QN(oc3_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[2]  (.CLK(clk_i),
    .D(n_12469),
    .QN(oc0_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[30]  (.CLK(clk_i),
    .D(n_12438),
    .QN(oc3_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[31]  (.CLK(clk_i),
    .D(n_12444),
    .QN(u13_occ0_r[31]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[3]  (.CLK(clk_i),
    .D(n_12468),
    .QN(oc0_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[4]  (.CLK(clk_i),
    .D(n_69029),
    .QN(oc0_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[5]  (.CLK(clk_i),
    .D(n_19068),
    .QN(oc0_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[6]  (.CLK(clk_i),
    .D(n_12454),
    .QN(oc0_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[7]  (.CLK(clk_i),
    .D(n_12452),
    .QN(u13_occ0_r[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[8]  (.CLK(clk_i),
    .D(n_29661),
    .QN(oc1_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ0_r_reg[9]  (.CLK(clk_i),
    .D(n_12466),
    .QN(oc1_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[0]  (.CLK(clk_i),
    .D(n_21312),
    .QN(oc4_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[10]  (.CLK(clk_i),
    .D(n_66830),
    .QN(oc5_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[11]  (.CLK(clk_i),
    .D(n_10963),
    .QN(oc5_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[12]  (.CLK(clk_i),
    .D(n_10962),
    .QN(oc5_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[13]  (.CLK(clk_i),
    .D(n_10960),
    .QN(oc5_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[14]  (.CLK(clk_i),
    .D(n_15274),
    .QN(oc5_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[15]  (.CLK(clk_i),
    .D(n_15271),
    .QN(u13_occ1_r[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[1]  (.CLK(clk_i),
    .D(n_10959),
    .QN(oc4_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[2]  (.CLK(clk_i),
    .D(n_10970),
    .QN(oc4_cfg[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[3]  (.CLK(clk_i),
    .D(n_10969),
    .QN(oc4_cfg[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[4]  (.CLK(clk_i),
    .D(n_69017),
    .QN(oc4_cfg[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[5]  (.CLK(clk_i),
    .D(n_10961),
    .QN(oc4_cfg[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[6]  (.CLK(clk_i),
    .D(n_24670),
    .QN(oc4_cfg[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[7]  (.CLK(clk_i),
    .D(n_10971),
    .QN(u13_occ1_r[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[8]  (.CLK(clk_i),
    .D(n_15300),
    .QN(oc5_cfg[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u13_occ1_r_reg[9]  (.CLK(clk_i),
    .D(n_35654),
    .QN(oc5_cfg[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_L u13_resume_req_reg (.CLK(clk_i),
    .D(n_10910),
    .QN(resume_req));
 SDFHx1_ASAP7_75t_SL u14_crac_valid_r_reg (.CLK(clk_i),
    .QN(out_slt0[14]),
    .D(n_112),
    .SE(n_62919),
    .SI(n_280));
 DFFHQNx2_ASAP7_75t_SL u14_crac_wr_r_reg (.CLK(clk_i),
    .D(n_36097),
    .QN(out_slt0[13]));
 DFFHQNx1_ASAP7_75t_SL u14_u0_en_out_l2_reg (.CLK(clk_i),
    .D(n_36103),
    .QN(u14_u0_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u0_en_out_l_reg (.CLK(clk_i),
    .D(n_37111),
    .QN(out_slt0[12]));
 DFFHQNx1_ASAP7_75t_SL u14_u0_full_empty_r_reg (.CLK(clk_i),
    .D(n_36102),
    .QN(u14_u0_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u1_en_out_l2_reg (.CLK(clk_i),
    .D(n_36089),
    .QN(u14_u1_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u1_en_out_l_reg (.CLK(clk_i),
    .D(n_36077),
    .QN(out_slt0[11]));
 DFFHQNx2_ASAP7_75t_SL u14_u1_full_empty_r_reg (.CLK(clk_i),
    .D(n_36081),
    .QN(u14_u1_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u2_en_out_l2_reg (.CLK(clk_i),
    .D(n_62920),
    .QN(u14_u2_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u2_en_out_l_reg (.CLK(clk_i),
    .D(n_36098),
    .QN(out_slt0[9]));
 DFFHQNx2_ASAP7_75t_SL u14_u2_full_empty_r_reg (.CLK(clk_i),
    .D(n_36079),
    .QN(u14_u2_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u3_en_out_l2_reg (.CLK(clk_i),
    .D(n_36094),
    .QN(u14_u3_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u3_en_out_l_reg (.CLK(clk_i),
    .D(n_36080),
    .QN(out_slt0[8]));
 DFFHQNx2_ASAP7_75t_SL u14_u3_full_empty_r_reg (.CLK(clk_i),
    .D(n_36083),
    .QN(u14_u3_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u4_en_out_l2_reg (.CLK(clk_i),
    .D(n_36092),
    .QN(u14_u4_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u4_en_out_l_reg (.CLK(clk_i),
    .D(n_38760),
    .QN(out_slt0[7]));
 DFFHQNx1_ASAP7_75t_SL u14_u4_full_empty_r_reg (.CLK(clk_i),
    .D(n_36101),
    .QN(u14_u4_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u5_en_out_l2_reg (.CLK(clk_i),
    .D(n_36076),
    .QN(u14_u5_en_out_l2));
 DFFHQNx2_ASAP7_75t_SL u14_u5_en_out_l_reg (.CLK(clk_i),
    .D(n_13777),
    .QN(out_slt0[6]));
 DFFHQNx1_ASAP7_75t_SL u14_u5_full_empty_r_reg (.CLK(clk_i),
    .D(n_36086),
    .QN(u14_u5_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u6_en_out_l2_reg (.CLK(clk_i),
    .D(n_7582),
    .QN(u14_u6_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u6_en_out_l_reg (.CLK(clk_i),
    .D(n_13597),
    .QN(u14_u6_en_out_l_44));
 DFFHQNx1_ASAP7_75t_L u14_u6_full_empty_r_reg (.CLK(clk_i),
    .D(n_4070),
    .QN(u14_u6_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u7_en_out_l2_reg (.CLK(clk_i),
    .D(n_12117),
    .QN(u14_u7_en_out_l2));
 DFFHQNx1_ASAP7_75t_SL u14_u7_en_out_l_reg (.CLK(clk_i),
    .D(n_41769),
    .QN(u14_u7_en_out_l_44));
 DFFHQNx1_ASAP7_75t_SL u14_u7_full_empty_r_reg (.CLK(clk_i),
    .D(n_3909),
    .QN(u14_u7_full_empty_r));
 DFFHQNx1_ASAP7_75t_SL u14_u8_en_out_l2_reg (.CLK(clk_i),
    .D(n_28850),
    .QN(u14_u8_en_out_l2));
 DFFHQNx2_ASAP7_75t_SL u14_u8_en_out_l_reg (.CLK(clk_i),
    .D(n_28849),
    .QN(u14_u8_en_out_l_44));
 DFFHQNx1_ASAP7_75t_L u14_u8_full_empty_r_reg (.CLK(clk_i),
    .D(n_3993),
    .QN(u14_u8_full_empty_r));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[0]  (.CLK(clk_i),
    .D(n_42731),
    .QN(crac_din[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[10]  (.CLK(clk_i),
    .D(n_42738),
    .QN(crac_din[10]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[11]  (.CLK(clk_i),
    .D(n_42734),
    .QN(crac_din[11]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[12]  (.CLK(clk_i),
    .D(n_42725),
    .QN(crac_din[12]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[13]  (.CLK(clk_i),
    .D(n_42730),
    .QN(crac_din[13]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[14]  (.CLK(clk_i),
    .D(n_42726),
    .QN(crac_din[14]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[15]  (.CLK(clk_i),
    .D(n_42732),
    .QN(crac_din[15]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[1]  (.CLK(clk_i),
    .D(n_42733),
    .QN(crac_din[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[2]  (.CLK(clk_i),
    .D(n_42739),
    .QN(crac_din[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[3]  (.CLK(clk_i),
    .D(n_42735),
    .QN(crac_din[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[4]  (.CLK(clk_i),
    .D(n_42737),
    .QN(crac_din[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[5]  (.CLK(clk_i),
    .D(n_42727),
    .QN(crac_din[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[6]  (.CLK(clk_i),
    .D(n_42723),
    .QN(crac_din[6]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[7]  (.CLK(clk_i),
    .D(n_42728),
    .QN(crac_din[7]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[8]  (.CLK(clk_i),
    .D(n_42724),
    .QN(crac_din[8]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u15_crac_din_reg[9]  (.CLK(clk_i),
    .D(n_42740),
    .QN(crac_din[9]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQx4_ASAP7_75t_SL u15_crac_rd_done_reg (.CLK(clk_i),
    .D(n_36085),
    .Q(crac_rd_done));
 DFFASRHQNx1_ASAP7_75t_SL u15_crac_rd_reg (.CLK(clk_i),
    .D(n_14816),
    .QN(u15_crac_rd),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx2_ASAP7_75t_SL u15_crac_we_r_reg (.CLK(clk_i),
    .D(n_28367),
    .QN(u15_crac_we_r));
 DFFASRHQNx1_ASAP7_75t_SL u15_crac_wr_reg (.CLK(clk_i),
    .D(n_21515),
    .QN(crac_wr),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL u15_rdd1_reg (.CLK(clk_i),
    .D(n_36084),
    .QN(u15_rdd1),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL u15_rdd2_reg (.CLK(clk_i),
    .D(n_4591),
    .QN(u15_rdd2),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL u15_rdd3_reg (.CLK(clk_i),
    .D(n_36090),
    .QN(u15_rdd3),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx2_ASAP7_75t_SL u15_valid_r_reg (.CLK(clk_i),
    .D(n_36082),
    .QN(u15_valid_r));
 DFFHQNx3_ASAP7_75t_SL u16_u0_dma_req_r1_reg (.CLK(clk_i),
    .D(n_18871),
    .QN(u16_u0_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u0_dma_req_reg (.CLK(clk_i),
    .D(n_23101),
    .QN(u16_u0_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx3_ASAP7_75t_SL u16_u1_dma_req_r1_reg (.CLK(clk_i),
    .D(n_18875),
    .QN(u16_u1_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u1_dma_req_reg (.CLK(clk_i),
    .D(n_22933),
    .QN(u16_u1_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx3_ASAP7_75t_SL u16_u2_dma_req_r1_reg (.CLK(clk_i),
    .D(n_28881),
    .QN(u16_u2_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u2_dma_req_reg (.CLK(clk_i),
    .D(n_31129),
    .QN(u16_u2_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx2_ASAP7_75t_SL u16_u3_dma_req_r1_reg (.CLK(clk_i),
    .D(n_31740),
    .QN(u16_u3_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u3_dma_req_reg (.CLK(clk_i),
    .D(n_26714),
    .QN(u16_u3_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx3_ASAP7_75t_SL u16_u4_dma_req_r1_reg (.CLK(clk_i),
    .D(n_41611),
    .QN(u16_u4_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u4_dma_req_reg (.CLK(clk_i),
    .D(n_28595),
    .QN(u16_u4_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_L u16_u5_dma_req_r1_reg (.CLK(clk_i),
    .D(n_70201),
    .QN(u16_u5_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u5_dma_req_reg (.CLK(clk_i),
    .D(n_22924),
    .QN(u16_u5_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_L u16_u6_dma_req_r1_reg (.CLK(clk_i),
    .D(n_31272),
    .QN(u16_u6_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u6_dma_req_reg (.CLK(clk_i),
    .D(n_28663),
    .QN(u16_u6_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_L u16_u7_dma_req_r1_reg (.CLK(clk_i),
    .D(n_29938),
    .QN(u16_u7_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u7_dma_req_reg (.CLK(clk_i),
    .D(n_4161),
    .QN(u16_u7_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_L u16_u8_dma_req_r1_reg (.CLK(clk_i),
    .D(n_18872),
    .QN(u16_u8_dma_req_r1));
 DFFASRHQNx1_ASAP7_75t_SL u16_u8_dma_req_reg (.CLK(clk_i),
    .D(n_4162),
    .QN(u16_u8_dma_req_52),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u17_int_set_reg[0]  (.CLK(clk_i),
    .D(n_34536),
    .QN(oc0_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u17_int_set_reg[1]  (.CLK(clk_i),
    .D(n_36072),
    .QN(oc0_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u17_int_set_reg[2]  (.CLK(clk_i),
    .D(n_49143),
    .QN(oc0_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u18_int_set_reg[0]  (.CLK(clk_i),
    .D(n_15023),
    .QN(oc1_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u18_int_set_reg[1]  (.CLK(clk_i),
    .D(n_46640),
    .QN(oc1_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u18_int_set_reg[2]  (.CLK(clk_i),
    .D(n_58735),
    .QN(oc1_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u19_int_set_reg[0]  (.CLK(clk_i),
    .D(n_24536),
    .QN(oc2_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u19_int_set_reg[1]  (.CLK(clk_i),
    .D(n_36100),
    .QN(oc2_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u19_int_set_reg[2]  (.CLK(clk_i),
    .D(n_19623),
    .QN(oc2_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_R u1_sdata_in_r_reg (.CLK(n_434),
    .D(n_107),
    .QN(u1_sdata_in_r));
 DFFHQNx1_ASAP7_75t_R \u1_slt0_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5290),
    .QN(in_slt0[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt0_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5297),
    .QN(in_slt0[12]));
 DFFHQNx1_ASAP7_75t_R \u1_slt0_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5317),
    .QN(in_slt0[15]));
 DFFHQNx1_ASAP7_75t_R \u1_slt0_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5278),
    .QN(in_slt0[9]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5285),
    .QN(in_slt1[10]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5291),
    .QN(in_slt1[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_4207),
    .QN(in_slt1[5]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4533),
    .QN(in_slt1[6]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5221),
    .QN(in_slt1[7]));
 DFFHQNx1_ASAP7_75t_R \u1_slt1_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5272),
    .QN(in_slt1[8]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5286),
    .QN(in_slt2[10]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5288),
    .QN(in_slt2[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5298),
    .QN(in_slt2[12]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5305),
    .QN(in_slt2[13]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5311),
    .QN(in_slt2[14]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5315),
    .QN(in_slt2[15]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5322),
    .QN(in_slt2[16]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5329),
    .QN(in_slt2[17]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5337),
    .QN(in_slt2[18]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5345),
    .QN(in_slt2[19]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_3906),
    .QN(in_slt2[4]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_4156),
    .QN(in_slt2[5]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4534),
    .QN(in_slt2[6]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5222),
    .QN(in_slt2[7]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5271),
    .QN(in_slt2[8]));
 DFFHQNx1_ASAP7_75t_R \u1_slt2_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5277),
    .QN(in_slt2[9]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2275),
    .QN(in_slt3[0]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5281),
    .QN(in_slt3[10]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5289),
    .QN(in_slt3[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5299),
    .QN(in_slt3[12]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5306),
    .QN(in_slt3[13]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5312),
    .QN(in_slt3[14]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5318),
    .QN(in_slt3[15]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5323),
    .QN(in_slt3[16]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5330),
    .QN(in_slt3[17]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5340),
    .QN(in_slt3[18]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5346),
    .QN(in_slt3[19]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_2274),
    .QN(in_slt3[1]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2651),
    .QN(in_slt3[2]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_2948),
    .QN(in_slt3[3]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_3948),
    .QN(in_slt3[4]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_4208),
    .QN(in_slt3[5]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4535),
    .QN(in_slt3[6]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5223),
    .QN(in_slt3[7]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5267),
    .QN(in_slt3[8]));
 DFFHQNx1_ASAP7_75t_R \u1_slt3_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5276),
    .QN(in_slt3[9]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2479),
    .QN(in_slt4[0]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5282),
    .QN(in_slt4[10]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5292),
    .QN(in_slt4[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5300),
    .QN(in_slt4[12]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5307),
    .QN(in_slt4[13]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5310),
    .QN(in_slt4[14]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5319),
    .QN(in_slt4[15]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5324),
    .QN(in_slt4[16]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5328),
    .QN(in_slt4[17]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5343),
    .QN(in_slt4[18]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5347),
    .QN(in_slt4[19]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_2478),
    .QN(in_slt4[1]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2576),
    .QN(in_slt4[2]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_2941),
    .QN(in_slt4[3]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_3947),
    .QN(in_slt4[4]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_4177),
    .QN(in_slt4[5]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4536),
    .QN(in_slt4[6]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5224),
    .QN(in_slt4[7]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5268),
    .QN(in_slt4[8]));
 DFFHQNx1_ASAP7_75t_R \u1_slt4_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5275),
    .QN(in_slt4[9]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2575),
    .QN(in_slt6[0]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5283),
    .QN(in_slt6[10]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5294),
    .QN(in_slt6[11]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5301),
    .QN(in_slt6[12]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5304),
    .QN(in_slt6[13]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5309),
    .QN(in_slt6[14]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5316),
    .QN(in_slt6[15]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5321),
    .QN(in_slt6[16]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5327),
    .QN(in_slt6[17]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5335),
    .QN(in_slt6[18]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5344),
    .QN(in_slt6[19]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_2574),
    .QN(in_slt6[1]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2612),
    .QN(in_slt6[2]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_2940),
    .QN(in_slt6[3]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_3907),
    .QN(in_slt6[4]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_4155),
    .QN(in_slt6[5]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4537),
    .QN(in_slt6[6]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_5225),
    .QN(in_slt6[7]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_5269),
    .QN(in_slt6[8]));
 DFFHQNx1_ASAP7_75t_R \u1_slt6_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5274),
    .QN(in_slt6[9]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_560),
    .QN(u1_sr[0]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[10]  (.CLK(bit_clk_pad_i),
    .D(n_5273),
    .QN(u1_sr[10]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[11]  (.CLK(bit_clk_pad_i),
    .D(n_5280),
    .QN(u1_sr[11]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[12]  (.CLK(bit_clk_pad_i),
    .D(n_5287),
    .QN(u1_sr[12]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[13]  (.CLK(bit_clk_pad_i),
    .D(n_5295),
    .QN(u1_sr[13]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[14]  (.CLK(bit_clk_pad_i),
    .D(n_5302),
    .QN(u1_sr[14]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[15]  (.CLK(bit_clk_pad_i),
    .D(n_5308),
    .QN(u1_sr[15]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[16]  (.CLK(bit_clk_pad_i),
    .D(n_5313),
    .QN(u1_sr[16]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[17]  (.CLK(bit_clk_pad_i),
    .D(n_5320),
    .QN(u1_sr[17]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[18]  (.CLK(bit_clk_pad_i),
    .D(n_5326),
    .QN(u1_sr[18]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[19]  (.CLK(bit_clk_pad_i),
    .D(n_5331),
    .QN(u1_sr[19]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_1231),
    .QN(u1_sr[1]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2136),
    .QN(u1_sr[2]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_2292),
    .QN(u1_sr[3]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_2684),
    .QN(u1_sr[4]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_2974),
    .QN(u1_sr[5]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_4003),
    .QN(u1_sr[6]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_4230),
    .QN(u1_sr[7]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[8]  (.CLK(bit_clk_pad_i),
    .D(n_4624),
    .QN(u1_sr[8]));
 DFFHQNx1_ASAP7_75t_R \u1_sr_reg[9]  (.CLK(bit_clk_pad_i),
    .D(n_5263),
    .QN(u1_sr[9]));
 DFFASRHQNx1_ASAP7_75t_SL \u20_int_set_reg[0]  (.CLK(clk_i),
    .D(n_4280),
    .QN(oc3_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u20_int_set_reg[1]  (.CLK(clk_i),
    .D(n_36099),
    .QN(oc3_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u20_int_set_reg[2]  (.CLK(clk_i),
    .D(n_12226),
    .QN(oc3_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u21_int_set_reg[0]  (.CLK(clk_i),
    .D(n_15040),
    .QN(oc4_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u21_int_set_reg[1]  (.CLK(clk_i),
    .D(n_36091),
    .QN(oc4_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u21_int_set_reg[2]  (.CLK(clk_i),
    .D(n_43078),
    .QN(oc4_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u22_int_set_reg[0]  (.CLK(clk_i),
    .D(n_15054),
    .QN(oc5_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u22_int_set_reg[1]  (.CLK(clk_i),
    .D(n_37460),
    .QN(oc5_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u22_int_set_reg[2]  (.CLK(clk_i),
    .D(n_78934),
    .QN(oc5_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u23_int_set_reg[0]  (.CLK(clk_i),
    .D(n_24532),
    .QN(ic0_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_L \u23_int_set_reg[1]  (.CLK(clk_i),
    .D(n_2564),
    .QN(ic0_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u23_int_set_reg[2]  (.CLK(clk_i),
    .D(n_17401),
    .QN(ic0_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u24_int_set_reg[0]  (.CLK(clk_i),
    .D(n_29939),
    .QN(ic1_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_L \u24_int_set_reg[1]  (.CLK(clk_i),
    .D(n_2566),
    .QN(ic1_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u24_int_set_reg[2]  (.CLK(clk_i),
    .D(n_4077),
    .QN(ic1_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u25_int_set_reg[0]  (.CLK(clk_i),
    .D(n_15034),
    .QN(ic2_int_set[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_L \u25_int_set_reg[1]  (.CLK(clk_i),
    .D(n_2565),
    .QN(ic2_int_set[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u25_int_set_reg[2]  (.CLK(clk_i),
    .D(n_35399),
    .QN(ic2_int_set[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL u26_ac97_rst__reg (.CLK(clk_i),
    .D(n_2955),
    .QN(u26_ac97_rst_104),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_cnt_reg[0]  (.CLK(clk_i),
    .D(n_21865),
    .QN(u26_cnt[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_cnt_reg[1]  (.CLK(clk_i),
    .D(n_24762),
    .QN(u26_cnt[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_cnt_reg[2]  (.CLK(clk_i),
    .D(n_4505),
    .QN(u26_cnt[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[0]  (.CLK(clk_i),
    .D(n_76056),
    .QN(u26_ps_cnt[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[1]  (.CLK(clk_i),
    .D(n_42618),
    .QN(u26_ps_cnt[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[2]  (.CLK(clk_i),
    .D(n_21871),
    .QN(u26_ps_cnt[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[3]  (.CLK(clk_i),
    .D(n_21872),
    .QN(u26_ps_cnt[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[4]  (.CLK(clk_i),
    .D(n_64000),
    .QN(u26_ps_cnt[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u26_ps_cnt_reg[5]  (.CLK(clk_i),
    .D(n_21867),
    .QN(u26_ps_cnt[5]),
    .RESETN(one_),
    .SETN(rst_i));
 SDFHx1_ASAP7_75t_SL u2_bit_clk_e_reg (.CLK(clk_i),
    .QN(u2_bit_clk_e),
    .D(n_806),
    .SE(u2_bit_clk_r1),
    .SI(u2_bit_clk_r));
 DFFHQNx1_ASAP7_75t_R u2_bit_clk_r1_reg (.CLK(clk_i),
    .D(n_806),
    .QN(u2_bit_clk_r1));
 DFFHQNx1_ASAP7_75t_L u2_bit_clk_r_reg (.CLK(clk_i),
    .D(n_434),
    .QN(u2_bit_clk_r));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2289),
    .QN(u2_cnt[0]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_2466),
    .QN(u2_cnt[1]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2291),
    .QN(u2_cnt[2]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_2464),
    .QN(u2_cnt[3]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_2468),
    .QN(u2_cnt[4]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_2331),
    .QN(u2_cnt[5]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[6]  (.CLK(bit_clk_pad_i),
    .D(n_2560),
    .QN(u2_cnt[6]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFASRHQNx1_ASAP7_75t_R \u2_cnt_reg[7]  (.CLK(bit_clk_pad_i),
    .D(n_2567),
    .QN(u2_cnt[7]),
    .RESETN(rst_i),
    .SETN(one_));
 DFFHQNx1_ASAP7_75t_R \u2_in_valid_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2120),
    .QN(in_valid[0]));
 DFFHQNx1_ASAP7_75t_R \u2_in_valid_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_1646),
    .QN(in_valid[1]));
 DFFHQNx1_ASAP7_75t_R \u2_in_valid_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_1904),
    .QN(in_valid[2]));
 DFFHQNx1_ASAP7_75t_R u2_ld_reg (.CLK(bit_clk_pad_i),
    .D(n_1337),
    .QN(ld));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[0]  (.CLK(bit_clk_pad_i),
    .D(n_2129),
    .QN(out_le[0]));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[1]  (.CLK(bit_clk_pad_i),
    .D(n_1194),
    .QN(out_le[1]));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[2]  (.CLK(bit_clk_pad_i),
    .D(n_2223),
    .QN(out_le[2]));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[3]  (.CLK(bit_clk_pad_i),
    .D(n_1089),
    .QN(out_le[3]));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[4]  (.CLK(bit_clk_pad_i),
    .D(n_1510),
    .QN(out_le[4]));
 DFFHQNx1_ASAP7_75t_R \u2_out_le_reg[5]  (.CLK(bit_clk_pad_i),
    .D(n_1915),
    .QN(out_le[5]));
 DFFHQNx2_ASAP7_75t_SL \u2_res_cnt_reg[0]  (.CLK(clk_i),
    .D(n_2251),
    .QN(u2_res_cnt[0]));
 DFFHQNx1_ASAP7_75t_SL \u2_res_cnt_reg[1]  (.CLK(clk_i),
    .D(n_2519),
    .QN(u2_res_cnt[1]));
 DFFHQNx2_ASAP7_75t_SL \u2_res_cnt_reg[2]  (.CLK(clk_i),
    .D(n_2652),
    .QN(u2_res_cnt[2]));
 DFFHQNx2_ASAP7_75t_SL \u2_res_cnt_reg[3]  (.CLK(clk_i),
    .D(n_2817),
    .QN(u2_res_cnt[3]));
 DFFHQNx1_ASAP7_75t_SL u2_suspended_reg (.CLK(clk_i),
    .D(n_19578),
    .QN(u13_csr[1]));
 DFFHQNx1_ASAP7_75t_R u2_sync_beat_reg (.CLK(bit_clk_pad_i),
    .D(n_529),
    .QN(u2_sync_beat));
 DFFASRHQNx1_ASAP7_75t_SL u2_sync_resume_reg (.CLK(clk_i),
    .D(n_2976),
    .QN(u2_sync_resume),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[0]  (.CLK(clk_i),
    .D(n_2302),
    .QN(u2_to_cnt[0]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[1]  (.CLK(clk_i),
    .D(n_17079),
    .QN(u2_to_cnt[1]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[2]  (.CLK(clk_i),
    .D(n_14945),
    .QN(u2_to_cnt[2]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[3]  (.CLK(clk_i),
    .D(n_43469),
    .QN(u2_to_cnt[3]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[4]  (.CLK(clk_i),
    .D(n_17441),
    .QN(u2_to_cnt[4]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFASRHQNx1_ASAP7_75t_SL \u2_to_cnt_reg[5]  (.CLK(clk_i),
    .D(n_2702),
    .QN(u2_to_cnt[5]),
    .RESETN(one_),
    .SETN(rst_i));
 DFFHQNx1_ASAP7_75t_R u2_valid_reg (.CLK(bit_clk_pad_i),
    .D(n_1651),
    .QN(valid));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[0]  (.CLK(clk_i),
    .D(n_14008),
    .QN(out_slt3[0]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[10]  (.CLK(clk_i),
    .D(n_8008),
    .QN(out_slt3[10]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[11]  (.CLK(clk_i),
    .D(n_8006),
    .QN(out_slt3[11]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[12]  (.CLK(clk_i),
    .D(n_4927),
    .QN(out_slt3[12]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[13]  (.CLK(clk_i),
    .D(n_8119),
    .QN(out_slt3[13]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[14]  (.CLK(clk_i),
    .D(n_31865),
    .QN(out_slt3[14]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[15]  (.CLK(clk_i),
    .D(n_31867),
    .QN(out_slt3[15]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[16]  (.CLK(clk_i),
    .D(n_5023),
    .QN(out_slt3[16]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[17]  (.CLK(clk_i),
    .D(n_5022),
    .QN(out_slt3[17]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[18]  (.CLK(clk_i),
    .D(n_5021),
    .QN(out_slt3[18]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[19]  (.CLK(clk_i),
    .D(n_5054),
    .QN(out_slt3[19]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[1]  (.CLK(clk_i),
    .D(n_4516),
    .QN(out_slt3[1]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[2]  (.CLK(clk_i),
    .D(n_24596),
    .QN(out_slt3[2]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[3]  (.CLK(clk_i),
    .D(n_4794),
    .QN(out_slt3[3]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[4]  (.CLK(clk_i),
    .D(n_5036),
    .QN(out_slt3[4]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[5]  (.CLK(clk_i),
    .D(n_14418),
    .QN(out_slt3[5]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[6]  (.CLK(clk_i),
    .D(n_7491),
    .QN(out_slt3[6]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[7]  (.CLK(clk_i),
    .D(n_7527),
    .QN(out_slt3[7]));
 DFFHQNx2_ASAP7_75t_SL \u3_dout_reg[8]  (.CLK(clk_i),
    .D(n_5081),
    .QN(out_slt3[8]));
 DFFHQNx1_ASAP7_75t_SL \u3_dout_reg[9]  (.CLK(clk_i),
    .D(n_5082),
    .QN(out_slt3[9]));
 DFFHQNx1_ASAP7_75t_SL u3_empty_reg (.CLK(clk_i),
    .D(n_75795),
    .QN(o3_empty));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_52913),
    .QN(\u3_mem[0] [0]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_66835),
    .QN(\u3_mem[0] [10]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_52900),
    .QN(\u3_mem[0] [11]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_52926),
    .QN(\u3_mem[0] [12]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_52907),
    .QN(\u3_mem[0] [13]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_52922),
    .QN(\u3_mem[0] [14]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_52920),
    .QN(\u3_mem[0] [15]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_52919),
    .QN(\u3_mem[0] [16]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_52901),
    .QN(\u3_mem[0] [17]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_52915),
    .QN(\u3_mem[0] [18]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_52918),
    .QN(\u3_mem[0] [19]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_52896),
    .QN(\u3_mem[0] [1]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_52905),
    .QN(\u3_mem[0] [20]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_52897),
    .QN(\u3_mem[0] [21]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_66805),
    .QN(\u3_mem[0] [22]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_52921),
    .QN(\u3_mem[0] [23]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_52903),
    .QN(\u3_mem[0] [24]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_52906),
    .QN(\u3_mem[0] [25]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_52912),
    .QN(\u3_mem[0] [26]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_52910),
    .QN(\u3_mem[0] [27]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_52914),
    .QN(\u3_mem[0] [28]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_52917),
    .QN(\u3_mem[0] [29]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_52924),
    .QN(\u3_mem[0] [2]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_52908),
    .QN(\u3_mem[0] [30]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_52916),
    .QN(\u3_mem[0] [31]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_52895),
    .QN(\u3_mem[0] [3]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_68231),
    .QN(\u3_mem[0] [4]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_52923),
    .QN(\u3_mem[0] [5]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_52899),
    .QN(\u3_mem[0] [6]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_52902),
    .QN(\u3_mem[0] [7]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_52909),
    .QN(\u3_mem[0] [8]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_52911),
    .QN(\u3_mem[0] [9]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_15496),
    .QN(\u3_mem[1] [0]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_66825),
    .QN(\u3_mem[1] [10]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_16304),
    .QN(\u3_mem[1] [11]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_15515),
    .QN(\u3_mem[1] [12]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_15473),
    .QN(\u3_mem[1] [13]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_15487),
    .QN(\u3_mem[1] [14]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_16593),
    .QN(\u3_mem[1] [15]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_15481),
    .QN(\u3_mem[1] [16]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_15521),
    .QN(\u3_mem[1] [17]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_15534),
    .QN(\u3_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_16427),
    .QN(\u3_mem[1] [19]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_3621),
    .QN(\u3_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_15145),
    .QN(\u3_mem[1] [20]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_10259),
    .QN(\u3_mem[1] [21]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_66816),
    .QN(\u3_mem[1] [22]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_15775),
    .QN(\u3_mem[1] [23]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_15475),
    .QN(\u3_mem[1] [24]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_16031),
    .QN(\u3_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_15854),
    .QN(\u3_mem[1] [26]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_15771),
    .QN(\u3_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_15773),
    .QN(\u3_mem[1] [28]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_22371),
    .QN(\u3_mem[1] [29]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_16416),
    .QN(\u3_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_22506),
    .QN(\u3_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_15426),
    .QN(\u3_mem[1] [31]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_22578),
    .QN(\u3_mem[1] [3]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_69028),
    .QN(\u3_mem[1] [4]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_15166),
    .QN(\u3_mem[1] [5]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_22311),
    .QN(\u3_mem[1] [6]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_15483),
    .QN(\u3_mem[1] [7]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_15469),
    .QN(\u3_mem[1] [8]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_15506),
    .QN(\u3_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_24812),
    .QN(\u3_mem[2] [0]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_24824),
    .QN(\u3_mem[2] [10]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_24821),
    .QN(\u3_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_24820),
    .QN(\u3_mem[2] [12]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_24830),
    .QN(\u3_mem[2] [13]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_24816),
    .QN(\u3_mem[2] [14]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_24811),
    .QN(\u3_mem[2] [15]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_24825),
    .QN(\u3_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_24815),
    .QN(\u3_mem[2] [17]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_24826),
    .QN(\u3_mem[2] [18]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_24813),
    .QN(\u3_mem[2] [19]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_24819),
    .QN(\u3_mem[2] [1]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_24814),
    .QN(\u3_mem[2] [20]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_24833),
    .QN(\u3_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_66812),
    .QN(\u3_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_24810),
    .QN(\u3_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_24809),
    .QN(\u3_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_24808),
    .QN(\u3_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_24838),
    .QN(\u3_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_24835),
    .QN(\u3_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_24807),
    .QN(\u3_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_24837),
    .QN(\u3_mem[2] [29]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_24822),
    .QN(\u3_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_24828),
    .QN(\u3_mem[2] [30]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_24827),
    .QN(\u3_mem[2] [31]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_24818),
    .QN(\u3_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_68219),
    .QN(\u3_mem[2] [4]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_24823),
    .QN(\u3_mem[2] [5]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_24831),
    .QN(\u3_mem[2] [6]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_24817),
    .QN(\u3_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_24829),
    .QN(\u3_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_24832),
    .QN(\u3_mem[2] [9]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_13094),
    .QN(\u3_mem[3] [0]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_13085),
    .QN(\u3_mem[3] [10]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_13084),
    .QN(\u3_mem[3] [11]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_13083),
    .QN(\u3_mem[3] [12]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_13082),
    .QN(\u3_mem[3] [13]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_13081),
    .QN(\u3_mem[3] [14]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_13080),
    .QN(\u3_mem[3] [15]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_13079),
    .QN(\u3_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_48431),
    .QN(\u3_mem[3] [17]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_13077),
    .QN(\u3_mem[3] [18]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_13076),
    .QN(\u3_mem[3] [19]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_13095),
    .QN(\u3_mem[3] [1]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_13075),
    .QN(\u3_mem[3] [20]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_48434),
    .QN(\u3_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_13072),
    .QN(\u3_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_13069),
    .QN(\u3_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_13066),
    .QN(\u3_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_13065),
    .QN(\u3_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_13064),
    .QN(\u3_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_13063),
    .QN(\u3_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_13067),
    .QN(\u3_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_13071),
    .QN(\u3_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_13093),
    .QN(\u3_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_13070),
    .QN(\u3_mem[3] [30]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_13068),
    .QN(\u3_mem[3] [31]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_13092),
    .QN(\u3_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_69027),
    .QN(\u3_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_13090),
    .QN(\u3_mem[3] [5]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_13089),
    .QN(\u3_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_13088),
    .QN(\u3_mem[3] [7]));
 DFFHQNx1_ASAP7_75t_SL \u3_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_13087),
    .QN(\u3_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u3_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_13086),
    .QN(\u3_mem[3] [9]));
 SDFHx4_ASAP7_75t_SL \u3_rp_reg[0]  (.CLK(clk_i),
    .D(n_29312),
    .QN(u3_rp[0]),
    .SE(u3_rp[0]),
    .SI(n_21234));
 DFFHQx4_ASAP7_75t_SL \u3_rp_reg[1]  (.CLK(clk_i),
    .D(n_27237),
    .Q(u3_rp[1]));
 DFFHQx4_ASAP7_75t_SL \u3_rp_reg[2]  (.CLK(clk_i),
    .D(n_29313),
    .Q(u3_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u3_rp_reg[3]  (.CLK(clk_i),
    .D(n_21795),
    .QN(u3_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u3_status_reg[0]  (.CLK(clk_i),
    .D(n_40420),
    .QN(o3_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u3_status_reg[1]  (.CLK(clk_i),
    .D(n_5847),
    .QN(o3_status[1]));
 DFFHQx4_ASAP7_75t_SL \u3_wp_reg[0]  (.CLK(clk_i),
    .D(n_2983),
    .Q(u3_wp[0]));
 DFFHQNx1_ASAP7_75t_SL \u3_wp_reg[1]  (.CLK(clk_i),
    .D(n_3913),
    .QN(u3_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u3_wp_reg[2]  (.CLK(clk_i),
    .D(n_3081),
    .QN(u3_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[0]  (.CLK(clk_i),
    .D(n_43096),
    .QN(out_slt4[0]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[10]  (.CLK(clk_i),
    .D(n_64856),
    .QN(out_slt4[10]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[11]  (.CLK(clk_i),
    .D(n_32587),
    .QN(out_slt4[11]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[12]  (.CLK(clk_i),
    .D(n_32588),
    .QN(out_slt4[12]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[13]  (.CLK(clk_i),
    .D(n_32597),
    .QN(out_slt4[13]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[14]  (.CLK(clk_i),
    .D(n_32599),
    .QN(out_slt4[14]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[15]  (.CLK(clk_i),
    .D(n_32595),
    .QN(out_slt4[15]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[16]  (.CLK(clk_i),
    .D(n_32593),
    .QN(out_slt4[16]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[17]  (.CLK(clk_i),
    .D(n_32589),
    .QN(out_slt4[17]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[18]  (.CLK(clk_i),
    .D(n_34634),
    .QN(out_slt4[18]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[19]  (.CLK(clk_i),
    .D(n_32601),
    .QN(out_slt4[19]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[1]  (.CLK(clk_i),
    .D(n_43092),
    .QN(out_slt4[1]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[2]  (.CLK(clk_i),
    .D(n_43095),
    .QN(out_slt4[2]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[3]  (.CLK(clk_i),
    .D(n_43094),
    .QN(out_slt4[3]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[4]  (.CLK(clk_i),
    .D(n_32600),
    .QN(out_slt4[4]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[5]  (.CLK(clk_i),
    .D(n_52934),
    .QN(out_slt4[5]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[6]  (.CLK(clk_i),
    .D(n_32592),
    .QN(out_slt4[6]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[7]  (.CLK(clk_i),
    .D(n_32591),
    .QN(out_slt4[7]));
 DFFHQNx1_ASAP7_75t_SL \u4_dout_reg[8]  (.CLK(clk_i),
    .D(n_32590),
    .QN(out_slt4[8]));
 DFFHQNx2_ASAP7_75t_SL \u4_dout_reg[9]  (.CLK(clk_i),
    .D(n_32584),
    .QN(out_slt4[9]));
 DFFHQNx1_ASAP7_75t_SL u4_empty_reg (.CLK(clk_i),
    .D(n_65329),
    .QN(o4_empty));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_33684),
    .QN(\u4_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_66832),
    .QN(\u4_mem[0] [10]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_33667),
    .QN(\u4_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_33666),
    .QN(\u4_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_33659),
    .QN(\u4_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_33661),
    .QN(\u4_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_33673),
    .QN(\u4_mem[0] [15]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_33665),
    .QN(\u4_mem[0] [16]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_33664),
    .QN(\u4_mem[0] [17]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_33658),
    .QN(\u4_mem[0] [18]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_33682),
    .QN(\u4_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_33685),
    .QN(\u4_mem[0] [1]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_33663),
    .QN(\u4_mem[0] [20]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_33681),
    .QN(\u4_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_66815),
    .QN(\u4_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_33662),
    .QN(\u4_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_33656),
    .QN(\u4_mem[0] [24]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_33677),
    .QN(\u4_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_33676),
    .QN(\u4_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_33675),
    .QN(\u4_mem[0] [27]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_33678),
    .QN(\u4_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_33686),
    .QN(\u4_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_33660),
    .QN(\u4_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_33674),
    .QN(\u4_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_33679),
    .QN(\u4_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_33671),
    .QN(\u4_mem[0] [3]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_69015),
    .QN(\u4_mem[0] [4]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_33683),
    .QN(\u4_mem[0] [5]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_33687),
    .QN(\u4_mem[0] [6]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_33672),
    .QN(\u4_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_33670),
    .QN(\u4_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_33668),
    .QN(\u4_mem[0] [9]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_65251),
    .QN(\u4_mem[1] [0]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_65764),
    .QN(\u4_mem[1] [10]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_65255),
    .QN(\u4_mem[1] [11]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_65263),
    .QN(\u4_mem[1] [12]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_65244),
    .QN(\u4_mem[1] [13]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_65247),
    .QN(\u4_mem[1] [14]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_65268),
    .QN(\u4_mem[1] [15]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_65256),
    .QN(\u4_mem[1] [16]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_65257),
    .QN(\u4_mem[1] [17]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_65252),
    .QN(\u4_mem[1] [18]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_65258),
    .QN(\u4_mem[1] [19]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_65269),
    .QN(\u4_mem[1] [1]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_65250),
    .QN(\u4_mem[1] [20]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_65249),
    .QN(\u4_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_65267),
    .QN(\u4_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_65243),
    .QN(\u4_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_65242),
    .QN(\u4_mem[1] [24]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_65248),
    .QN(\u4_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_65238),
    .QN(\u4_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_65240),
    .QN(\u4_mem[1] [27]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_65260),
    .QN(\u4_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_65270),
    .QN(\u4_mem[1] [29]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_65246),
    .QN(\u4_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_65253),
    .QN(\u4_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_65241),
    .QN(\u4_mem[1] [31]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_65245),
    .QN(\u4_mem[1] [3]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_69024),
    .QN(\u4_mem[1] [4]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_65265),
    .QN(\u4_mem[1] [5]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_65261),
    .QN(\u4_mem[1] [6]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_65262),
    .QN(\u4_mem[1] [7]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_65254),
    .QN(\u4_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_65266),
    .QN(\u4_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_10918),
    .QN(\u4_mem[2] [0]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_66827),
    .QN(\u4_mem[2] [10]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_10018),
    .QN(\u4_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_10047),
    .QN(\u4_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_10104),
    .QN(\u4_mem[2] [13]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_9756),
    .QN(\u4_mem[2] [14]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_9785),
    .QN(\u4_mem[2] [15]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_10133),
    .QN(\u4_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_10161),
    .QN(\u4_mem[2] [17]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_10187),
    .QN(\u4_mem[2] [18]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_10214),
    .QN(\u4_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_10896),
    .QN(\u4_mem[2] [1]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_10241),
    .QN(\u4_mem[2] [20]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_10268),
    .QN(\u4_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_66810),
    .QN(\u4_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_10324),
    .QN(\u4_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_10430),
    .QN(\u4_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_10456),
    .QN(\u4_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_10482),
    .QN(\u4_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_10507),
    .QN(\u4_mem[2] [27]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_10378),
    .QN(\u4_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_10681),
    .QN(\u4_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_9844),
    .QN(\u4_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_10657),
    .QN(\u4_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_10351),
    .QN(\u4_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_9874),
    .QN(\u4_mem[2] [3]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_69023),
    .QN(\u4_mem[2] [4]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_10076),
    .QN(\u4_mem[2] [5]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_9727),
    .QN(\u4_mem[2] [6]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_9815),
    .QN(\u4_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_9903),
    .QN(\u4_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_9958),
    .QN(\u4_mem[2] [9]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_3933),
    .QN(\u4_mem[3] [0]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_30254),
    .QN(\u4_mem[3] [10]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_3703),
    .QN(\u4_mem[3] [11]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_3702),
    .QN(\u4_mem[3] [12]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_3701),
    .QN(\u4_mem[3] [13]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_3700),
    .QN(\u4_mem[3] [14]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_3699),
    .QN(\u4_mem[3] [15]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_3698),
    .QN(\u4_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_3697),
    .QN(\u4_mem[3] [17]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_11191),
    .QN(\u4_mem[3] [18]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_11190),
    .QN(\u4_mem[3] [19]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_3934),
    .QN(\u4_mem[3] [1]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_47334),
    .QN(\u4_mem[3] [20]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_11188),
    .QN(\u4_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_11187),
    .QN(\u4_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_11186),
    .QN(\u4_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_11185),
    .QN(\u4_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_11184),
    .QN(\u4_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_11183),
    .QN(\u4_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_26054),
    .QN(\u4_mem[3] [27]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_26057),
    .QN(\u4_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_30247),
    .QN(\u4_mem[3] [29]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_3935),
    .QN(\u4_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_30235),
    .QN(\u4_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_26055),
    .QN(\u4_mem[3] [31]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_3941),
    .QN(\u4_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_69022),
    .QN(\u4_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_47322),
    .QN(\u4_mem[3] [5]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_47255),
    .QN(\u4_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_47391),
    .QN(\u4_mem[3] [7]));
 DFFHQNx1_ASAP7_75t_SL \u4_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_3955),
    .QN(\u4_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u4_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_3956),
    .QN(\u4_mem[3] [9]));
 SDFHx4_ASAP7_75t_SL \u4_rp_reg[0]  (.CLK(clk_i),
    .D(n_43097),
    .QN(u4_rp[0]),
    .SE(n_71390),
    .SI(n_24641));
 DFFHQx4_ASAP7_75t_SL \u4_rp_reg[1]  (.CLK(clk_i),
    .D(n_50602),
    .Q(u4_rp[1]));
 DFFHQNx2_ASAP7_75t_SL \u4_rp_reg[2]  (.CLK(clk_i),
    .D(n_43091),
    .QN(u4_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u4_rp_reg[3]  (.CLK(clk_i),
    .D(n_22829),
    .QN(u4_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u4_status_reg[0]  (.CLK(clk_i),
    .D(n_71393),
    .QN(o4_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u4_status_reg[1]  (.CLK(clk_i),
    .D(n_5846),
    .QN(o4_status[1]));
 DFFHQx4_ASAP7_75t_SL \u4_wp_reg[0]  (.CLK(clk_i),
    .D(n_2985),
    .Q(u4_wp[0]));
 DFFHQNx1_ASAP7_75t_SL \u4_wp_reg[1]  (.CLK(clk_i),
    .D(n_29662),
    .QN(u4_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u4_wp_reg[2]  (.CLK(clk_i),
    .D(n_41379),
    .QN(u4_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[0]  (.CLK(clk_i),
    .D(n_66683),
    .QN(out_slt6[0]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[10]  (.CLK(clk_i),
    .D(n_43761),
    .QN(out_slt6[10]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[11]  (.CLK(clk_i),
    .D(n_23394),
    .QN(out_slt6[11]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[12]  (.CLK(clk_i),
    .D(n_7251),
    .QN(out_slt6[12]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[13]  (.CLK(clk_i),
    .D(n_7997),
    .QN(out_slt6[13]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[14]  (.CLK(clk_i),
    .D(n_7942),
    .QN(out_slt6[14]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[15]  (.CLK(clk_i),
    .D(n_47683),
    .QN(out_slt6[15]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[16]  (.CLK(clk_i),
    .D(n_29630),
    .QN(out_slt6[16]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[17]  (.CLK(clk_i),
    .D(n_17304),
    .QN(out_slt6[17]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[18]  (.CLK(clk_i),
    .D(n_73174),
    .QN(out_slt6[18]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[19]  (.CLK(clk_i),
    .D(n_66663),
    .QN(out_slt6[19]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[1]  (.CLK(clk_i),
    .D(n_66681),
    .QN(out_slt6[1]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[2]  (.CLK(clk_i),
    .D(n_66665),
    .QN(out_slt6[2]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[3]  (.CLK(clk_i),
    .D(n_66679),
    .QN(out_slt6[3]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[4]  (.CLK(clk_i),
    .D(n_52940),
    .QN(out_slt6[4]));
 DFFHQNx1_ASAP7_75t_SL \u5_dout_reg[5]  (.CLK(clk_i),
    .D(n_54566),
    .QN(out_slt6[5]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[6]  (.CLK(clk_i),
    .D(n_7288),
    .QN(out_slt6[6]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[7]  (.CLK(clk_i),
    .D(n_7308),
    .QN(out_slt6[7]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[8]  (.CLK(clk_i),
    .D(n_8013),
    .QN(out_slt6[8]));
 DFFHQNx2_ASAP7_75t_SL \u5_dout_reg[9]  (.CLK(clk_i),
    .D(n_7995),
    .QN(out_slt6[9]));
 DFFHQNx1_ASAP7_75t_SL u5_empty_reg (.CLK(clk_i),
    .D(n_23154),
    .QN(o6_empty));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_26419),
    .QN(\u5_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_26399),
    .QN(\u5_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_26404),
    .QN(\u5_mem[0] [11]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_26409),
    .QN(\u5_mem[0] [12]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_26395),
    .QN(\u5_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_26417),
    .QN(\u5_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_26416),
    .QN(\u5_mem[0] [15]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_26394),
    .QN(\u5_mem[0] [16]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_26393),
    .QN(\u5_mem[0] [17]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_26392),
    .QN(\u5_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_26391),
    .QN(\u5_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_26418),
    .QN(\u5_mem[0] [1]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_26415),
    .QN(\u5_mem[0] [20]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_26411),
    .QN(\u5_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_26405),
    .QN(\u5_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_26407),
    .QN(\u5_mem[0] [23]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_26412),
    .QN(\u5_mem[0] [24]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_26408),
    .QN(\u5_mem[0] [25]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_26414),
    .QN(\u5_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_26406),
    .QN(\u5_mem[0] [27]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_26413),
    .QN(\u5_mem[0] [28]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_26387),
    .QN(\u5_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_26410),
    .QN(\u5_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_26388),
    .QN(\u5_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_26390),
    .QN(\u5_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_26401),
    .QN(\u5_mem[0] [3]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_69019),
    .QN(\u5_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_26396),
    .QN(\u5_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_26403),
    .QN(\u5_mem[0] [6]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_26402),
    .QN(\u5_mem[0] [7]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_26400),
    .QN(\u5_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_26398),
    .QN(\u5_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_3638),
    .QN(\u5_mem[1] [0]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_66819),
    .QN(\u5_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_10007),
    .QN(\u5_mem[1] [11]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_10036),
    .QN(\u5_mem[1] [12]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_10094),
    .QN(\u5_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_9745),
    .QN(\u5_mem[1] [14]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_9774),
    .QN(\u5_mem[1] [15]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_10122),
    .QN(\u5_mem[1] [16]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_10151),
    .QN(\u5_mem[1] [17]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_10177),
    .QN(\u5_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_10204),
    .QN(\u5_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_3635),
    .QN(\u5_mem[1] [1]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_10231),
    .QN(\u5_mem[1] [20]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_10260),
    .QN(\u5_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_66807),
    .QN(\u5_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_10315),
    .QN(\u5_mem[1] [23]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_10420),
    .QN(\u5_mem[1] [24]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_10446),
    .QN(\u5_mem[1] [25]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_10471),
    .QN(\u5_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_10497),
    .QN(\u5_mem[1] [27]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_10370),
    .QN(\u5_mem[1] [28]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_10670),
    .QN(\u5_mem[1] [29]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_9834),
    .QN(\u5_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_10651),
    .QN(\u5_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_10344),
    .QN(\u5_mem[1] [31]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_9863),
    .QN(\u5_mem[1] [3]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_69020),
    .QN(\u5_mem[1] [4]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_10065),
    .QN(\u5_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_9717),
    .QN(\u5_mem[1] [6]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_9804),
    .QN(\u5_mem[1] [7]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_9892),
    .QN(\u5_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_9949),
    .QN(\u5_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_10921),
    .QN(\u5_mem[2] [0]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_66826),
    .QN(\u5_mem[2] [10]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_10014),
    .QN(\u5_mem[2] [11]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_10043),
    .QN(\u5_mem[2] [12]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_10100),
    .QN(\u5_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_9752),
    .QN(\u5_mem[2] [14]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_9781),
    .QN(\u5_mem[2] [15]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_10129),
    .QN(\u5_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_10157),
    .QN(\u5_mem[2] [17]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_10183),
    .QN(\u5_mem[2] [18]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_10210),
    .QN(\u5_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_10894),
    .QN(\u5_mem[2] [1]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_10238),
    .QN(\u5_mem[2] [20]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_10265),
    .QN(\u5_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_10292),
    .QN(\u5_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_10321),
    .QN(\u5_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_10426),
    .QN(\u5_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_10452),
    .QN(\u5_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_10477),
    .QN(\u5_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_10503),
    .QN(\u5_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_10376),
    .QN(\u5_mem[2] [28]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_10679),
    .QN(\u5_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_9841),
    .QN(\u5_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_10641),
    .QN(\u5_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_10335),
    .QN(\u5_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_9870),
    .QN(\u5_mem[2] [3]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_69021),
    .QN(\u5_mem[2] [4]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_10072),
    .QN(\u5_mem[2] [5]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_9723),
    .QN(\u5_mem[2] [6]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_9811),
    .QN(\u5_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_9899),
    .QN(\u5_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_9960),
    .QN(\u5_mem[2] [9]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_3862),
    .QN(\u5_mem[3] [0]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_9914),
    .QN(\u5_mem[3] [10]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_10001),
    .QN(\u5_mem[3] [11]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_10030),
    .QN(\u5_mem[3] [12]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_10089),
    .QN(\u5_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_9738),
    .QN(\u5_mem[3] [14]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_9767),
    .QN(\u5_mem[3] [15]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_11129),
    .QN(\u5_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_11127),
    .QN(\u5_mem[3] [17]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_11144),
    .QN(\u5_mem[3] [18]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_11143),
    .QN(\u5_mem[3] [19]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_3858),
    .QN(\u5_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_11142),
    .QN(\u5_mem[3] [20]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_11141),
    .QN(\u5_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_11140),
    .QN(\u5_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_11139),
    .QN(\u5_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_11138),
    .QN(\u5_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_11137),
    .QN(\u5_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_11136),
    .QN(\u5_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_3959),
    .QN(\u5_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_11134),
    .QN(\u5_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_11133),
    .QN(\u5_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_9828),
    .QN(\u5_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_11132),
    .QN(\u5_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_11131),
    .QN(\u5_mem[3] [31]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_9857),
    .QN(\u5_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_68229),
    .QN(\u5_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_10061),
    .QN(\u5_mem[3] [5]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_9711),
    .QN(\u5_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_9800),
    .QN(\u5_mem[3] [7]));
 DFFHQNx1_ASAP7_75t_SL \u5_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_9886),
    .QN(\u5_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u5_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_9944),
    .QN(\u5_mem[3] [9]));
 SDFHx4_ASAP7_75t_SL \u5_rp_reg[0]  (.CLK(clk_i),
    .D(n_66675),
    .QN(u5_rp[0]),
    .SE(n_13405),
    .SI(n_58650));
 DFFHQx4_ASAP7_75t_SL \u5_rp_reg[1]  (.CLK(clk_i),
    .D(n_22532),
    .Q(u5_rp[1]));
 DFFHQx4_ASAP7_75t_SL \u5_rp_reg[2]  (.CLK(clk_i),
    .D(n_64851),
    .Q(u5_rp[2]));
 DFFHQNx2_ASAP7_75t_SL \u5_rp_reg[3]  (.CLK(clk_i),
    .D(n_66661),
    .QN(u5_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u5_status_reg[0]  (.CLK(clk_i),
    .D(n_19620),
    .QN(o6_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u5_status_reg[1]  (.CLK(clk_i),
    .D(n_5848),
    .QN(o6_status[1]));
 DFFHQx4_ASAP7_75t_SL \u5_wp_reg[0]  (.CLK(clk_i),
    .D(n_41761),
    .Q(u5_wp[0]));
 DFFHQNx1_ASAP7_75t_SL \u5_wp_reg[1]  (.CLK(clk_i),
    .D(n_17575),
    .QN(u5_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u5_wp_reg[2]  (.CLK(clk_i),
    .D(n_11130),
    .QN(u5_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[0]  (.CLK(clk_i),
    .D(n_46188),
    .QN(out_slt7[0]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[10]  (.CLK(clk_i),
    .D(n_36366),
    .QN(out_slt7[10]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[11]  (.CLK(clk_i),
    .D(n_36367),
    .QN(out_slt7[11]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[12]  (.CLK(clk_i),
    .D(n_25961),
    .QN(out_slt7[12]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[13]  (.CLK(clk_i),
    .D(n_79168),
    .QN(out_slt7[13]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[14]  (.CLK(clk_i),
    .D(n_30357),
    .QN(out_slt7[14]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[15]  (.CLK(clk_i),
    .D(n_29948),
    .QN(out_slt7[15]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[16]  (.CLK(clk_i),
    .D(n_25967),
    .QN(out_slt7[16]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[17]  (.CLK(clk_i),
    .D(n_43291),
    .QN(out_slt7[17]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[18]  (.CLK(clk_i),
    .D(n_25965),
    .QN(out_slt7[18]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[19]  (.CLK(clk_i),
    .D(n_48225),
    .QN(out_slt7[19]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[1]  (.CLK(clk_i),
    .D(n_46191),
    .QN(out_slt7[1]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[2]  (.CLK(clk_i),
    .D(n_13976),
    .QN(out_slt7[2]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[3]  (.CLK(clk_i),
    .D(n_27132),
    .QN(out_slt7[3]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[4]  (.CLK(clk_i),
    .D(n_26103),
    .QN(out_slt7[4]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[5]  (.CLK(clk_i),
    .D(n_25964),
    .QN(out_slt7[5]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[6]  (.CLK(clk_i),
    .D(n_29970),
    .QN(out_slt7[6]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[7]  (.CLK(clk_i),
    .D(n_29949),
    .QN(out_slt7[7]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[8]  (.CLK(clk_i),
    .D(n_25955),
    .QN(out_slt7[8]));
 DFFHQNx2_ASAP7_75t_SL \u6_dout_reg[9]  (.CLK(clk_i),
    .D(n_37141),
    .QN(out_slt7[9]));
 DFFHQNx1_ASAP7_75t_SL u6_empty_reg (.CLK(clk_i),
    .D(n_18668),
    .QN(o7_empty));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_10929),
    .QN(\u6_mem[0] [0]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_66828),
    .QN(\u6_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_10005),
    .QN(\u6_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_10034),
    .QN(\u6_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_10092),
    .QN(\u6_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_9742),
    .QN(\u6_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_9772),
    .QN(\u6_mem[0] [15]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_10119),
    .QN(\u6_mem[0] [16]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_10146),
    .QN(\u6_mem[0] [17]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_10175),
    .QN(\u6_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_10202),
    .QN(\u6_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_10902),
    .QN(\u6_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_10230),
    .QN(\u6_mem[0] [20]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_10257),
    .QN(\u6_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_66803),
    .QN(\u6_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_10310),
    .QN(\u6_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_10414),
    .QN(\u6_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_10442),
    .QN(\u6_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_10467),
    .QN(\u6_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_10493),
    .QN(\u6_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_10366),
    .QN(\u6_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_10669),
    .QN(\u6_mem[0] [29]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_9832),
    .QN(\u6_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_10649),
    .QN(\u6_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_10339),
    .QN(\u6_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_9860),
    .QN(\u6_mem[0] [3]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_69018),
    .QN(\u6_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_10057),
    .QN(\u6_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_9713),
    .QN(\u6_mem[0] [6]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_9802),
    .QN(\u6_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_9889),
    .QN(\u6_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_9941),
    .QN(\u6_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_14390),
    .QN(\u6_mem[1] [0]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_9922),
    .QN(\u6_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_10009),
    .QN(\u6_mem[1] [11]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_10038),
    .QN(\u6_mem[1] [12]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_14399),
    .QN(\u6_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_9747),
    .QN(\u6_mem[1] [14]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_9776),
    .QN(\u6_mem[1] [15]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_10124),
    .QN(\u6_mem[1] [16]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_14400),
    .QN(\u6_mem[1] [17]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_14401),
    .QN(\u6_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_14402),
    .QN(\u6_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_14405),
    .QN(\u6_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_10234),
    .QN(\u6_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_14403),
    .QN(\u6_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_10288),
    .QN(\u6_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_10317),
    .QN(\u6_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_10422),
    .QN(\u6_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_78411),
    .QN(\u6_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_10473),
    .QN(\u6_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_10499),
    .QN(\u6_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_10372),
    .QN(\u6_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_10676),
    .QN(\u6_mem[1] [29]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_14393),
    .QN(\u6_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_10654),
    .QN(\u6_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_10346),
    .QN(\u6_mem[1] [31]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_14394),
    .QN(\u6_mem[1] [3]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_68211),
    .QN(\u6_mem[1] [4]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_14398),
    .QN(\u6_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_14391),
    .QN(\u6_mem[1] [6]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_14392),
    .QN(\u6_mem[1] [7]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_14395),
    .QN(\u6_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_14396),
    .QN(\u6_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_70056),
    .QN(\u6_mem[2] [0]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_70057),
    .QN(\u6_mem[2] [10]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_70070),
    .QN(\u6_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_70066),
    .QN(\u6_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_70068),
    .QN(\u6_mem[2] [13]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_70043),
    .QN(\u6_mem[2] [14]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_70054),
    .QN(\u6_mem[2] [15]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_70060),
    .QN(\u6_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_70071),
    .QN(\u6_mem[2] [17]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_70042),
    .QN(\u6_mem[2] [18]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_70055),
    .QN(\u6_mem[2] [19]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_78045),
    .QN(\u6_mem[2] [1]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_70053),
    .QN(\u6_mem[2] [20]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_70051),
    .QN(\u6_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_70072),
    .QN(\u6_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_70044),
    .QN(\u6_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_70052),
    .QN(\u6_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_70048),
    .QN(\u6_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_70064),
    .QN(\u6_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_70047),
    .QN(\u6_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_70045),
    .QN(\u6_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_70063),
    .QN(\u6_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_70058),
    .QN(\u6_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_70050),
    .QN(\u6_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_70067),
    .QN(\u6_mem[2] [31]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_70062),
    .QN(\u6_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_70040),
    .QN(\u6_mem[2] [4]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_70046),
    .QN(\u6_mem[2] [5]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_70065),
    .QN(\u6_mem[2] [6]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_70069),
    .QN(\u6_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_70059),
    .QN(\u6_mem[2] [8]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_70061),
    .QN(\u6_mem[2] [9]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_44456),
    .QN(\u6_mem[3] [0]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_66821),
    .QN(\u6_mem[3] [10]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_44440),
    .QN(\u6_mem[3] [11]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_77234),
    .QN(\u6_mem[3] [12]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_49641),
    .QN(\u6_mem[3] [13]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_60588),
    .QN(\u6_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_46422),
    .QN(\u6_mem[3] [15]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_22315),
    .QN(\u6_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_25333),
    .QN(\u6_mem[3] [17]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_25332),
    .QN(\u6_mem[3] [18]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_25331),
    .QN(\u6_mem[3] [19]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_11295),
    .QN(\u6_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_25330),
    .QN(\u6_mem[3] [20]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_29355),
    .QN(\u6_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_29356),
    .QN(\u6_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_29358),
    .QN(\u6_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_47164),
    .QN(\u6_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_47127),
    .QN(\u6_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_19241),
    .QN(\u6_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_64862),
    .QN(\u6_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_22642),
    .QN(\u6_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_19234),
    .QN(\u6_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_76778),
    .QN(\u6_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_19235),
    .QN(\u6_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_19237),
    .QN(\u6_mem[3] [31]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_45388),
    .QN(\u6_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_69013),
    .QN(\u6_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_44452),
    .QN(\u6_mem[3] [5]));
 DFFHQNx2_ASAP7_75t_SL \u6_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_76986),
    .QN(\u6_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_61229),
    .QN(\u6_mem[3] [7]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_44447),
    .QN(\u6_mem[3] [8]));
 DFFHQNx1_ASAP7_75t_SL \u6_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_44864),
    .QN(\u6_mem[3] [9]));
 SDFHx4_ASAP7_75t_SL \u6_rp_reg[0]  (.CLK(clk_i),
    .D(n_4645),
    .QN(u6_rp[0]),
    .SE(u6_rp[0]),
    .SI(n_4312));
 DFFHQx4_ASAP7_75t_SL \u6_rp_reg[1]  (.CLK(clk_i),
    .D(n_12099),
    .Q(u6_rp[1]));
 DFFHQx4_ASAP7_75t_SL \u6_rp_reg[2]  (.CLK(clk_i),
    .D(n_4646),
    .Q(u6_rp[2]));
 DFFHQNx2_ASAP7_75t_SL \u6_rp_reg[3]  (.CLK(clk_i),
    .D(n_28111),
    .QN(u6_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u6_status_reg[0]  (.CLK(clk_i),
    .D(n_12225),
    .QN(o7_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u6_status_reg[1]  (.CLK(clk_i),
    .D(n_5845),
    .QN(o7_status[1]));
 DFFHQx4_ASAP7_75t_SL \u6_wp_reg[0]  (.CLK(clk_i),
    .D(n_57966),
    .Q(u6_wp[0]));
 DFFHQNx1_ASAP7_75t_SL \u6_wp_reg[1]  (.CLK(clk_i),
    .D(n_28529),
    .QN(u6_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u6_wp_reg[2]  (.CLK(clk_i),
    .D(n_72087),
    .QN(u6_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[0]  (.CLK(clk_i),
    .D(n_42260),
    .QN(out_slt8[0]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[10]  (.CLK(clk_i),
    .D(n_5073),
    .QN(out_slt8[10]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[11]  (.CLK(clk_i),
    .D(n_5074),
    .QN(out_slt8[11]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[12]  (.CLK(clk_i),
    .D(n_17254),
    .QN(out_slt8[12]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[13]  (.CLK(clk_i),
    .D(n_46567),
    .QN(out_slt8[13]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[14]  (.CLK(clk_i),
    .D(n_17110),
    .QN(out_slt8[14]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[15]  (.CLK(clk_i),
    .D(n_22257),
    .QN(out_slt8[15]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[16]  (.CLK(clk_i),
    .D(n_4933),
    .QN(out_slt8[16]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[17]  (.CLK(clk_i),
    .D(n_62718),
    .QN(out_slt8[17]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[18]  (.CLK(clk_i),
    .D(n_42263),
    .QN(out_slt8[18]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[19]  (.CLK(clk_i),
    .D(n_27373),
    .QN(out_slt8[19]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[1]  (.CLK(clk_i),
    .D(n_56869),
    .QN(out_slt8[1]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[2]  (.CLK(clk_i),
    .D(n_19688),
    .QN(out_slt8[2]));
 DFFHQNx1_ASAP7_75t_SL \u7_dout_reg[3]  (.CLK(clk_i),
    .D(n_56870),
    .QN(out_slt8[3]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[4]  (.CLK(clk_i),
    .D(n_5041),
    .QN(out_slt8[4]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[5]  (.CLK(clk_i),
    .D(n_42262),
    .QN(out_slt8[5]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[6]  (.CLK(clk_i),
    .D(n_42261),
    .QN(out_slt8[6]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[7]  (.CLK(clk_i),
    .D(n_42264),
    .QN(out_slt8[7]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[8]  (.CLK(clk_i),
    .D(n_5071),
    .QN(out_slt8[8]));
 DFFHQNx2_ASAP7_75t_SL \u7_dout_reg[9]  (.CLK(clk_i),
    .D(n_5072),
    .QN(out_slt8[9]));
 DFFHQNx1_ASAP7_75t_SL u7_empty_reg (.CLK(clk_i),
    .D(n_18660),
    .QN(o8_empty));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_12404),
    .QN(\u7_mem[0] [0]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_66829),
    .QN(\u7_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_12429),
    .QN(\u7_mem[0] [11]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_12428),
    .QN(\u7_mem[0] [12]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_12414),
    .QN(\u7_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_12419),
    .QN(\u7_mem[0] [14]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_12418),
    .QN(\u7_mem[0] [15]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_12413),
    .QN(\u7_mem[0] [16]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_12412),
    .QN(\u7_mem[0] [17]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_12411),
    .QN(\u7_mem[0] [18]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_12410),
    .QN(\u7_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_12405),
    .QN(\u7_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_12427),
    .QN(\u7_mem[0] [20]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_12409),
    .QN(\u7_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_66813),
    .QN(\u7_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_12408),
    .QN(\u7_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_12406),
    .QN(\u7_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_12424),
    .QN(\u7_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_12423),
    .QN(\u7_mem[0] [26]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_12422),
    .QN(\u7_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_12425),
    .QN(\u7_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_12420),
    .QN(\u7_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_12433),
    .QN(\u7_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_12421),
    .QN(\u7_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_12407),
    .QN(\u7_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_12432),
    .QN(\u7_mem[0] [3]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_68215),
    .QN(\u7_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_12415),
    .QN(\u7_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_12435),
    .QN(\u7_mem[0] [6]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_12434),
    .QN(\u7_mem[0] [7]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_12417),
    .QN(\u7_mem[0] [8]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_12431),
    .QN(\u7_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_50225),
    .QN(\u7_mem[1] [0]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_66833),
    .QN(\u7_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_50229),
    .QN(\u7_mem[1] [11]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_50231),
    .QN(\u7_mem[1] [12]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_50242),
    .QN(\u7_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_50240),
    .QN(\u7_mem[1] [14]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_50233),
    .QN(\u7_mem[1] [15]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_50245),
    .QN(\u7_mem[1] [16]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_50235),
    .QN(\u7_mem[1] [17]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_50228),
    .QN(\u7_mem[1] [18]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_50232),
    .QN(\u7_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_50219),
    .QN(\u7_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_50237),
    .QN(\u7_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_50221),
    .QN(\u7_mem[1] [21]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_66809),
    .QN(\u7_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_50238),
    .QN(\u7_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_50241),
    .QN(\u7_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_50227),
    .QN(\u7_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_50243),
    .QN(\u7_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_50224),
    .QN(\u7_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_50251),
    .QN(\u7_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_50222),
    .QN(\u7_mem[1] [29]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_50239),
    .QN(\u7_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_50226),
    .QN(\u7_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_50250),
    .QN(\u7_mem[1] [31]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_50247),
    .QN(\u7_mem[1] [3]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_68221),
    .QN(\u7_mem[1] [4]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_50223),
    .QN(\u7_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_50236),
    .QN(\u7_mem[1] [6]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_50234),
    .QN(\u7_mem[1] [7]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_50246),
    .QN(\u7_mem[1] [8]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_50230),
    .QN(\u7_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_10919),
    .QN(\u7_mem[2] [0]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_9930),
    .QN(\u7_mem[2] [10]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_10017),
    .QN(\u7_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_10046),
    .QN(\u7_mem[2] [12]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_10103),
    .QN(\u7_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_9755),
    .QN(\u7_mem[2] [14]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_9784),
    .QN(\u7_mem[2] [15]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_10132),
    .QN(\u7_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_10160),
    .QN(\u7_mem[2] [17]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_10186),
    .QN(\u7_mem[2] [18]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_10213),
    .QN(\u7_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_10895),
    .QN(\u7_mem[2] [1]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_10240),
    .QN(\u7_mem[2] [20]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_10267),
    .QN(\u7_mem[2] [21]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_66802),
    .QN(\u7_mem[2] [22]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_10323),
    .QN(\u7_mem[2] [23]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_10429),
    .QN(\u7_mem[2] [24]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_10455),
    .QN(\u7_mem[2] [25]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_10481),
    .QN(\u7_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_10506),
    .QN(\u7_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_10377),
    .QN(\u7_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_10680),
    .QN(\u7_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_9843),
    .QN(\u7_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_10656),
    .QN(\u7_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_10350),
    .QN(\u7_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_9873),
    .QN(\u7_mem[2] [3]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_69016),
    .QN(\u7_mem[2] [4]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_10075),
    .QN(\u7_mem[2] [5]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_9726),
    .QN(\u7_mem[2] [6]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_9814),
    .QN(\u7_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_9902),
    .QN(\u7_mem[2] [8]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_9957),
    .QN(\u7_mem[2] [9]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_25381),
    .QN(\u7_mem[3] [0]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_3717),
    .QN(\u7_mem[3] [10]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_3716),
    .QN(\u7_mem[3] [11]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_14030),
    .QN(\u7_mem[3] [12]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_3714),
    .QN(\u7_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_3713),
    .QN(\u7_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_3712),
    .QN(\u7_mem[3] [15]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_43533),
    .QN(\u7_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_3710),
    .QN(\u7_mem[3] [17]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_3709),
    .QN(\u7_mem[3] [18]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_25382),
    .QN(\u7_mem[3] [19]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_25390),
    .QN(\u7_mem[3] [1]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_25388),
    .QN(\u7_mem[3] [20]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_25383),
    .QN(\u7_mem[3] [21]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_25391),
    .QN(\u7_mem[3] [22]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_25389),
    .QN(\u7_mem[3] [23]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_25394),
    .QN(\u7_mem[3] [24]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_25395),
    .QN(\u7_mem[3] [25]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_25379),
    .QN(\u7_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_25380),
    .QN(\u7_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_25386),
    .QN(\u7_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_25385),
    .QN(\u7_mem[3] [29]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_25392),
    .QN(\u7_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_25384),
    .QN(\u7_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u7_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_25393),
    .QN(\u7_mem[3] [31]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_11259),
    .QN(\u7_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_69026),
    .QN(\u7_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_3722),
    .QN(\u7_mem[3] [5]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_3721),
    .QN(\u7_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_3720),
    .QN(\u7_mem[3] [7]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_3719),
    .QN(\u7_mem[3] [8]));
 DFFHQNx1_ASAP7_75t_SL \u7_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_3718),
    .QN(\u7_mem[3] [9]));
 SDFHx1_ASAP7_75t_SL \u7_rp_reg[0]  (.CLK(clk_i),
    .QN(u7_rp[0]),
    .D(n_52770),
    .SE(u7_rp[0]),
    .SI(n_4443));
 DFFHQx4_ASAP7_75t_SL \u7_rp_reg[1]  (.CLK(clk_i),
    .D(n_16899),
    .Q(u7_rp[1]));
 DFFHQx4_ASAP7_75t_SL \u7_rp_reg[2]  (.CLK(clk_i),
    .D(n_4644),
    .Q(u7_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u7_rp_reg[3]  (.CLK(clk_i),
    .D(n_43607),
    .QN(u7_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u7_status_reg[0]  (.CLK(clk_i),
    .D(n_1372),
    .QN(o8_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u7_status_reg[1]  (.CLK(clk_i),
    .D(n_17672),
    .QN(o8_status[1]));
 DFFHQx4_ASAP7_75t_SL \u7_wp_reg[0]  (.CLK(clk_i),
    .D(n_57760),
    .Q(u7_wp[0]));
 DFFHQNx2_ASAP7_75t_SL \u7_wp_reg[1]  (.CLK(clk_i),
    .D(n_33112),
    .QN(u7_wp[1]));
 DFFHQNx1_ASAP7_75t_SL \u7_wp_reg[2]  (.CLK(clk_i),
    .D(n_3077),
    .QN(u7_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[0]  (.CLK(clk_i),
    .D(n_73302),
    .QN(out_slt9[0]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[10]  (.CLK(clk_i),
    .D(n_43282),
    .QN(out_slt9[10]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[11]  (.CLK(clk_i),
    .D(n_50707),
    .QN(out_slt9[11]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[12]  (.CLK(clk_i),
    .D(n_5093),
    .QN(out_slt9[12]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[13]  (.CLK(clk_i),
    .D(n_14425),
    .QN(out_slt9[13]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[14]  (.CLK(clk_i),
    .D(n_73308),
    .QN(out_slt9[14]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[15]  (.CLK(clk_i),
    .D(n_50541),
    .QN(out_slt9[15]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[16]  (.CLK(clk_i),
    .D(n_7999),
    .QN(out_slt9[16]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[17]  (.CLK(clk_i),
    .D(n_7744),
    .QN(out_slt9[17]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[18]  (.CLK(clk_i),
    .D(n_4990),
    .QN(out_slt9[18]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[19]  (.CLK(clk_i),
    .D(n_72308),
    .QN(out_slt9[19]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[1]  (.CLK(clk_i),
    .D(n_73303),
    .QN(out_slt9[1]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[2]  (.CLK(clk_i),
    .D(n_40905),
    .QN(out_slt9[2]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[3]  (.CLK(clk_i),
    .D(n_4798),
    .QN(out_slt9[3]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[4]  (.CLK(clk_i),
    .D(n_73311),
    .QN(out_slt9[4]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[5]  (.CLK(clk_i),
    .D(n_73314),
    .QN(out_slt9[5]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[6]  (.CLK(clk_i),
    .D(n_73309),
    .QN(out_slt9[6]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[7]  (.CLK(clk_i),
    .D(n_73310),
    .QN(out_slt9[7]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[8]  (.CLK(clk_i),
    .D(n_5087),
    .QN(out_slt9[8]));
 DFFHQNx2_ASAP7_75t_SL \u8_dout_reg[9]  (.CLK(clk_i),
    .D(n_5088),
    .QN(out_slt9[9]));
 DFFHQNx1_ASAP7_75t_SL u8_empty_reg (.CLK(clk_i),
    .D(n_31455),
    .QN(o9_empty));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_10923),
    .QN(\u8_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_66818),
    .QN(\u8_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_10019),
    .QN(\u8_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_10048),
    .QN(\u8_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_10105),
    .QN(\u8_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_9757),
    .QN(\u8_mem[0] [14]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_9786),
    .QN(\u8_mem[0] [15]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_10134),
    .QN(\u8_mem[0] [16]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_10162),
    .QN(\u8_mem[0] [17]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_10188),
    .QN(\u8_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_10215),
    .QN(\u8_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_10906),
    .QN(\u8_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_10242),
    .QN(\u8_mem[0] [20]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_10269),
    .QN(\u8_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_66806),
    .QN(\u8_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_10326),
    .QN(\u8_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_10431),
    .QN(\u8_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_10457),
    .QN(\u8_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_10483),
    .QN(\u8_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_10509),
    .QN(\u8_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_10379),
    .QN(\u8_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_10665),
    .QN(\u8_mem[0] [29]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_9838),
    .QN(\u8_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_10644),
    .QN(\u8_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_10352),
    .QN(\u8_mem[0] [31]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_9867),
    .QN(\u8_mem[0] [3]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_69011),
    .QN(\u8_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_10069),
    .QN(\u8_mem[0] [5]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_9721),
    .QN(\u8_mem[0] [6]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_9808),
    .QN(\u8_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_9896),
    .QN(\u8_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_9959),
    .QN(\u8_mem[0] [9]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_75736),
    .QN(\u8_mem[1] [0]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_66822),
    .QN(\u8_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_40992),
    .QN(\u8_mem[1] [11]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_40983),
    .QN(\u8_mem[1] [12]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_40985),
    .QN(\u8_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_40989),
    .QN(\u8_mem[1] [14]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_40982),
    .QN(\u8_mem[1] [15]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_16314),
    .QN(\u8_mem[1] [16]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_46289),
    .QN(\u8_mem[1] [17]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_73400),
    .QN(\u8_mem[1] [18]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_10203),
    .QN(\u8_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_40993),
    .QN(\u8_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_15931),
    .QN(\u8_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_73999),
    .QN(\u8_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_16680),
    .QN(\u8_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_16684),
    .QN(\u8_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_15927),
    .QN(\u8_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_15915),
    .QN(\u8_mem[1] [25]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_10470),
    .QN(\u8_mem[1] [26]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_10496),
    .QN(\u8_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_10369),
    .QN(\u8_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_22718),
    .QN(\u8_mem[1] [29]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_40986),
    .QN(\u8_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_47403),
    .QN(\u8_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_15923),
    .QN(\u8_mem[1] [31]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_15869),
    .QN(\u8_mem[1] [3]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_68217),
    .QN(\u8_mem[1] [4]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_40990),
    .QN(\u8_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_49387),
    .QN(\u8_mem[1] [6]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_40987),
    .QN(\u8_mem[1] [7]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_40988),
    .QN(\u8_mem[1] [8]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_73388),
    .QN(\u8_mem[1] [9]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_10922),
    .QN(\u8_mem[2] [0]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_9926),
    .QN(\u8_mem[2] [10]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_10013),
    .QN(\u8_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_10042),
    .QN(\u8_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_10099),
    .QN(\u8_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_9751),
    .QN(\u8_mem[2] [14]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_9780),
    .QN(\u8_mem[2] [15]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_10128),
    .QN(\u8_mem[2] [16]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_10156),
    .QN(\u8_mem[2] [17]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_10182),
    .QN(\u8_mem[2] [18]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_10209),
    .QN(\u8_mem[2] [19]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_10892),
    .QN(\u8_mem[2] [1]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_10227),
    .QN(\u8_mem[2] [20]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_10254),
    .QN(\u8_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_66808),
    .QN(\u8_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_10306),
    .QN(\u8_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_10413),
    .QN(\u8_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_10439),
    .QN(\u8_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_10464),
    .QN(\u8_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_10490),
    .QN(\u8_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_10363),
    .QN(\u8_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_10666),
    .QN(\u8_mem[2] [29]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_9840),
    .QN(\u8_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_10642),
    .QN(\u8_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_10336),
    .QN(\u8_mem[2] [31]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_9869),
    .QN(\u8_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_69014),
    .QN(\u8_mem[2] [4]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_10071),
    .QN(\u8_mem[2] [5]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_9722),
    .QN(\u8_mem[2] [6]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_9810),
    .QN(\u8_mem[2] [7]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_9898),
    .QN(\u8_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_9954),
    .QN(\u8_mem[2] [9]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_22508),
    .QN(\u8_mem[3] [0]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_17801),
    .QN(\u8_mem[3] [10]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_18060),
    .QN(\u8_mem[3] [11]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_18491),
    .QN(\u8_mem[3] [12]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_17778),
    .QN(\u8_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_18195),
    .QN(\u8_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_18448),
    .QN(\u8_mem[3] [15]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_17787),
    .QN(\u8_mem[3] [16]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_11197),
    .QN(\u8_mem[3] [17]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_23971),
    .QN(\u8_mem[3] [18]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_11212),
    .QN(\u8_mem[3] [19]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_3900),
    .QN(\u8_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_47415),
    .QN(\u8_mem[3] [20]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_47261),
    .QN(\u8_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_47348),
    .QN(\u8_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_47340),
    .QN(\u8_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_47373),
    .QN(\u8_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_47184),
    .QN(\u8_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_47287),
    .QN(\u8_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_47192),
    .QN(\u8_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_47157),
    .QN(\u8_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_47266),
    .QN(\u8_mem[3] [29]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_18289),
    .QN(\u8_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_47121),
    .QN(\u8_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_47217),
    .QN(\u8_mem[3] [31]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_18058),
    .QN(\u8_mem[3] [3]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_68212),
    .QN(\u8_mem[3] [4]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_17979),
    .QN(\u8_mem[3] [5]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_17809),
    .QN(\u8_mem[3] [6]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_18018),
    .QN(\u8_mem[3] [7]));
 DFFHQNx2_ASAP7_75t_SL \u8_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_17785),
    .QN(\u8_mem[3] [8]));
 DFFHQNx1_ASAP7_75t_SL \u8_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_17938),
    .QN(\u8_mem[3] [9]));
 SDFHx4_ASAP7_75t_SL \u8_rp_reg[0]  (.CLK(clk_i),
    .D(n_79204),
    .QN(u8_rp[0]),
    .SE(u8_rp[0]),
    .SI(n_4439));
 DFFHQx4_ASAP7_75t_SL \u8_rp_reg[1]  (.CLK(clk_i),
    .D(n_78141),
    .Q(u8_rp[1]));
 DFFHQx4_ASAP7_75t_SL \u8_rp_reg[2]  (.CLK(clk_i),
    .D(n_72061),
    .Q(u8_rp[2]));
 DFFHQNx2_ASAP7_75t_SL \u8_rp_reg[3]  (.CLK(clk_i),
    .D(n_31191),
    .QN(u8_rp[3]));
 DFFHQNx1_ASAP7_75t_SL \u8_status_reg[0]  (.CLK(clk_i),
    .D(n_78935),
    .QN(o9_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u8_status_reg[1]  (.CLK(clk_i),
    .D(n_58150),
    .QN(o9_status[1]));
 DFFHQx4_ASAP7_75t_SL \u8_wp_reg[0]  (.CLK(clk_i),
    .D(n_2984),
    .Q(u8_wp[0]));
 DFFHQNx1_ASAP7_75t_SL \u8_wp_reg[1]  (.CLK(clk_i),
    .D(n_40994),
    .QN(u8_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u8_wp_reg[2]  (.CLK(clk_i),
    .D(n_72909),
    .QN(u8_wp[2]));
 DFFHQNx2_ASAP7_75t_SL \u9_din_tmp1_reg[0]  (.CLK(clk_i),
    .D(n_29554),
    .QN(u9_din_tmp1[0]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[10]  (.CLK(clk_i),
    .D(n_34499),
    .QN(u9_din_tmp1[10]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[11]  (.CLK(clk_i),
    .D(n_34503),
    .QN(u9_din_tmp1[11]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[12]  (.CLK(clk_i),
    .D(n_29558),
    .QN(u9_din_tmp1[12]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[13]  (.CLK(clk_i),
    .D(n_34507),
    .QN(u9_din_tmp1[13]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[14]  (.CLK(clk_i),
    .D(n_29534),
    .QN(u9_din_tmp1[14]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[15]  (.CLK(clk_i),
    .D(n_29532),
    .QN(u9_din_tmp1[15]));
 DFFHQNx2_ASAP7_75t_SL \u9_din_tmp1_reg[1]  (.CLK(clk_i),
    .D(n_29556),
    .QN(u9_din_tmp1[1]));
 DFFHQNx2_ASAP7_75t_SL \u9_din_tmp1_reg[2]  (.CLK(clk_i),
    .D(n_29528),
    .QN(u9_din_tmp1[2]));
 DFFHQNx2_ASAP7_75t_SL \u9_din_tmp1_reg[3]  (.CLK(clk_i),
    .D(n_29530),
    .QN(u9_din_tmp1[3]));
 DFFHQNx2_ASAP7_75t_SL \u9_din_tmp1_reg[4]  (.CLK(clk_i),
    .D(n_34491),
    .QN(u9_din_tmp1[4]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[5]  (.CLK(clk_i),
    .D(n_29550),
    .QN(u9_din_tmp1[5]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[6]  (.CLK(clk_i),
    .D(n_29548),
    .QN(u9_din_tmp1[6]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[7]  (.CLK(clk_i),
    .D(n_29546),
    .QN(u9_din_tmp1[7]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[8]  (.CLK(clk_i),
    .D(n_29544),
    .QN(u9_din_tmp1[8]));
 DFFHQNx1_ASAP7_75t_SL \u9_din_tmp1_reg[9]  (.CLK(clk_i),
    .D(n_34495),
    .QN(u9_din_tmp1[9]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[0]  (.CLK(clk_i),
    .D(n_1629),
    .Q(i3_dout[0]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[10]  (.CLK(clk_i),
    .D(n_1620),
    .Q(i3_dout[10]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[11]  (.CLK(clk_i),
    .D(n_1619),
    .Q(i3_dout[11]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[12]  (.CLK(clk_i),
    .D(n_1618),
    .Q(i3_dout[12]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[13]  (.CLK(clk_i),
    .D(n_1617),
    .Q(i3_dout[13]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[14]  (.CLK(clk_i),
    .D(n_1616),
    .Q(i3_dout[14]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[15]  (.CLK(clk_i),
    .D(n_1615),
    .Q(i3_dout[15]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[16]  (.CLK(clk_i),
    .D(n_1614),
    .Q(i3_dout[16]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[17]  (.CLK(clk_i),
    .D(n_1530),
    .Q(i3_dout[17]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[18]  (.CLK(clk_i),
    .D(n_1613),
    .Q(i3_dout[18]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[19]  (.CLK(clk_i),
    .D(n_1612),
    .Q(i3_dout[19]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[1]  (.CLK(clk_i),
    .D(n_1628),
    .Q(i3_dout[1]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[20]  (.CLK(clk_i),
    .D(n_1611),
    .Q(i3_dout[20]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[21]  (.CLK(clk_i),
    .D(n_1609),
    .Q(i3_dout[21]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[22]  (.CLK(clk_i),
    .D(n_1608),
    .Q(i3_dout[22]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[23]  (.CLK(clk_i),
    .D(n_1547),
    .Q(i3_dout[23]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[24]  (.CLK(clk_i),
    .D(n_1607),
    .Q(i3_dout[24]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[25]  (.CLK(clk_i),
    .D(n_1606),
    .Q(i3_dout[25]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[26]  (.CLK(clk_i),
    .D(n_1605),
    .Q(i3_dout[26]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[27]  (.CLK(clk_i),
    .D(n_1604),
    .Q(i3_dout[27]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[28]  (.CLK(clk_i),
    .D(n_1603),
    .Q(i3_dout[28]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[29]  (.CLK(clk_i),
    .D(n_1602),
    .Q(i3_dout[29]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[2]  (.CLK(clk_i),
    .D(n_1627),
    .Q(i3_dout[2]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[30]  (.CLK(clk_i),
    .D(n_1601),
    .Q(i3_dout[30]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[31]  (.CLK(clk_i),
    .D(n_1600),
    .Q(i3_dout[31]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[3]  (.CLK(clk_i),
    .D(n_1626),
    .Q(i3_dout[3]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[4]  (.CLK(clk_i),
    .D(n_1625),
    .Q(i3_dout[4]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[5]  (.CLK(clk_i),
    .D(n_1624),
    .Q(i3_dout[5]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[6]  (.CLK(clk_i),
    .D(n_1623),
    .Q(i3_dout[6]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[7]  (.CLK(clk_i),
    .D(n_1622),
    .Q(i3_dout[7]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[8]  (.CLK(clk_i),
    .D(n_1621),
    .Q(i3_dout[8]));
 DFFHQx4_ASAP7_75t_SL \u9_dout_reg[9]  (.CLK(clk_i),
    .D(n_1531),
    .Q(i3_dout[9]));
 DFFHQNx1_ASAP7_75t_SL u9_empty_reg (.CLK(clk_i),
    .D(n_48632),
    .QN(i3_empty));
 DFFHQNx1_ASAP7_75t_SL u9_full_reg (.CLK(clk_i),
    .D(n_50427),
    .QN(i3_full));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][0]  (.CLK(clk_i),
    .D(n_46588),
    .QN(\u9_mem[0] [0]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][10]  (.CLK(clk_i),
    .D(n_5008),
    .QN(\u9_mem[0] [10]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][11]  (.CLK(clk_i),
    .D(n_5009),
    .QN(\u9_mem[0] [11]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][12]  (.CLK(clk_i),
    .D(n_5010),
    .QN(\u9_mem[0] [12]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][13]  (.CLK(clk_i),
    .D(n_5011),
    .QN(\u9_mem[0] [13]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][14]  (.CLK(clk_i),
    .D(n_5012),
    .QN(\u9_mem[0] [14]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][15]  (.CLK(clk_i),
    .D(n_5014),
    .QN(\u9_mem[0] [15]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][16]  (.CLK(clk_i),
    .D(n_5015),
    .QN(\u9_mem[0] [16]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][17]  (.CLK(clk_i),
    .D(n_5016),
    .QN(\u9_mem[0] [17]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][18]  (.CLK(clk_i),
    .D(n_17927),
    .QN(\u9_mem[0] [18]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][19]  (.CLK(clk_i),
    .D(n_5020),
    .QN(\u9_mem[0] [19]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][1]  (.CLK(clk_i),
    .D(n_4998),
    .QN(\u9_mem[0] [1]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][20]  (.CLK(clk_i),
    .D(n_4876),
    .QN(\u9_mem[0] [20]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][21]  (.CLK(clk_i),
    .D(n_4873),
    .QN(\u9_mem[0] [21]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][22]  (.CLK(clk_i),
    .D(n_4872),
    .QN(\u9_mem[0] [22]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][23]  (.CLK(clk_i),
    .D(n_4871),
    .QN(\u9_mem[0] [23]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][24]  (.CLK(clk_i),
    .D(n_4868),
    .QN(\u9_mem[0] [24]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][25]  (.CLK(clk_i),
    .D(n_4867),
    .QN(\u9_mem[0] [25]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][26]  (.CLK(clk_i),
    .D(n_4865),
    .QN(\u9_mem[0] [26]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][27]  (.CLK(clk_i),
    .D(n_4864),
    .QN(\u9_mem[0] [27]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][28]  (.CLK(clk_i),
    .D(n_4862),
    .QN(\u9_mem[0] [28]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][29]  (.CLK(clk_i),
    .D(n_4861),
    .QN(\u9_mem[0] [29]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][2]  (.CLK(clk_i),
    .D(n_4999),
    .QN(\u9_mem[0] [2]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][30]  (.CLK(clk_i),
    .D(n_4859),
    .QN(\u9_mem[0] [30]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][31]  (.CLK(clk_i),
    .D(n_4858),
    .QN(\u9_mem[0] [31]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][3]  (.CLK(clk_i),
    .D(n_5000),
    .QN(\u9_mem[0] [3]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][4]  (.CLK(clk_i),
    .D(n_5002),
    .QN(\u9_mem[0] [4]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][5]  (.CLK(clk_i),
    .D(n_5003),
    .QN(\u9_mem[0] [5]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][6]  (.CLK(clk_i),
    .D(n_5004),
    .QN(\u9_mem[0] [6]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][7]  (.CLK(clk_i),
    .D(n_5005),
    .QN(\u9_mem[0] [7]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][8]  (.CLK(clk_i),
    .D(n_24891),
    .QN(\u9_mem[0] [8]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[0][9]  (.CLK(clk_i),
    .D(n_5007),
    .QN(\u9_mem[0] [9]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][0]  (.CLK(clk_i),
    .D(n_5121),
    .QN(\u9_mem[1] [0]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][10]  (.CLK(clk_i),
    .D(n_5143),
    .QN(\u9_mem[1] [10]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][11]  (.CLK(clk_i),
    .D(n_22694),
    .QN(\u9_mem[1] [11]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][12]  (.CLK(clk_i),
    .D(n_22629),
    .QN(\u9_mem[1] [12]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][13]  (.CLK(clk_i),
    .D(n_5149),
    .QN(\u9_mem[1] [13]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][14]  (.CLK(clk_i),
    .D(n_5152),
    .QN(\u9_mem[1] [14]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][15]  (.CLK(clk_i),
    .D(n_5153),
    .QN(\u9_mem[1] [15]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][16]  (.CLK(clk_i),
    .D(n_5154),
    .QN(\u9_mem[1] [16]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][17]  (.CLK(clk_i),
    .D(n_5156),
    .QN(\u9_mem[1] [17]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][18]  (.CLK(clk_i),
    .D(n_5157),
    .QN(\u9_mem[1] [18]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][19]  (.CLK(clk_i),
    .D(n_5158),
    .QN(\u9_mem[1] [19]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][1]  (.CLK(clk_i),
    .D(n_60874),
    .QN(\u9_mem[1] [1]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][20]  (.CLK(clk_i),
    .D(n_5195),
    .QN(\u9_mem[1] [20]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][21]  (.CLK(clk_i),
    .D(n_5196),
    .QN(\u9_mem[1] [21]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][22]  (.CLK(clk_i),
    .D(n_5197),
    .QN(\u9_mem[1] [22]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][23]  (.CLK(clk_i),
    .D(n_5198),
    .QN(\u9_mem[1] [23]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][24]  (.CLK(clk_i),
    .D(n_5199),
    .QN(\u9_mem[1] [24]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][25]  (.CLK(clk_i),
    .D(n_5200),
    .QN(\u9_mem[1] [25]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][26]  (.CLK(clk_i),
    .D(n_5201),
    .QN(\u9_mem[1] [26]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][27]  (.CLK(clk_i),
    .D(n_5202),
    .QN(\u9_mem[1] [27]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][28]  (.CLK(clk_i),
    .D(n_5203),
    .QN(\u9_mem[1] [28]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][29]  (.CLK(clk_i),
    .D(n_5204),
    .QN(\u9_mem[1] [29]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][2]  (.CLK(clk_i),
    .D(n_5125),
    .QN(\u9_mem[1] [2]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][30]  (.CLK(clk_i),
    .D(n_5207),
    .QN(\u9_mem[1] [30]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][31]  (.CLK(clk_i),
    .D(n_5208),
    .QN(\u9_mem[1] [31]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][3]  (.CLK(clk_i),
    .D(n_5127),
    .QN(\u9_mem[1] [3]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][4]  (.CLK(clk_i),
    .D(n_5129),
    .QN(\u9_mem[1] [4]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][5]  (.CLK(clk_i),
    .D(n_22635),
    .QN(\u9_mem[1] [5]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][6]  (.CLK(clk_i),
    .D(n_5133),
    .QN(\u9_mem[1] [6]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][7]  (.CLK(clk_i),
    .D(n_5135),
    .QN(\u9_mem[1] [7]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][8]  (.CLK(clk_i),
    .D(n_24892),
    .QN(\u9_mem[1] [8]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[1][9]  (.CLK(clk_i),
    .D(n_5139),
    .QN(\u9_mem[1] [9]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][0]  (.CLK(clk_i),
    .D(n_12896),
    .QN(\u9_mem[2] [0]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][10]  (.CLK(clk_i),
    .D(n_12889),
    .QN(\u9_mem[2] [10]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][11]  (.CLK(clk_i),
    .D(n_12893),
    .QN(\u9_mem[2] [11]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][12]  (.CLK(clk_i),
    .D(n_12902),
    .QN(\u9_mem[2] [12]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][13]  (.CLK(clk_i),
    .D(n_12892),
    .QN(\u9_mem[2] [13]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][14]  (.CLK(clk_i),
    .D(n_12875),
    .QN(\u9_mem[2] [14]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][15]  (.CLK(clk_i),
    .D(n_12895),
    .QN(\u9_mem[2] [15]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][16]  (.CLK(clk_i),
    .D(n_12874),
    .QN(\u9_mem[2] [16]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][17]  (.CLK(clk_i),
    .D(n_12891),
    .QN(\u9_mem[2] [17]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][18]  (.CLK(clk_i),
    .D(n_12888),
    .QN(\u9_mem[2] [18]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][19]  (.CLK(clk_i),
    .D(n_12870),
    .QN(\u9_mem[2] [19]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][1]  (.CLK(clk_i),
    .D(n_12897),
    .QN(\u9_mem[2] [1]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][20]  (.CLK(clk_i),
    .D(n_12886),
    .QN(\u9_mem[2] [20]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][21]  (.CLK(clk_i),
    .D(n_12885),
    .QN(\u9_mem[2] [21]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][22]  (.CLK(clk_i),
    .D(n_12884),
    .QN(\u9_mem[2] [22]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][23]  (.CLK(clk_i),
    .D(n_12883),
    .QN(\u9_mem[2] [23]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][24]  (.CLK(clk_i),
    .D(n_12882),
    .QN(\u9_mem[2] [24]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][25]  (.CLK(clk_i),
    .D(n_12881),
    .QN(\u9_mem[2] [25]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][26]  (.CLK(clk_i),
    .D(n_12880),
    .QN(\u9_mem[2] [26]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][27]  (.CLK(clk_i),
    .D(n_12879),
    .QN(\u9_mem[2] [27]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][28]  (.CLK(clk_i),
    .D(n_12872),
    .QN(\u9_mem[2] [28]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][29]  (.CLK(clk_i),
    .D(n_12878),
    .QN(\u9_mem[2] [29]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][2]  (.CLK(clk_i),
    .D(n_12898),
    .QN(\u9_mem[2] [2]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][30]  (.CLK(clk_i),
    .D(n_12877),
    .QN(\u9_mem[2] [30]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][31]  (.CLK(clk_i),
    .D(n_12876),
    .QN(\u9_mem[2] [31]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][3]  (.CLK(clk_i),
    .D(n_12899),
    .QN(\u9_mem[2] [3]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][4]  (.CLK(clk_i),
    .D(n_12887),
    .QN(\u9_mem[2] [4]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][5]  (.CLK(clk_i),
    .D(n_12900),
    .QN(\u9_mem[2] [5]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][6]  (.CLK(clk_i),
    .D(n_12873),
    .QN(\u9_mem[2] [6]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][7]  (.CLK(clk_i),
    .D(n_12901),
    .QN(\u9_mem[2] [7]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][8]  (.CLK(clk_i),
    .D(n_24890),
    .QN(\u9_mem[2] [8]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[2][9]  (.CLK(clk_i),
    .D(n_12890),
    .QN(\u9_mem[2] [9]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][0]  (.CLK(clk_i),
    .D(n_5118),
    .QN(\u9_mem[3] [0]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][10]  (.CLK(clk_i),
    .D(n_21536),
    .QN(\u9_mem[3] [10]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][11]  (.CLK(clk_i),
    .D(n_15694),
    .QN(\u9_mem[3] [11]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][12]  (.CLK(clk_i),
    .D(n_5106),
    .QN(\u9_mem[3] [12]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][13]  (.CLK(clk_i),
    .D(n_5105),
    .QN(\u9_mem[3] [13]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][14]  (.CLK(clk_i),
    .D(n_5104),
    .QN(\u9_mem[3] [14]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][15]  (.CLK(clk_i),
    .D(n_5103),
    .QN(\u9_mem[3] [15]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][16]  (.CLK(clk_i),
    .D(n_5101),
    .QN(\u9_mem[3] [16]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][17]  (.CLK(clk_i),
    .D(n_5100),
    .QN(\u9_mem[3] [17]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][18]  (.CLK(clk_i),
    .D(n_49626),
    .QN(\u9_mem[3] [18]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][19]  (.CLK(clk_i),
    .D(n_5212),
    .QN(\u9_mem[3] [19]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][1]  (.CLK(clk_i),
    .D(n_22432),
    .QN(\u9_mem[3] [1]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][20]  (.CLK(clk_i),
    .D(n_5159),
    .QN(\u9_mem[3] [20]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][21]  (.CLK(clk_i),
    .D(n_5160),
    .QN(\u9_mem[3] [21]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][22]  (.CLK(clk_i),
    .D(n_5161),
    .QN(\u9_mem[3] [22]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][23]  (.CLK(clk_i),
    .D(n_22407),
    .QN(\u9_mem[3] [23]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][24]  (.CLK(clk_i),
    .D(n_22413),
    .QN(\u9_mem[3] [24]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][25]  (.CLK(clk_i),
    .D(n_22964),
    .QN(\u9_mem[3] [25]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][26]  (.CLK(clk_i),
    .D(n_5172),
    .QN(\u9_mem[3] [26]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][27]  (.CLK(clk_i),
    .D(n_5178),
    .QN(\u9_mem[3] [27]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][28]  (.CLK(clk_i),
    .D(n_22415),
    .QN(\u9_mem[3] [28]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][29]  (.CLK(clk_i),
    .D(n_22424),
    .QN(\u9_mem[3] [29]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][2]  (.CLK(clk_i),
    .D(n_46559),
    .QN(\u9_mem[3] [2]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][30]  (.CLK(clk_i),
    .D(n_22482),
    .QN(\u9_mem[3] [30]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][31]  (.CLK(clk_i),
    .D(n_22430),
    .QN(\u9_mem[3] [31]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][3]  (.CLK(clk_i),
    .D(n_46563),
    .QN(\u9_mem[3] [3]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][4]  (.CLK(clk_i),
    .D(n_5114),
    .QN(\u9_mem[3] [4]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][5]  (.CLK(clk_i),
    .D(n_5113),
    .QN(\u9_mem[3] [5]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][6]  (.CLK(clk_i),
    .D(n_5112),
    .QN(\u9_mem[3] [6]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][7]  (.CLK(clk_i),
    .D(n_5111),
    .QN(\u9_mem[3] [7]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][8]  (.CLK(clk_i),
    .D(n_24889),
    .QN(\u9_mem[3] [8]));
 DFFHQNx2_ASAP7_75t_SL \u9_mem_reg[3][9]  (.CLK(clk_i),
    .D(n_21532),
    .QN(\u9_mem[3] [9]));
 DFFHQx4_ASAP7_75t_SL \u9_rp_reg[0]  (.CLK(clk_i),
    .D(n_2708),
    .Q(u9_rp[0]));
 DFFHQNx2_ASAP7_75t_SL \u9_rp_reg[1]  (.CLK(clk_i),
    .D(n_11513),
    .QN(u9_rp[1]));
 DFFHQNx2_ASAP7_75t_SL \u9_rp_reg[2]  (.CLK(clk_i),
    .D(n_2956),
    .QN(u9_rp[2]));
 DFFHQNx1_ASAP7_75t_SL \u9_status_reg[0]  (.CLK(clk_i),
    .D(n_703),
    .QN(i3_status[0]));
 DFFHQNx1_ASAP7_75t_SL \u9_status_reg[1]  (.CLK(clk_i),
    .D(n_21599),
    .QN(i3_status[1]));
 DFFHQNx1_ASAP7_75t_SL \u9_wp_reg[0]  (.CLK(clk_i),
    .D(n_4826),
    .QN(u9_wp[0]));
 DFFHQx4_ASAP7_75t_SL \u9_wp_reg[1]  (.CLK(clk_i),
    .D(n_24733),
    .Q(u9_wp[1]));
 DFFHQNx2_ASAP7_75t_SL \u9_wp_reg[2]  (.CLK(clk_i),
    .D(n_21264),
    .QN(u9_wp[2]));
 DFFHQx4_ASAP7_75t_SL \u9_wp_reg[3]  (.CLK(clk_i),
    .D(n_4827),
    .Q(u9_wp[3]));
 DFFHQNx1_ASAP7_75t_R valid_s1_reg (.CLK(clk_i),
    .D(n_2190),
    .QN(valid_s1));
 DFFHQNx1_ASAP7_75t_SL valid_s_reg (.CLK(clk_i),
    .D(n_2571),
    .QN(valid_s));
endmodule
